magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755253277
<< metal1 >>
rect 1152 84692 20352 84716
rect 1152 84652 3688 84692
rect 3728 84652 3770 84692
rect 3810 84652 3852 84692
rect 3892 84652 3934 84692
rect 3974 84652 4016 84692
rect 4056 84652 18808 84692
rect 18848 84652 18890 84692
rect 18930 84652 18972 84692
rect 19012 84652 19054 84692
rect 19094 84652 19136 84692
rect 19176 84652 20352 84692
rect 1152 84628 20352 84652
rect 4299 84440 4341 84449
rect 4299 84400 4300 84440
rect 4340 84400 4341 84440
rect 4299 84391 4341 84400
rect 4483 84356 4541 84357
rect 4483 84316 4492 84356
rect 4532 84316 4541 84356
rect 4483 84315 4541 84316
rect 1152 83936 20452 83960
rect 1152 83896 4928 83936
rect 4968 83896 5010 83936
rect 5050 83896 5092 83936
rect 5132 83896 5174 83936
rect 5214 83896 5256 83936
rect 5296 83896 20048 83936
rect 20088 83896 20130 83936
rect 20170 83896 20212 83936
rect 20252 83896 20294 83936
rect 20334 83896 20376 83936
rect 20416 83896 20452 83936
rect 1152 83872 20452 83896
rect 1707 83768 1749 83777
rect 1707 83728 1708 83768
rect 1748 83728 1749 83768
rect 1707 83719 1749 83728
rect 1899 83768 1941 83777
rect 1899 83728 1900 83768
rect 1940 83728 1941 83768
rect 1899 83719 1941 83728
rect 2283 83768 2325 83777
rect 2283 83728 2284 83768
rect 2324 83728 2325 83768
rect 2283 83719 2325 83728
rect 2667 83768 2709 83777
rect 2667 83728 2668 83768
rect 2708 83728 2709 83768
rect 2667 83719 2709 83728
rect 3051 83768 3093 83777
rect 3051 83728 3052 83768
rect 3092 83728 3093 83768
rect 3051 83719 3093 83728
rect 3435 83768 3477 83777
rect 3435 83728 3436 83768
rect 3476 83728 3477 83768
rect 3435 83719 3477 83728
rect 3819 83768 3861 83777
rect 3819 83728 3820 83768
rect 3860 83728 3861 83768
rect 3819 83719 3861 83728
rect 4203 83768 4245 83777
rect 4203 83728 4204 83768
rect 4244 83728 4245 83768
rect 4203 83719 4245 83728
rect 4587 83768 4629 83777
rect 4587 83728 4588 83768
rect 4628 83728 4629 83768
rect 4587 83719 4629 83728
rect 4971 83768 5013 83777
rect 4971 83728 4972 83768
rect 5012 83728 5013 83768
rect 4971 83719 5013 83728
rect 5355 83768 5397 83777
rect 5355 83728 5356 83768
rect 5396 83728 5397 83768
rect 5355 83719 5397 83728
rect 5931 83768 5973 83777
rect 5931 83728 5932 83768
rect 5972 83728 5973 83768
rect 5931 83719 5973 83728
rect 6699 83768 6741 83777
rect 6699 83728 6700 83768
rect 6740 83728 6741 83768
rect 6699 83719 6741 83728
rect 7179 83768 7221 83777
rect 7179 83728 7180 83768
rect 7220 83728 7221 83768
rect 7179 83719 7221 83728
rect 7563 83768 7605 83777
rect 7563 83728 7564 83768
rect 7604 83728 7605 83768
rect 7563 83719 7605 83728
rect 7755 83768 7797 83777
rect 7755 83728 7756 83768
rect 7796 83728 7797 83768
rect 7755 83719 7797 83728
rect 8331 83768 8373 83777
rect 8331 83728 8332 83768
rect 8372 83728 8373 83768
rect 8331 83719 8373 83728
rect 8523 83768 8565 83777
rect 8523 83728 8524 83768
rect 8564 83728 8565 83768
rect 8523 83719 8565 83728
rect 13323 83768 13365 83777
rect 13323 83728 13324 83768
rect 13364 83728 13365 83768
rect 13323 83719 13365 83728
rect 14955 83768 14997 83777
rect 14955 83728 14956 83768
rect 14996 83728 14997 83768
rect 14955 83719 14997 83728
rect 15531 83768 15573 83777
rect 15531 83728 15532 83768
rect 15572 83728 15573 83768
rect 15531 83719 15573 83728
rect 15723 83768 15765 83777
rect 15723 83728 15724 83768
rect 15764 83728 15765 83768
rect 15723 83719 15765 83728
rect 18123 83768 18165 83777
rect 18123 83728 18124 83768
rect 18164 83728 18165 83768
rect 18123 83719 18165 83728
rect 19179 83768 19221 83777
rect 19179 83728 19180 83768
rect 19220 83728 19221 83768
rect 19179 83719 19221 83728
rect 19563 83768 19605 83777
rect 19563 83728 19564 83768
rect 19604 83728 19605 83768
rect 19563 83719 19605 83728
rect 1507 83516 1565 83517
rect 1507 83476 1516 83516
rect 1556 83476 1565 83516
rect 1507 83475 1565 83476
rect 2083 83516 2141 83517
rect 2083 83476 2092 83516
rect 2132 83476 2141 83516
rect 2083 83475 2141 83476
rect 2467 83516 2525 83517
rect 2467 83476 2476 83516
rect 2516 83476 2525 83516
rect 2467 83475 2525 83476
rect 2851 83516 2909 83517
rect 2851 83476 2860 83516
rect 2900 83476 2909 83516
rect 2851 83475 2909 83476
rect 3235 83516 3293 83517
rect 3235 83476 3244 83516
rect 3284 83476 3293 83516
rect 3235 83475 3293 83476
rect 3619 83516 3677 83517
rect 3619 83476 3628 83516
rect 3668 83476 3677 83516
rect 3619 83475 3677 83476
rect 4003 83516 4061 83517
rect 4003 83476 4012 83516
rect 4052 83476 4061 83516
rect 4003 83475 4061 83476
rect 4387 83516 4445 83517
rect 4387 83476 4396 83516
rect 4436 83476 4445 83516
rect 4387 83475 4445 83476
rect 4771 83516 4829 83517
rect 4771 83476 4780 83516
rect 4820 83476 4829 83516
rect 4771 83475 4829 83476
rect 5155 83516 5213 83517
rect 5155 83476 5164 83516
rect 5204 83476 5213 83516
rect 5155 83475 5213 83476
rect 5539 83516 5597 83517
rect 5539 83476 5548 83516
rect 5588 83476 5597 83516
rect 5539 83475 5597 83476
rect 6115 83516 6173 83517
rect 6115 83476 6124 83516
rect 6164 83476 6173 83516
rect 6115 83475 6173 83476
rect 6499 83516 6557 83517
rect 6499 83476 6508 83516
rect 6548 83476 6557 83516
rect 6499 83475 6557 83476
rect 6979 83516 7037 83517
rect 6979 83476 6988 83516
rect 7028 83476 7037 83516
rect 6979 83475 7037 83476
rect 7363 83516 7421 83517
rect 7363 83476 7372 83516
rect 7412 83476 7421 83516
rect 7363 83475 7421 83476
rect 7939 83516 7997 83517
rect 7939 83476 7948 83516
rect 7988 83476 7997 83516
rect 7939 83475 7997 83476
rect 8131 83516 8189 83517
rect 8131 83476 8140 83516
rect 8180 83476 8189 83516
rect 8131 83475 8189 83476
rect 8707 83516 8765 83517
rect 8707 83476 8716 83516
rect 8756 83476 8765 83516
rect 8707 83475 8765 83476
rect 13507 83516 13565 83517
rect 13507 83476 13516 83516
rect 13556 83476 13565 83516
rect 13507 83475 13565 83476
rect 15139 83516 15197 83517
rect 15139 83476 15148 83516
rect 15188 83476 15197 83516
rect 15139 83475 15197 83476
rect 15331 83516 15389 83517
rect 15331 83476 15340 83516
rect 15380 83476 15389 83516
rect 15331 83475 15389 83476
rect 15907 83516 15965 83517
rect 15907 83476 15916 83516
rect 15956 83476 15965 83516
rect 15907 83475 15965 83476
rect 18307 83516 18365 83517
rect 18307 83476 18316 83516
rect 18356 83476 18365 83516
rect 18307 83475 18365 83476
rect 18979 83516 19037 83517
rect 18979 83476 18988 83516
rect 19028 83476 19037 83516
rect 18979 83475 19037 83476
rect 19363 83516 19421 83517
rect 19363 83476 19372 83516
rect 19412 83476 19421 83516
rect 19363 83475 19421 83476
rect 1152 83180 20352 83204
rect 1152 83140 3688 83180
rect 3728 83140 3770 83180
rect 3810 83140 3852 83180
rect 3892 83140 3934 83180
rect 3974 83140 4016 83180
rect 4056 83140 18808 83180
rect 18848 83140 18890 83180
rect 18930 83140 18972 83180
rect 19012 83140 19054 83180
rect 19094 83140 19136 83180
rect 19176 83140 20352 83180
rect 1152 83116 20352 83140
rect 2667 83012 2709 83021
rect 2667 82972 2668 83012
rect 2708 82972 2709 83012
rect 2667 82963 2709 82972
rect 3051 83012 3093 83021
rect 3051 82972 3052 83012
rect 3092 82972 3093 83012
rect 3051 82963 3093 82972
rect 3435 83012 3477 83021
rect 3435 82972 3436 83012
rect 3476 82972 3477 83012
rect 3435 82963 3477 82972
rect 3915 83012 3957 83021
rect 3915 82972 3916 83012
rect 3956 82972 3957 83012
rect 3915 82963 3957 82972
rect 4587 83012 4629 83021
rect 4587 82972 4588 83012
rect 4628 82972 4629 83012
rect 4587 82963 4629 82972
rect 19179 83012 19221 83021
rect 19179 82972 19180 83012
rect 19220 82972 19221 83012
rect 19179 82963 19221 82972
rect 19563 83012 19605 83021
rect 19563 82972 19564 83012
rect 19604 82972 19605 83012
rect 19563 82963 19605 82972
rect 2851 82844 2909 82845
rect 2851 82804 2860 82844
rect 2900 82804 2909 82844
rect 2851 82803 2909 82804
rect 3235 82844 3293 82845
rect 3235 82804 3244 82844
rect 3284 82804 3293 82844
rect 3235 82803 3293 82804
rect 3619 82844 3677 82845
rect 3619 82804 3628 82844
rect 3668 82804 3677 82844
rect 3619 82803 3677 82804
rect 4099 82844 4157 82845
rect 4099 82804 4108 82844
rect 4148 82804 4157 82844
rect 4099 82803 4157 82804
rect 4771 82844 4829 82845
rect 4771 82804 4780 82844
rect 4820 82804 4829 82844
rect 4771 82803 4829 82804
rect 18979 82844 19037 82845
rect 18979 82804 18988 82844
rect 19028 82804 19037 82844
rect 18979 82803 19037 82804
rect 19363 82844 19421 82845
rect 19363 82804 19372 82844
rect 19412 82804 19421 82844
rect 19363 82803 19421 82804
rect 1152 82424 20452 82448
rect 1152 82384 4928 82424
rect 4968 82384 5010 82424
rect 5050 82384 5092 82424
rect 5132 82384 5174 82424
rect 5214 82384 5256 82424
rect 5296 82384 20048 82424
rect 20088 82384 20130 82424
rect 20170 82384 20212 82424
rect 20252 82384 20294 82424
rect 20334 82384 20376 82424
rect 20416 82384 20452 82424
rect 1152 82360 20452 82384
rect 14283 82256 14325 82265
rect 14283 82216 14284 82256
rect 14324 82216 14325 82256
rect 14283 82207 14325 82216
rect 15723 82256 15765 82265
rect 15723 82216 15724 82256
rect 15764 82216 15765 82256
rect 15723 82207 15765 82216
rect 14083 82004 14141 82005
rect 14083 81964 14092 82004
rect 14132 81964 14141 82004
rect 14083 81963 14141 81964
rect 15523 82004 15581 82005
rect 15523 81964 15532 82004
rect 15572 81964 15581 82004
rect 15523 81963 15581 81964
rect 1152 81668 20352 81692
rect 1152 81628 3688 81668
rect 3728 81628 3770 81668
rect 3810 81628 3852 81668
rect 3892 81628 3934 81668
rect 3974 81628 4016 81668
rect 4056 81628 18808 81668
rect 18848 81628 18890 81668
rect 18930 81628 18972 81668
rect 19012 81628 19054 81668
rect 19094 81628 19136 81668
rect 19176 81628 20352 81668
rect 1152 81604 20352 81628
rect 19563 81500 19605 81509
rect 19563 81460 19564 81500
rect 19604 81460 19605 81500
rect 19563 81451 19605 81460
rect 19179 81416 19221 81425
rect 19179 81376 19180 81416
rect 19220 81376 19221 81416
rect 19179 81367 19221 81376
rect 18979 81332 19037 81333
rect 18979 81292 18988 81332
rect 19028 81292 19037 81332
rect 18979 81291 19037 81292
rect 19363 81332 19421 81333
rect 19363 81292 19372 81332
rect 19412 81292 19421 81332
rect 19363 81291 19421 81292
rect 1152 80912 20452 80936
rect 1152 80872 4928 80912
rect 4968 80872 5010 80912
rect 5050 80872 5092 80912
rect 5132 80872 5174 80912
rect 5214 80872 5256 80912
rect 5296 80872 20048 80912
rect 20088 80872 20130 80912
rect 20170 80872 20212 80912
rect 20252 80872 20294 80912
rect 20334 80872 20376 80912
rect 20416 80872 20452 80912
rect 1152 80848 20452 80872
rect 13219 80576 13277 80577
rect 13219 80536 13228 80576
rect 13268 80536 13277 80576
rect 13219 80535 13277 80536
rect 14467 80576 14525 80577
rect 14467 80536 14476 80576
rect 14516 80536 14525 80576
rect 14467 80535 14525 80536
rect 18691 80492 18749 80493
rect 18691 80452 18700 80492
rect 18740 80452 18749 80492
rect 18691 80451 18749 80452
rect 19363 80492 19421 80493
rect 19363 80452 19372 80492
rect 19412 80452 19421 80492
rect 19363 80451 19421 80452
rect 19747 80492 19805 80493
rect 19747 80452 19756 80492
rect 19796 80452 19805 80492
rect 19747 80451 19805 80452
rect 18891 80408 18933 80417
rect 18891 80368 18892 80408
rect 18932 80368 18933 80408
rect 18891 80359 18933 80368
rect 19947 80408 19989 80417
rect 19947 80368 19948 80408
rect 19988 80368 19989 80408
rect 19947 80359 19989 80368
rect 14667 80324 14709 80333
rect 14667 80284 14668 80324
rect 14708 80284 14709 80324
rect 14667 80275 14709 80284
rect 19563 80324 19605 80333
rect 19563 80284 19564 80324
rect 19604 80284 19605 80324
rect 19563 80275 19605 80284
rect 1152 80156 20352 80180
rect 1152 80116 3688 80156
rect 3728 80116 3770 80156
rect 3810 80116 3852 80156
rect 3892 80116 3934 80156
rect 3974 80116 4016 80156
rect 4056 80116 18808 80156
rect 18848 80116 18890 80156
rect 18930 80116 18972 80156
rect 19012 80116 19054 80156
rect 19094 80116 19136 80156
rect 19176 80116 20352 80156
rect 1152 80092 20352 80116
rect 15723 79988 15765 79997
rect 15723 79948 15724 79988
rect 15764 79948 15765 79988
rect 15723 79939 15765 79948
rect 15915 79988 15957 79997
rect 15915 79948 15916 79988
rect 15956 79948 15957 79988
rect 15915 79939 15957 79948
rect 16683 79988 16725 79997
rect 16683 79948 16684 79988
rect 16724 79948 16725 79988
rect 16683 79939 16725 79948
rect 19179 79988 19221 79997
rect 19179 79948 19180 79988
rect 19220 79948 19221 79988
rect 19179 79939 19221 79948
rect 15523 79820 15581 79821
rect 15523 79780 15532 79820
rect 15572 79780 15581 79820
rect 15523 79779 15581 79780
rect 16099 79820 16157 79821
rect 16099 79780 16108 79820
rect 16148 79780 16157 79820
rect 16099 79779 16157 79780
rect 16483 79820 16541 79821
rect 16483 79780 16492 79820
rect 16532 79780 16541 79820
rect 16483 79779 16541 79780
rect 18979 79820 19037 79821
rect 18979 79780 18988 79820
rect 19028 79780 19037 79820
rect 18979 79779 19037 79780
rect 19363 79820 19421 79821
rect 19363 79780 19372 79820
rect 19412 79780 19421 79820
rect 19363 79779 19421 79780
rect 19747 79820 19805 79821
rect 19747 79780 19756 79820
rect 19796 79780 19805 79820
rect 19747 79779 19805 79780
rect 11011 79736 11069 79737
rect 11011 79696 11020 79736
rect 11060 79696 11069 79736
rect 11011 79695 11069 79696
rect 12259 79736 12317 79737
rect 12259 79696 12268 79736
rect 12308 79696 12317 79736
rect 12259 79695 12317 79696
rect 13411 79736 13469 79737
rect 13411 79696 13420 79736
rect 13460 79696 13469 79736
rect 13411 79695 13469 79696
rect 14659 79736 14717 79737
rect 14659 79696 14668 79736
rect 14708 79696 14717 79736
rect 14659 79695 14717 79696
rect 10731 79568 10773 79577
rect 10731 79528 10732 79568
rect 10772 79528 10773 79568
rect 10731 79519 10773 79528
rect 12459 79568 12501 79577
rect 12459 79528 12460 79568
rect 12500 79528 12501 79568
rect 12459 79519 12501 79528
rect 14859 79568 14901 79577
rect 14859 79528 14860 79568
rect 14900 79528 14901 79568
rect 14859 79519 14901 79528
rect 19563 79568 19605 79577
rect 19563 79528 19564 79568
rect 19604 79528 19605 79568
rect 19563 79519 19605 79528
rect 19947 79568 19989 79577
rect 19947 79528 19948 79568
rect 19988 79528 19989 79568
rect 19947 79519 19989 79528
rect 1152 79400 20452 79424
rect 1152 79360 4928 79400
rect 4968 79360 5010 79400
rect 5050 79360 5092 79400
rect 5132 79360 5174 79400
rect 5214 79360 5256 79400
rect 5296 79360 20048 79400
rect 20088 79360 20130 79400
rect 20170 79360 20212 79400
rect 20252 79360 20294 79400
rect 20334 79360 20376 79400
rect 20416 79360 20452 79400
rect 1152 79336 20452 79360
rect 19179 79232 19221 79241
rect 19179 79192 19180 79232
rect 19220 79192 19221 79232
rect 19179 79183 19221 79192
rect 10539 79148 10581 79157
rect 10539 79108 10540 79148
rect 10580 79108 10581 79148
rect 10539 79099 10581 79108
rect 12555 79148 12597 79157
rect 12555 79108 12556 79148
rect 12596 79108 12597 79148
rect 12555 79099 12597 79108
rect 14859 79148 14901 79157
rect 14859 79108 14860 79148
rect 14900 79108 14901 79148
rect 14859 79099 14901 79108
rect 9091 79064 9149 79065
rect 9091 79024 9100 79064
rect 9140 79024 9149 79064
rect 9091 79023 9149 79024
rect 10339 79064 10397 79065
rect 10339 79024 10348 79064
rect 10388 79024 10397 79064
rect 10339 79023 10397 79024
rect 10827 79064 10869 79073
rect 10827 79024 10828 79064
rect 10868 79024 10869 79064
rect 10827 79015 10869 79024
rect 10923 79064 10965 79073
rect 10923 79024 10924 79064
rect 10964 79024 10965 79064
rect 10923 79015 10965 79024
rect 11403 79064 11445 79073
rect 11403 79024 11404 79064
rect 11444 79024 11445 79064
rect 11403 79015 11445 79024
rect 11875 79064 11933 79065
rect 11875 79024 11884 79064
rect 11924 79024 11933 79064
rect 13131 79064 13173 79073
rect 11875 79023 11933 79024
rect 12411 79054 12453 79063
rect 12411 79014 12412 79054
rect 12452 79014 12453 79054
rect 13131 79024 13132 79064
rect 13172 79024 13173 79064
rect 13131 79015 13173 79024
rect 13227 79064 13269 79073
rect 13227 79024 13228 79064
rect 13268 79024 13269 79064
rect 13227 79015 13269 79024
rect 13707 79064 13749 79073
rect 13707 79024 13708 79064
rect 13748 79024 13749 79064
rect 13707 79015 13749 79024
rect 14179 79064 14237 79065
rect 14179 79024 14188 79064
rect 14228 79024 14237 79064
rect 15331 79064 15389 79065
rect 14179 79023 14237 79024
rect 14715 79054 14757 79063
rect 12411 79005 12453 79014
rect 14715 79014 14716 79054
rect 14756 79014 14757 79054
rect 15331 79024 15340 79064
rect 15380 79024 15389 79064
rect 15331 79023 15389 79024
rect 16579 79064 16637 79065
rect 16579 79024 16588 79064
rect 16628 79024 16637 79064
rect 16579 79023 16637 79024
rect 14715 79005 14757 79014
rect 11307 78980 11349 78989
rect 11307 78940 11308 78980
rect 11348 78940 11349 78980
rect 11307 78931 11349 78940
rect 13611 78980 13653 78989
rect 13611 78940 13612 78980
rect 13652 78940 13653 78980
rect 13611 78931 13653 78940
rect 18979 78980 19037 78981
rect 18979 78940 18988 78980
rect 19028 78940 19037 78980
rect 18979 78939 19037 78940
rect 19363 78980 19421 78981
rect 19363 78940 19372 78980
rect 19412 78940 19421 78980
rect 19363 78939 19421 78940
rect 19747 78980 19805 78981
rect 19747 78940 19756 78980
rect 19796 78940 19805 78980
rect 19747 78939 19805 78940
rect 16779 78812 16821 78821
rect 16779 78772 16780 78812
rect 16820 78772 16821 78812
rect 16779 78763 16821 78772
rect 19563 78812 19605 78821
rect 19563 78772 19564 78812
rect 19604 78772 19605 78812
rect 19563 78763 19605 78772
rect 19947 78812 19989 78821
rect 19947 78772 19948 78812
rect 19988 78772 19989 78812
rect 19947 78763 19989 78772
rect 1152 78644 20352 78668
rect 1152 78604 3688 78644
rect 3728 78604 3770 78644
rect 3810 78604 3852 78644
rect 3892 78604 3934 78644
rect 3974 78604 4016 78644
rect 4056 78604 18808 78644
rect 18848 78604 18890 78644
rect 18930 78604 18972 78644
rect 19012 78604 19054 78644
rect 19094 78604 19136 78644
rect 19176 78604 20352 78644
rect 1152 78580 20352 78604
rect 13131 78476 13173 78485
rect 13131 78436 13132 78476
rect 13172 78436 13173 78476
rect 13131 78427 13173 78436
rect 18795 78476 18837 78485
rect 18795 78436 18796 78476
rect 18836 78436 18837 78476
rect 18795 78427 18837 78436
rect 19179 78476 19221 78485
rect 19179 78436 19180 78476
rect 19220 78436 19221 78476
rect 19179 78427 19221 78436
rect 8427 78392 8469 78401
rect 8427 78352 8428 78392
rect 8468 78352 8469 78392
rect 8427 78343 8469 78352
rect 19563 78392 19605 78401
rect 19563 78352 19564 78392
rect 19604 78352 19605 78392
rect 19563 78343 19605 78352
rect 18595 78308 18653 78309
rect 16539 78266 16581 78275
rect 18595 78268 18604 78308
rect 18644 78268 18653 78308
rect 18595 78267 18653 78268
rect 18979 78308 19037 78309
rect 18979 78268 18988 78308
rect 19028 78268 19037 78308
rect 18979 78267 19037 78268
rect 19363 78308 19421 78309
rect 19363 78268 19372 78308
rect 19412 78268 19421 78308
rect 19363 78267 19421 78268
rect 19747 78308 19805 78309
rect 19747 78268 19756 78308
rect 19796 78268 19805 78308
rect 19747 78267 19805 78268
rect 11683 78224 11741 78225
rect 11683 78184 11692 78224
rect 11732 78184 11741 78224
rect 11683 78183 11741 78184
rect 12931 78224 12989 78225
rect 12931 78184 12940 78224
rect 12980 78184 12989 78224
rect 12931 78183 12989 78184
rect 14955 78224 14997 78233
rect 14955 78184 14956 78224
rect 14996 78184 14997 78224
rect 14955 78175 14997 78184
rect 15051 78224 15093 78233
rect 15051 78184 15052 78224
rect 15092 78184 15093 78224
rect 15051 78175 15093 78184
rect 15435 78224 15477 78233
rect 15435 78184 15436 78224
rect 15476 78184 15477 78224
rect 15435 78175 15477 78184
rect 15531 78224 15573 78233
rect 16539 78226 16540 78266
rect 16580 78226 16581 78266
rect 15531 78184 15532 78224
rect 15572 78184 15573 78224
rect 15531 78175 15573 78184
rect 16003 78224 16061 78225
rect 16003 78184 16012 78224
rect 16052 78184 16061 78224
rect 16539 78217 16581 78226
rect 16003 78183 16061 78184
rect 10731 78140 10773 78149
rect 10731 78100 10732 78140
rect 10772 78100 10773 78140
rect 10731 78091 10773 78100
rect 16683 78056 16725 78065
rect 16683 78016 16684 78056
rect 16724 78016 16725 78056
rect 16683 78007 16725 78016
rect 19947 78056 19989 78065
rect 19947 78016 19948 78056
rect 19988 78016 19989 78056
rect 19947 78007 19989 78016
rect 1152 77888 20452 77912
rect 1152 77848 4928 77888
rect 4968 77848 5010 77888
rect 5050 77848 5092 77888
rect 5132 77848 5174 77888
rect 5214 77848 5256 77888
rect 5296 77848 20048 77888
rect 20088 77848 20130 77888
rect 20170 77848 20212 77888
rect 20252 77848 20294 77888
rect 20334 77848 20376 77888
rect 20416 77848 20452 77888
rect 1152 77824 20452 77848
rect 8427 77720 8469 77729
rect 8427 77680 8428 77720
rect 8468 77680 8469 77720
rect 8427 77671 8469 77680
rect 16683 77720 16725 77729
rect 16683 77680 16684 77720
rect 16724 77680 16725 77720
rect 16683 77671 16725 77680
rect 17067 77720 17109 77729
rect 17067 77680 17068 77720
rect 17108 77680 17109 77720
rect 17067 77671 17109 77680
rect 8803 77552 8861 77553
rect 8803 77512 8812 77552
rect 8852 77512 8861 77552
rect 8803 77511 8861 77512
rect 10051 77552 10109 77553
rect 10051 77512 10060 77552
rect 10100 77512 10109 77552
rect 10051 77511 10109 77512
rect 10627 77552 10685 77553
rect 10627 77512 10636 77552
rect 10676 77512 10685 77552
rect 10627 77511 10685 77512
rect 11875 77552 11933 77553
rect 11875 77512 11884 77552
rect 11924 77512 11933 77552
rect 11875 77511 11933 77512
rect 13027 77552 13085 77553
rect 13027 77512 13036 77552
rect 13076 77512 13085 77552
rect 13027 77511 13085 77512
rect 14275 77552 14333 77553
rect 14275 77512 14284 77552
rect 14324 77512 14333 77552
rect 14275 77511 14333 77512
rect 15043 77552 15101 77553
rect 15043 77512 15052 77552
rect 15092 77512 15101 77552
rect 15043 77511 15101 77512
rect 16291 77552 16349 77553
rect 16291 77512 16300 77552
rect 16340 77512 16349 77552
rect 16291 77511 16349 77512
rect 17731 77552 17789 77553
rect 17731 77512 17740 77552
rect 17780 77512 17789 77552
rect 17731 77511 17789 77512
rect 18979 77552 19037 77553
rect 18979 77512 18988 77552
rect 19028 77512 19037 77552
rect 18979 77511 19037 77512
rect 19353 77481 19395 77490
rect 16867 77468 16925 77469
rect 16867 77428 16876 77468
rect 16916 77428 16925 77468
rect 16867 77427 16925 77428
rect 17251 77468 17309 77469
rect 17251 77428 17260 77468
rect 17300 77428 17309 77468
rect 19353 77441 19354 77481
rect 19394 77441 19395 77481
rect 19353 77432 19395 77441
rect 19747 77468 19805 77469
rect 17251 77427 17309 77428
rect 19747 77428 19756 77468
rect 19796 77428 19805 77468
rect 19747 77427 19805 77428
rect 10251 77300 10293 77309
rect 10251 77260 10252 77300
rect 10292 77260 10293 77300
rect 10251 77251 10293 77260
rect 12075 77300 12117 77309
rect 12075 77260 12076 77300
rect 12116 77260 12117 77300
rect 12075 77251 12117 77260
rect 14475 77300 14517 77309
rect 14475 77260 14476 77300
rect 14516 77260 14517 77300
rect 14475 77251 14517 77260
rect 16491 77300 16533 77309
rect 16491 77260 16492 77300
rect 16532 77260 16533 77300
rect 16491 77251 16533 77260
rect 19179 77300 19221 77309
rect 19179 77260 19180 77300
rect 19220 77260 19221 77300
rect 19179 77251 19221 77260
rect 19563 77300 19605 77309
rect 19563 77260 19564 77300
rect 19604 77260 19605 77300
rect 19563 77251 19605 77260
rect 19947 77300 19989 77309
rect 19947 77260 19948 77300
rect 19988 77260 19989 77300
rect 19947 77251 19989 77260
rect 1152 77132 20352 77156
rect 1152 77092 3688 77132
rect 3728 77092 3770 77132
rect 3810 77092 3852 77132
rect 3892 77092 3934 77132
rect 3974 77092 4016 77132
rect 4056 77092 18808 77132
rect 18848 77092 18890 77132
rect 18930 77092 18972 77132
rect 19012 77092 19054 77132
rect 19094 77092 19136 77132
rect 19176 77092 20352 77132
rect 1152 77068 20352 77092
rect 8907 76796 8949 76805
rect 8907 76756 8908 76796
rect 8948 76756 8949 76796
rect 8907 76747 8949 76756
rect 10923 76796 10965 76805
rect 10923 76756 10924 76796
rect 10964 76756 10965 76796
rect 15627 76796 15669 76805
rect 10923 76747 10965 76756
rect 12027 76754 12069 76763
rect 6691 76712 6749 76713
rect 6691 76672 6700 76712
rect 6740 76672 6749 76712
rect 6691 76671 6749 76672
rect 7939 76712 7997 76713
rect 7939 76672 7948 76712
rect 7988 76672 7997 76712
rect 7939 76671 7997 76672
rect 8427 76712 8469 76721
rect 8427 76672 8428 76712
rect 8468 76672 8469 76712
rect 8427 76663 8469 76672
rect 8523 76712 8565 76721
rect 8523 76672 8524 76712
rect 8564 76672 8565 76712
rect 8523 76663 8565 76672
rect 9003 76712 9045 76721
rect 9963 76717 10005 76726
rect 9003 76672 9004 76712
rect 9044 76672 9045 76712
rect 9003 76663 9045 76672
rect 9475 76712 9533 76713
rect 9475 76672 9484 76712
rect 9524 76672 9533 76712
rect 9475 76671 9533 76672
rect 9963 76677 9964 76717
rect 10004 76677 10005 76717
rect 9963 76668 10005 76677
rect 10443 76712 10485 76721
rect 10443 76672 10444 76712
rect 10484 76672 10485 76712
rect 10443 76663 10485 76672
rect 10539 76712 10581 76721
rect 10539 76672 10540 76712
rect 10580 76672 10581 76712
rect 10539 76663 10581 76672
rect 11019 76712 11061 76721
rect 12027 76714 12028 76754
rect 12068 76714 12069 76754
rect 15627 76756 15628 76796
rect 15668 76756 15669 76796
rect 15627 76747 15669 76756
rect 18595 76796 18653 76797
rect 18595 76756 18604 76796
rect 18644 76756 18653 76796
rect 18595 76755 18653 76756
rect 18979 76796 19037 76797
rect 18979 76756 18988 76796
rect 19028 76756 19037 76796
rect 18979 76755 19037 76756
rect 19555 76796 19613 76797
rect 19555 76756 19564 76796
rect 19604 76756 19613 76796
rect 19555 76755 19613 76756
rect 19939 76796 19997 76797
rect 19939 76756 19948 76796
rect 19988 76756 19997 76796
rect 19939 76755 19997 76756
rect 14571 76726 14613 76735
rect 11019 76672 11020 76712
rect 11060 76672 11061 76712
rect 11019 76663 11061 76672
rect 11491 76712 11549 76713
rect 11491 76672 11500 76712
rect 11540 76672 11549 76712
rect 12027 76705 12069 76714
rect 13035 76712 13077 76721
rect 11491 76671 11549 76672
rect 13035 76672 13036 76712
rect 13076 76672 13077 76712
rect 13035 76663 13077 76672
rect 13131 76712 13173 76721
rect 13131 76672 13132 76712
rect 13172 76672 13173 76712
rect 13131 76663 13173 76672
rect 13515 76712 13557 76721
rect 13515 76672 13516 76712
rect 13556 76672 13557 76712
rect 13515 76663 13557 76672
rect 13611 76712 13653 76721
rect 13611 76672 13612 76712
rect 13652 76672 13653 76712
rect 13611 76663 13653 76672
rect 14083 76712 14141 76713
rect 14083 76672 14092 76712
rect 14132 76672 14141 76712
rect 14571 76686 14572 76726
rect 14612 76686 14613 76726
rect 16587 76726 16629 76735
rect 14571 76677 14613 76686
rect 15051 76712 15093 76721
rect 14083 76671 14141 76672
rect 15051 76672 15052 76712
rect 15092 76672 15093 76712
rect 15051 76663 15093 76672
rect 15147 76712 15189 76721
rect 15147 76672 15148 76712
rect 15188 76672 15189 76712
rect 15147 76663 15189 76672
rect 15531 76712 15573 76721
rect 15531 76672 15532 76712
rect 15572 76672 15573 76712
rect 15531 76663 15573 76672
rect 16099 76712 16157 76713
rect 16099 76672 16108 76712
rect 16148 76672 16157 76712
rect 16587 76686 16588 76726
rect 16628 76686 16629 76726
rect 16587 76677 16629 76686
rect 17155 76712 17213 76713
rect 16099 76671 16157 76672
rect 17155 76672 17164 76712
rect 17204 76672 17213 76712
rect 17155 76671 17213 76672
rect 18403 76712 18461 76713
rect 18403 76672 18412 76712
rect 18452 76672 18461 76712
rect 18403 76671 18461 76672
rect 8139 76628 8181 76637
rect 8139 76588 8140 76628
rect 8180 76588 8181 76628
rect 8139 76579 8181 76588
rect 10155 76544 10197 76553
rect 10155 76504 10156 76544
rect 10196 76504 10197 76544
rect 10155 76495 10197 76504
rect 12171 76544 12213 76553
rect 12171 76504 12172 76544
rect 12212 76504 12213 76544
rect 12171 76495 12213 76504
rect 14763 76544 14805 76553
rect 14763 76504 14764 76544
rect 14804 76504 14805 76544
rect 14763 76495 14805 76504
rect 16779 76544 16821 76553
rect 16779 76504 16780 76544
rect 16820 76504 16821 76544
rect 16779 76495 16821 76504
rect 16971 76544 17013 76553
rect 16971 76504 16972 76544
rect 17012 76504 17013 76544
rect 16971 76495 17013 76504
rect 18795 76544 18837 76553
rect 18795 76504 18796 76544
rect 18836 76504 18837 76544
rect 18795 76495 18837 76504
rect 19179 76544 19221 76553
rect 19179 76504 19180 76544
rect 19220 76504 19221 76544
rect 19179 76495 19221 76504
rect 19755 76544 19797 76553
rect 19755 76504 19756 76544
rect 19796 76504 19797 76544
rect 19755 76495 19797 76504
rect 20139 76544 20181 76553
rect 20139 76504 20140 76544
rect 20180 76504 20181 76544
rect 20139 76495 20181 76504
rect 1152 76376 20452 76400
rect 1152 76336 4928 76376
rect 4968 76336 5010 76376
rect 5050 76336 5092 76376
rect 5132 76336 5174 76376
rect 5214 76336 5256 76376
rect 5296 76336 20048 76376
rect 20088 76336 20130 76376
rect 20170 76336 20212 76376
rect 20252 76336 20294 76376
rect 20334 76336 20376 76376
rect 20416 76336 20452 76376
rect 1152 76312 20452 76336
rect 8427 76208 8469 76217
rect 8427 76168 8428 76208
rect 8468 76168 8469 76208
rect 8427 76159 8469 76168
rect 10155 76208 10197 76217
rect 10155 76168 10156 76208
rect 10196 76168 10197 76208
rect 10155 76159 10197 76168
rect 14763 76208 14805 76217
rect 14763 76168 14764 76208
rect 14804 76168 14805 76208
rect 14763 76159 14805 76168
rect 15435 76208 15477 76217
rect 15435 76168 15436 76208
rect 15476 76168 15477 76208
rect 15435 76159 15477 76168
rect 19371 76124 19413 76133
rect 19371 76084 19372 76124
rect 19412 76084 19413 76124
rect 19371 76075 19413 76084
rect 6691 76040 6749 76041
rect 6691 76000 6700 76040
rect 6740 76000 6749 76040
rect 6691 75999 6749 76000
rect 7939 76040 7997 76041
rect 7939 76000 7948 76040
rect 7988 76000 7997 76040
rect 7939 75999 7997 76000
rect 8707 76040 8765 76041
rect 8707 76000 8716 76040
rect 8756 76000 8765 76040
rect 8707 75999 8765 76000
rect 9955 76040 10013 76041
rect 9955 76000 9964 76040
rect 10004 76000 10013 76040
rect 9955 75999 10013 76000
rect 11491 76040 11549 76041
rect 11491 76000 11500 76040
rect 11540 76000 11549 76040
rect 11491 75999 11549 76000
rect 12739 76040 12797 76041
rect 12739 76000 12748 76040
rect 12788 76000 12797 76040
rect 12739 75999 12797 76000
rect 13315 76040 13373 76041
rect 13315 76000 13324 76040
rect 13364 76000 13373 76040
rect 13315 75999 13373 76000
rect 14563 76040 14621 76041
rect 14563 76000 14572 76040
rect 14612 76000 14621 76040
rect 14563 75999 14621 76000
rect 15619 76040 15677 76041
rect 15619 76000 15628 76040
rect 15668 76000 15677 76040
rect 15619 75999 15677 76000
rect 16867 76040 16925 76041
rect 16867 76000 16876 76040
rect 16916 76000 16925 76040
rect 16867 75999 16925 76000
rect 17643 76040 17685 76049
rect 17643 76000 17644 76040
rect 17684 76000 17685 76040
rect 17643 75991 17685 76000
rect 17739 76040 17781 76049
rect 17739 76000 17740 76040
rect 17780 76000 17781 76040
rect 17739 75991 17781 76000
rect 18219 76040 18261 76049
rect 18219 76000 18220 76040
rect 18260 76000 18261 76040
rect 18219 75991 18261 76000
rect 18691 76040 18749 76041
rect 18691 76000 18700 76040
rect 18740 76000 18749 76040
rect 18691 75999 18749 76000
rect 19227 76030 19269 76039
rect 19227 75990 19228 76030
rect 19268 75990 19269 76030
rect 19227 75981 19269 75990
rect 15235 75956 15293 75957
rect 15235 75916 15244 75956
rect 15284 75916 15293 75956
rect 15235 75915 15293 75916
rect 18123 75956 18165 75965
rect 18123 75916 18124 75956
rect 18164 75916 18165 75956
rect 18123 75907 18165 75916
rect 19555 75956 19613 75957
rect 19555 75916 19564 75956
rect 19604 75916 19613 75956
rect 19555 75915 19613 75916
rect 19939 75956 19997 75957
rect 19939 75916 19948 75956
rect 19988 75916 19997 75956
rect 19939 75915 19997 75916
rect 10347 75872 10389 75881
rect 10347 75832 10348 75872
rect 10388 75832 10389 75872
rect 10347 75823 10389 75832
rect 12939 75872 12981 75881
rect 12939 75832 12940 75872
rect 12980 75832 12981 75872
rect 12939 75823 12981 75832
rect 17259 75872 17301 75881
rect 17259 75832 17260 75872
rect 17300 75832 17301 75872
rect 17259 75823 17301 75832
rect 8139 75788 8181 75797
rect 8139 75748 8140 75788
rect 8180 75748 8181 75788
rect 8139 75739 8181 75748
rect 17067 75788 17109 75797
rect 17067 75748 17068 75788
rect 17108 75748 17109 75788
rect 17067 75739 17109 75748
rect 19755 75788 19797 75797
rect 19755 75748 19756 75788
rect 19796 75748 19797 75788
rect 19755 75739 19797 75748
rect 20139 75788 20181 75797
rect 20139 75748 20140 75788
rect 20180 75748 20181 75788
rect 20139 75739 20181 75748
rect 1152 75620 20352 75644
rect 1152 75580 3688 75620
rect 3728 75580 3770 75620
rect 3810 75580 3852 75620
rect 3892 75580 3934 75620
rect 3974 75580 4016 75620
rect 4056 75580 18808 75620
rect 18848 75580 18890 75620
rect 18930 75580 18972 75620
rect 19012 75580 19054 75620
rect 19094 75580 19136 75620
rect 19176 75580 20352 75620
rect 1152 75556 20352 75580
rect 8427 75368 8469 75377
rect 8427 75328 8428 75368
rect 8468 75328 8469 75368
rect 8427 75319 8469 75328
rect 18211 75242 18269 75243
rect 18211 75202 18220 75242
rect 18260 75202 18269 75242
rect 18211 75201 18269 75202
rect 6691 75200 6749 75201
rect 6691 75160 6700 75200
rect 6740 75160 6749 75200
rect 6691 75159 6749 75160
rect 7939 75200 7997 75201
rect 7939 75160 7948 75200
rect 7988 75160 7997 75200
rect 7939 75159 7997 75160
rect 9187 75200 9245 75201
rect 9187 75160 9196 75200
rect 9236 75160 9245 75200
rect 9187 75159 9245 75160
rect 10435 75200 10493 75201
rect 10435 75160 10444 75200
rect 10484 75160 10493 75200
rect 10435 75159 10493 75160
rect 10819 75200 10877 75201
rect 10819 75160 10828 75200
rect 10868 75160 10877 75200
rect 10819 75159 10877 75160
rect 12067 75200 12125 75201
rect 12067 75160 12076 75200
rect 12116 75160 12125 75200
rect 12067 75159 12125 75160
rect 13027 75200 13085 75201
rect 13027 75160 13036 75200
rect 13076 75160 13085 75200
rect 13027 75159 13085 75160
rect 14275 75200 14333 75201
rect 14275 75160 14284 75200
rect 14324 75160 14333 75200
rect 14275 75159 14333 75160
rect 15331 75200 15389 75201
rect 15331 75160 15340 75200
rect 15380 75160 15389 75200
rect 15331 75159 15389 75160
rect 16579 75200 16637 75201
rect 16579 75160 16588 75200
rect 16628 75160 16637 75200
rect 16579 75159 16637 75160
rect 16963 75200 17021 75201
rect 16963 75160 16972 75200
rect 17012 75160 17021 75200
rect 16963 75159 17021 75160
rect 18787 75200 18845 75201
rect 18787 75160 18796 75200
rect 18836 75160 18845 75200
rect 18787 75159 18845 75160
rect 20035 75200 20093 75201
rect 20035 75160 20044 75200
rect 20084 75160 20093 75200
rect 20035 75159 20093 75160
rect 8139 75032 8181 75041
rect 8139 74992 8140 75032
rect 8180 74992 8181 75032
rect 8139 74983 8181 74992
rect 8323 75032 8381 75033
rect 8323 74992 8332 75032
rect 8372 74992 8381 75032
rect 8323 74991 8381 74992
rect 10635 75032 10677 75041
rect 10635 74992 10636 75032
rect 10676 74992 10677 75032
rect 10635 74983 10677 74992
rect 12267 75032 12309 75041
rect 12267 74992 12268 75032
rect 12308 74992 12309 75032
rect 12267 74983 12309 74992
rect 14475 75032 14517 75041
rect 14475 74992 14476 75032
rect 14516 74992 14517 75032
rect 14475 74983 14517 74992
rect 16779 75032 16821 75041
rect 16779 74992 16780 75032
rect 16820 74992 16821 75032
rect 16779 74983 16821 74992
rect 18411 75032 18453 75041
rect 18411 74992 18412 75032
rect 18452 74992 18453 75032
rect 18411 74983 18453 74992
rect 18603 75032 18645 75041
rect 18603 74992 18604 75032
rect 18644 74992 18645 75032
rect 18603 74983 18645 74992
rect 1152 74864 20452 74888
rect 1152 74824 4928 74864
rect 4968 74824 5010 74864
rect 5050 74824 5092 74864
rect 5132 74824 5174 74864
rect 5214 74824 5256 74864
rect 5296 74824 20048 74864
rect 20088 74824 20130 74864
rect 20170 74824 20212 74864
rect 20252 74824 20294 74864
rect 20334 74824 20376 74864
rect 20416 74824 20452 74864
rect 1152 74800 20452 74824
rect 10251 74696 10293 74705
rect 10251 74656 10252 74696
rect 10292 74656 10293 74696
rect 10251 74647 10293 74656
rect 14379 74612 14421 74621
rect 14379 74572 14380 74612
rect 14420 74572 14421 74612
rect 14379 74563 14421 74572
rect 16971 74612 17013 74621
rect 16971 74572 16972 74612
rect 17012 74572 17013 74612
rect 16971 74563 17013 74572
rect 19275 74612 19317 74621
rect 19275 74572 19276 74612
rect 19316 74572 19317 74612
rect 19275 74563 19317 74572
rect 5155 74528 5213 74529
rect 5155 74488 5164 74528
rect 5204 74488 5213 74528
rect 5155 74487 5213 74488
rect 6403 74528 6461 74529
rect 6403 74488 6412 74528
rect 6452 74488 6461 74528
rect 6403 74487 6461 74488
rect 6787 74528 6845 74529
rect 6787 74488 6796 74528
rect 6836 74488 6845 74528
rect 6787 74487 6845 74488
rect 8035 74528 8093 74529
rect 8035 74488 8044 74528
rect 8084 74488 8093 74528
rect 8035 74487 8093 74488
rect 8523 74528 8565 74537
rect 8523 74488 8524 74528
rect 8564 74488 8565 74528
rect 8523 74479 8565 74488
rect 8619 74528 8661 74537
rect 8619 74488 8620 74528
rect 8660 74488 8661 74528
rect 8619 74479 8661 74488
rect 9003 74528 9045 74537
rect 9003 74488 9004 74528
rect 9044 74488 9045 74528
rect 9003 74479 9045 74488
rect 9571 74528 9629 74529
rect 9571 74488 9580 74528
rect 9620 74488 9629 74528
rect 9571 74487 9629 74488
rect 10059 74523 10101 74532
rect 10059 74483 10060 74523
rect 10100 74483 10101 74523
rect 10915 74528 10973 74529
rect 10915 74488 10924 74528
rect 10964 74488 10973 74528
rect 10915 74487 10973 74488
rect 12163 74528 12221 74529
rect 12163 74488 12172 74528
rect 12212 74488 12221 74528
rect 12163 74487 12221 74488
rect 12651 74528 12693 74537
rect 12651 74488 12652 74528
rect 12692 74488 12693 74528
rect 10059 74474 10101 74483
rect 12651 74479 12693 74488
rect 12747 74528 12789 74537
rect 12747 74488 12748 74528
rect 12788 74488 12789 74528
rect 12747 74479 12789 74488
rect 13699 74528 13757 74529
rect 13699 74488 13708 74528
rect 13748 74488 13757 74528
rect 15243 74528 15285 74537
rect 13699 74487 13757 74488
rect 14235 74518 14277 74527
rect 14235 74478 14236 74518
rect 14276 74478 14277 74518
rect 15243 74488 15244 74528
rect 15284 74488 15285 74528
rect 15243 74479 15285 74488
rect 15339 74528 15381 74537
rect 15339 74488 15340 74528
rect 15380 74488 15381 74528
rect 15339 74479 15381 74488
rect 15723 74528 15765 74537
rect 15723 74488 15724 74528
rect 15764 74488 15765 74528
rect 15723 74479 15765 74488
rect 16291 74528 16349 74529
rect 16291 74488 16300 74528
rect 16340 74488 16349 74528
rect 16291 74487 16349 74488
rect 16779 74523 16821 74532
rect 16779 74483 16780 74523
rect 16820 74483 16821 74523
rect 14235 74469 14277 74478
rect 16779 74474 16821 74483
rect 17547 74528 17589 74537
rect 17547 74488 17548 74528
rect 17588 74488 17589 74528
rect 17547 74479 17589 74488
rect 17643 74528 17685 74537
rect 17643 74488 17644 74528
rect 17684 74488 17685 74528
rect 17643 74479 17685 74488
rect 18027 74528 18069 74537
rect 18027 74488 18028 74528
rect 18068 74488 18069 74528
rect 18027 74479 18069 74488
rect 18595 74528 18653 74529
rect 18595 74488 18604 74528
rect 18644 74488 18653 74528
rect 18595 74487 18653 74488
rect 19083 74523 19125 74532
rect 19083 74483 19084 74523
rect 19124 74483 19125 74523
rect 19083 74474 19125 74483
rect 19449 74457 19491 74466
rect 9099 74444 9141 74453
rect 9099 74404 9100 74444
rect 9140 74404 9141 74444
rect 9099 74395 9141 74404
rect 13131 74444 13173 74453
rect 13131 74404 13132 74444
rect 13172 74404 13173 74444
rect 13131 74395 13173 74404
rect 13227 74444 13269 74453
rect 13227 74404 13228 74444
rect 13268 74404 13269 74444
rect 13227 74395 13269 74404
rect 15819 74444 15861 74453
rect 15819 74404 15820 74444
rect 15860 74404 15861 74444
rect 15819 74395 15861 74404
rect 18123 74444 18165 74453
rect 18123 74404 18124 74444
rect 18164 74404 18165 74444
rect 19449 74417 19450 74457
rect 19490 74417 19491 74457
rect 19449 74408 19491 74417
rect 19843 74444 19901 74445
rect 18123 74395 18165 74404
rect 19843 74404 19852 74444
rect 19892 74404 19901 74444
rect 19843 74403 19901 74404
rect 6603 74276 6645 74285
rect 6603 74236 6604 74276
rect 6644 74236 6645 74276
rect 6603 74227 6645 74236
rect 8235 74276 8277 74285
rect 8235 74236 8236 74276
rect 8276 74236 8277 74276
rect 8235 74227 8277 74236
rect 12363 74276 12405 74285
rect 12363 74236 12364 74276
rect 12404 74236 12405 74276
rect 12363 74227 12405 74236
rect 19659 74276 19701 74285
rect 19659 74236 19660 74276
rect 19700 74236 19701 74276
rect 19659 74227 19701 74236
rect 20043 74276 20085 74285
rect 20043 74236 20044 74276
rect 20084 74236 20085 74276
rect 20043 74227 20085 74236
rect 1152 74108 20352 74132
rect 1152 74068 3688 74108
rect 3728 74068 3770 74108
rect 3810 74068 3852 74108
rect 3892 74068 3934 74108
rect 3974 74068 4016 74108
rect 4056 74068 18808 74108
rect 18848 74068 18890 74108
rect 18930 74068 18972 74108
rect 19012 74068 19054 74108
rect 19094 74068 19136 74108
rect 19176 74068 20352 74108
rect 1152 74044 20352 74068
rect 14859 73940 14901 73949
rect 14859 73900 14860 73940
rect 14900 73900 14901 73940
rect 14859 73891 14901 73900
rect 19947 73940 19989 73949
rect 19947 73900 19948 73940
rect 19988 73900 19989 73940
rect 19947 73891 19989 73900
rect 5931 73772 5973 73781
rect 5931 73732 5932 73772
rect 5972 73732 5973 73772
rect 5931 73723 5973 73732
rect 9003 73772 9045 73781
rect 9003 73732 9004 73772
rect 9044 73732 9045 73772
rect 9003 73723 9045 73732
rect 11883 73772 11925 73781
rect 11883 73732 11884 73772
rect 11924 73732 11925 73772
rect 11883 73723 11925 73732
rect 11979 73772 12021 73781
rect 11979 73732 11980 73772
rect 12020 73732 12021 73772
rect 11979 73723 12021 73732
rect 18979 73772 19037 73773
rect 18979 73732 18988 73772
rect 19028 73732 19037 73772
rect 18979 73731 19037 73732
rect 19363 73772 19421 73773
rect 19363 73732 19372 73772
rect 19412 73732 19421 73772
rect 19363 73731 19421 73732
rect 19747 73772 19805 73773
rect 19747 73732 19756 73772
rect 19796 73732 19805 73772
rect 19747 73731 19805 73732
rect 6987 73702 7029 73711
rect 12939 73702 12981 73711
rect 3715 73688 3773 73689
rect 3715 73648 3724 73688
rect 3764 73648 3773 73688
rect 3715 73647 3773 73648
rect 4963 73688 5021 73689
rect 4963 73648 4972 73688
rect 5012 73648 5021 73688
rect 4963 73647 5021 73648
rect 5451 73688 5493 73697
rect 5451 73648 5452 73688
rect 5492 73648 5493 73688
rect 5451 73639 5493 73648
rect 5547 73688 5589 73697
rect 5547 73648 5548 73688
rect 5588 73648 5589 73688
rect 5547 73639 5589 73648
rect 6027 73688 6069 73697
rect 6027 73648 6028 73688
rect 6068 73648 6069 73688
rect 6027 73639 6069 73648
rect 6499 73688 6557 73689
rect 6499 73648 6508 73688
rect 6548 73648 6557 73688
rect 6987 73662 6988 73702
rect 7028 73662 7029 73702
rect 6987 73653 7029 73662
rect 8523 73688 8565 73697
rect 6499 73647 6557 73648
rect 8523 73648 8524 73688
rect 8564 73648 8565 73688
rect 8523 73639 8565 73648
rect 8619 73688 8661 73697
rect 8619 73648 8620 73688
rect 8660 73648 8661 73688
rect 8619 73639 8661 73648
rect 9099 73688 9141 73697
rect 10059 73693 10101 73702
rect 9099 73648 9100 73688
rect 9140 73648 9141 73688
rect 9099 73639 9141 73648
rect 9571 73688 9629 73689
rect 9571 73648 9580 73688
rect 9620 73648 9629 73688
rect 9571 73647 9629 73648
rect 10059 73653 10060 73693
rect 10100 73653 10101 73693
rect 10059 73644 10101 73653
rect 11403 73688 11445 73697
rect 11403 73648 11404 73688
rect 11444 73648 11445 73688
rect 11403 73639 11445 73648
rect 11499 73688 11541 73697
rect 11499 73648 11500 73688
rect 11540 73648 11541 73688
rect 11499 73639 11541 73648
rect 12451 73688 12509 73689
rect 12451 73648 12460 73688
rect 12500 73648 12509 73688
rect 12939 73662 12940 73702
rect 12980 73662 12981 73702
rect 16291 73709 16349 73710
rect 12939 73653 12981 73662
rect 13411 73688 13469 73689
rect 12451 73647 12509 73648
rect 13411 73648 13420 73688
rect 13460 73648 13469 73688
rect 13411 73647 13469 73648
rect 14659 73688 14717 73689
rect 14659 73648 14668 73688
rect 14708 73648 14717 73688
rect 14659 73647 14717 73648
rect 15043 73688 15101 73689
rect 15043 73648 15052 73688
rect 15092 73648 15101 73688
rect 16291 73669 16300 73709
rect 16340 73669 16349 73709
rect 16291 73668 16349 73669
rect 17155 73688 17213 73689
rect 15043 73647 15101 73648
rect 17155 73648 17164 73688
rect 17204 73648 17213 73688
rect 17155 73647 17213 73648
rect 18403 73688 18461 73689
rect 18403 73648 18412 73688
rect 18452 73648 18461 73688
rect 18403 73647 18461 73648
rect 5163 73604 5205 73613
rect 5163 73564 5164 73604
rect 5204 73564 5205 73604
rect 5163 73555 5205 73564
rect 13131 73604 13173 73613
rect 13131 73564 13132 73604
rect 13172 73564 13173 73604
rect 13131 73555 13173 73564
rect 7179 73520 7221 73529
rect 7179 73480 7180 73520
rect 7220 73480 7221 73520
rect 7179 73471 7221 73480
rect 10251 73520 10293 73529
rect 10251 73480 10252 73520
rect 10292 73480 10293 73520
rect 10251 73471 10293 73480
rect 16491 73520 16533 73529
rect 16491 73480 16492 73520
rect 16532 73480 16533 73520
rect 16491 73471 16533 73480
rect 18603 73520 18645 73529
rect 18603 73480 18604 73520
rect 18644 73480 18645 73520
rect 18603 73471 18645 73480
rect 19179 73520 19221 73529
rect 19179 73480 19180 73520
rect 19220 73480 19221 73520
rect 19179 73471 19221 73480
rect 19563 73520 19605 73529
rect 19563 73480 19564 73520
rect 19604 73480 19605 73520
rect 19563 73471 19605 73480
rect 1152 73352 20452 73376
rect 1152 73312 4928 73352
rect 4968 73312 5010 73352
rect 5050 73312 5092 73352
rect 5132 73312 5174 73352
rect 5214 73312 5256 73352
rect 5296 73312 20048 73352
rect 20088 73312 20130 73352
rect 20170 73312 20212 73352
rect 20252 73312 20294 73352
rect 20334 73312 20376 73352
rect 20416 73312 20452 73352
rect 1152 73288 20452 73312
rect 18411 73184 18453 73193
rect 18411 73144 18412 73184
rect 18452 73144 18453 73184
rect 18411 73135 18453 73144
rect 8523 73100 8565 73109
rect 8523 73060 8524 73100
rect 8564 73060 8565 73100
rect 8523 73051 8565 73060
rect 13803 73100 13845 73109
rect 13803 73060 13804 73100
rect 13844 73060 13845 73100
rect 13803 73051 13845 73060
rect 3907 73016 3965 73017
rect 3907 72976 3916 73016
rect 3956 72976 3965 73016
rect 3907 72975 3965 72976
rect 5155 73016 5213 73017
rect 5155 72976 5164 73016
rect 5204 72976 5213 73016
rect 5155 72975 5213 72976
rect 7075 73016 7133 73017
rect 7075 72976 7084 73016
rect 7124 72976 7133 73016
rect 7075 72975 7133 72976
rect 8707 73016 8765 73017
rect 8707 72976 8716 73016
rect 8756 72976 8765 73016
rect 8707 72975 8765 72976
rect 9955 73016 10013 73017
rect 9955 72976 9964 73016
rect 10004 72976 10013 73016
rect 9955 72975 10013 72976
rect 10339 73016 10397 73017
rect 10339 72976 10348 73016
rect 10388 72976 10397 73016
rect 10339 72975 10397 72976
rect 11587 73016 11645 73017
rect 11587 72976 11596 73016
rect 11636 72976 11645 73016
rect 11587 72975 11645 72976
rect 12075 73016 12117 73025
rect 12075 72976 12076 73016
rect 12116 72976 12117 73016
rect 8323 72974 8381 72975
rect 8323 72934 8332 72974
rect 8372 72934 8381 72974
rect 12075 72967 12117 72976
rect 12171 73016 12213 73025
rect 12171 72976 12172 73016
rect 12212 72976 12213 73016
rect 12171 72967 12213 72976
rect 13123 73016 13181 73017
rect 13123 72976 13132 73016
rect 13172 72976 13181 73016
rect 14947 73016 15005 73017
rect 13123 72975 13181 72976
rect 13611 73002 13653 73011
rect 13611 72962 13612 73002
rect 13652 72962 13653 73002
rect 14947 72976 14956 73016
rect 14996 72976 15005 73016
rect 14947 72975 15005 72976
rect 16195 73016 16253 73017
rect 16195 72976 16204 73016
rect 16244 72976 16253 73016
rect 16195 72975 16253 72976
rect 16683 73016 16725 73025
rect 16683 72976 16684 73016
rect 16724 72976 16725 73016
rect 16683 72967 16725 72976
rect 16779 73016 16821 73025
rect 16779 72976 16780 73016
rect 16820 72976 16821 73016
rect 16779 72967 16821 72976
rect 17163 73016 17205 73025
rect 17163 72976 17164 73016
rect 17204 72976 17205 73016
rect 17163 72967 17205 72976
rect 17731 73016 17789 73017
rect 17731 72976 17740 73016
rect 17780 72976 17789 73016
rect 17731 72975 17789 72976
rect 18267 73006 18309 73015
rect 13611 72953 13653 72962
rect 18267 72966 18268 73006
rect 18308 72966 18309 73006
rect 18267 72957 18309 72966
rect 8323 72933 8381 72934
rect 12555 72932 12597 72941
rect 12555 72892 12556 72932
rect 12596 72892 12597 72932
rect 12555 72883 12597 72892
rect 12651 72932 12693 72941
rect 12651 72892 12652 72932
rect 12692 72892 12693 72932
rect 12651 72883 12693 72892
rect 17259 72932 17301 72941
rect 17259 72892 17260 72932
rect 17300 72892 17301 72932
rect 17259 72883 17301 72892
rect 18595 72932 18653 72933
rect 18595 72892 18604 72932
rect 18644 72892 18653 72932
rect 18595 72891 18653 72892
rect 18979 72932 19037 72933
rect 18979 72892 18988 72932
rect 19028 72892 19037 72932
rect 18979 72891 19037 72892
rect 19363 72932 19421 72933
rect 19363 72892 19372 72932
rect 19412 72892 19421 72932
rect 19363 72891 19421 72892
rect 19747 72932 19805 72933
rect 19747 72892 19756 72932
rect 19796 72892 19805 72932
rect 19747 72891 19805 72892
rect 10155 72848 10197 72857
rect 10155 72808 10156 72848
rect 10196 72808 10197 72848
rect 10155 72799 10197 72808
rect 18795 72848 18837 72857
rect 18795 72808 18796 72848
rect 18836 72808 18837 72848
rect 18795 72799 18837 72808
rect 19179 72848 19221 72857
rect 19179 72808 19180 72848
rect 19220 72808 19221 72848
rect 19179 72799 19221 72808
rect 5355 72764 5397 72773
rect 5355 72724 5356 72764
rect 5396 72724 5397 72764
rect 5355 72715 5397 72724
rect 11787 72764 11829 72773
rect 11787 72724 11788 72764
rect 11828 72724 11829 72764
rect 11787 72715 11829 72724
rect 16395 72764 16437 72773
rect 16395 72724 16396 72764
rect 16436 72724 16437 72764
rect 16395 72715 16437 72724
rect 19563 72764 19605 72773
rect 19563 72724 19564 72764
rect 19604 72724 19605 72764
rect 19563 72715 19605 72724
rect 19947 72764 19989 72773
rect 19947 72724 19948 72764
rect 19988 72724 19989 72764
rect 19947 72715 19989 72724
rect 1152 72596 20352 72620
rect 1152 72556 3688 72596
rect 3728 72556 3770 72596
rect 3810 72556 3852 72596
rect 3892 72556 3934 72596
rect 3974 72556 4016 72596
rect 4056 72556 18808 72596
rect 18848 72556 18890 72596
rect 18930 72556 18972 72596
rect 19012 72556 19054 72596
rect 19094 72556 19136 72596
rect 19176 72556 20352 72596
rect 1152 72532 20352 72556
rect 19179 72428 19221 72437
rect 19179 72388 19180 72428
rect 19220 72388 19221 72428
rect 19179 72379 19221 72388
rect 18979 72260 19037 72261
rect 17259 72218 17301 72227
rect 1219 72176 1277 72177
rect 1219 72136 1228 72176
rect 1268 72136 1277 72176
rect 1219 72135 1277 72136
rect 2467 72176 2525 72177
rect 2467 72136 2476 72176
rect 2516 72136 2525 72176
rect 2467 72135 2525 72136
rect 4291 72176 4349 72177
rect 4291 72136 4300 72176
rect 4340 72136 4349 72176
rect 4291 72135 4349 72136
rect 5539 72176 5597 72177
rect 5539 72136 5548 72176
rect 5588 72136 5597 72176
rect 5539 72135 5597 72136
rect 5923 72176 5981 72177
rect 5923 72136 5932 72176
rect 5972 72136 5981 72176
rect 5923 72135 5981 72136
rect 7171 72176 7229 72177
rect 7171 72136 7180 72176
rect 7220 72136 7229 72176
rect 7171 72135 7229 72136
rect 7555 72176 7613 72177
rect 7555 72136 7564 72176
rect 7604 72136 7613 72176
rect 7555 72135 7613 72136
rect 8803 72176 8861 72177
rect 8803 72136 8812 72176
rect 8852 72136 8861 72176
rect 8803 72135 8861 72136
rect 10339 72176 10397 72177
rect 10339 72136 10348 72176
rect 10388 72136 10397 72176
rect 10339 72135 10397 72136
rect 11587 72176 11645 72177
rect 11587 72136 11596 72176
rect 11636 72136 11645 72176
rect 11587 72135 11645 72136
rect 11971 72176 12029 72177
rect 11971 72136 11980 72176
rect 12020 72136 12029 72176
rect 11971 72135 12029 72136
rect 13219 72176 13277 72177
rect 13219 72136 13228 72176
rect 13268 72136 13277 72176
rect 13219 72135 13277 72136
rect 13891 72176 13949 72177
rect 13891 72136 13900 72176
rect 13940 72136 13949 72176
rect 13891 72135 13949 72136
rect 15139 72176 15197 72177
rect 15139 72136 15148 72176
rect 15188 72136 15197 72176
rect 15139 72135 15197 72136
rect 16779 72176 16821 72185
rect 16779 72136 16780 72176
rect 16820 72136 16821 72176
rect 17259 72178 17260 72218
rect 17300 72178 17301 72218
rect 17259 72169 17301 72178
rect 17355 72218 17397 72227
rect 18979 72220 18988 72260
rect 19028 72220 19037 72260
rect 18979 72219 19037 72220
rect 19363 72260 19421 72261
rect 19363 72220 19372 72260
rect 19412 72220 19421 72260
rect 19363 72219 19421 72220
rect 19747 72260 19805 72261
rect 19747 72220 19756 72260
rect 19796 72220 19805 72260
rect 19747 72219 19805 72220
rect 17355 72178 17356 72218
rect 17396 72178 17397 72218
rect 17355 72169 17397 72178
rect 18363 72185 18405 72194
rect 17827 72176 17885 72177
rect 16779 72127 16821 72136
rect 16875 72156 16917 72165
rect 16875 72116 16876 72156
rect 16916 72116 16917 72156
rect 17827 72136 17836 72176
rect 17876 72136 17885 72176
rect 18363 72145 18364 72185
rect 18404 72145 18405 72185
rect 18363 72136 18405 72145
rect 17827 72135 17885 72136
rect 16875 72107 16917 72116
rect 2667 72008 2709 72017
rect 2667 71968 2668 72008
rect 2708 71968 2709 72008
rect 2667 71959 2709 71968
rect 5739 72008 5781 72017
rect 5739 71968 5740 72008
rect 5780 71968 5781 72008
rect 5739 71959 5781 71968
rect 7371 72008 7413 72017
rect 7371 71968 7372 72008
rect 7412 71968 7413 72008
rect 7371 71959 7413 71968
rect 9003 72008 9045 72017
rect 9003 71968 9004 72008
rect 9044 71968 9045 72008
rect 9003 71959 9045 71968
rect 11787 72008 11829 72017
rect 11787 71968 11788 72008
rect 11828 71968 11829 72008
rect 11787 71959 11829 71968
rect 13419 72008 13461 72017
rect 13419 71968 13420 72008
rect 13460 71968 13461 72008
rect 13419 71959 13461 71968
rect 15339 72008 15381 72017
rect 15339 71968 15340 72008
rect 15380 71968 15381 72008
rect 15339 71959 15381 71968
rect 18507 72008 18549 72017
rect 18507 71968 18508 72008
rect 18548 71968 18549 72008
rect 18507 71959 18549 71968
rect 19563 72008 19605 72017
rect 19563 71968 19564 72008
rect 19604 71968 19605 72008
rect 19563 71959 19605 71968
rect 19947 72008 19989 72017
rect 19947 71968 19948 72008
rect 19988 71968 19989 72008
rect 19947 71959 19989 71968
rect 1152 71840 20452 71864
rect 1152 71800 4928 71840
rect 4968 71800 5010 71840
rect 5050 71800 5092 71840
rect 5132 71800 5174 71840
rect 5214 71800 5256 71840
rect 5296 71800 20048 71840
rect 20088 71800 20130 71840
rect 20170 71800 20212 71840
rect 20252 71800 20294 71840
rect 20334 71800 20376 71840
rect 20416 71800 20452 71840
rect 1152 71776 20452 71800
rect 8331 71672 8373 71681
rect 8331 71632 8332 71672
rect 8372 71632 8373 71672
rect 8331 71623 8373 71632
rect 15723 71672 15765 71681
rect 15723 71632 15724 71672
rect 15764 71632 15765 71672
rect 15723 71623 15765 71632
rect 6315 71588 6357 71597
rect 6315 71548 6316 71588
rect 6356 71548 6357 71588
rect 6315 71539 6357 71548
rect 10731 71588 10773 71597
rect 10731 71548 10732 71588
rect 10772 71548 10773 71588
rect 10731 71539 10773 71548
rect 13707 71588 13749 71597
rect 13707 71548 13708 71588
rect 13748 71548 13749 71588
rect 13707 71539 13749 71548
rect 1507 71504 1565 71505
rect 1507 71464 1516 71504
rect 1556 71464 1565 71504
rect 1507 71463 1565 71464
rect 2755 71504 2813 71505
rect 2755 71464 2764 71504
rect 2804 71464 2813 71504
rect 2755 71463 2813 71464
rect 4587 71504 4629 71513
rect 4587 71464 4588 71504
rect 4628 71464 4629 71504
rect 4587 71455 4629 71464
rect 4683 71504 4725 71513
rect 4683 71464 4684 71504
rect 4724 71464 4725 71504
rect 4683 71455 4725 71464
rect 5067 71504 5109 71513
rect 5067 71464 5068 71504
rect 5108 71464 5109 71504
rect 5067 71455 5109 71464
rect 5635 71504 5693 71505
rect 5635 71464 5644 71504
rect 5684 71464 5693 71504
rect 6603 71504 6645 71513
rect 5635 71463 5693 71464
rect 6123 71490 6165 71499
rect 6123 71450 6124 71490
rect 6164 71450 6165 71490
rect 6603 71464 6604 71504
rect 6644 71464 6645 71504
rect 6603 71455 6645 71464
rect 6699 71504 6741 71513
rect 6699 71464 6700 71504
rect 6740 71464 6741 71504
rect 6699 71455 6741 71464
rect 7651 71504 7709 71505
rect 7651 71464 7660 71504
rect 7700 71464 7709 71504
rect 7651 71463 7709 71464
rect 8139 71499 8181 71508
rect 8139 71459 8140 71499
rect 8180 71459 8181 71499
rect 8139 71450 8181 71459
rect 9003 71504 9045 71513
rect 9003 71464 9004 71504
rect 9044 71464 9045 71504
rect 9003 71455 9045 71464
rect 9099 71504 9141 71513
rect 9099 71464 9100 71504
rect 9140 71464 9141 71504
rect 9099 71455 9141 71464
rect 10051 71504 10109 71505
rect 10051 71464 10060 71504
rect 10100 71464 10109 71504
rect 11979 71504 12021 71513
rect 10051 71463 10109 71464
rect 10539 71490 10581 71499
rect 10539 71450 10540 71490
rect 10580 71450 10581 71490
rect 11979 71464 11980 71504
rect 12020 71464 12021 71504
rect 11979 71455 12021 71464
rect 12075 71504 12117 71513
rect 12075 71464 12076 71504
rect 12116 71464 12117 71504
rect 12075 71455 12117 71464
rect 13027 71504 13085 71505
rect 13027 71464 13036 71504
rect 13076 71464 13085 71504
rect 13995 71504 14037 71513
rect 13027 71463 13085 71464
rect 13515 71490 13557 71499
rect 6123 71441 6165 71450
rect 10539 71441 10581 71450
rect 13515 71450 13516 71490
rect 13556 71450 13557 71490
rect 13995 71464 13996 71504
rect 14036 71464 14037 71504
rect 13995 71455 14037 71464
rect 14091 71504 14133 71513
rect 14091 71464 14092 71504
rect 14132 71464 14133 71504
rect 14091 71455 14133 71464
rect 14475 71504 14517 71513
rect 14475 71464 14476 71504
rect 14516 71464 14517 71504
rect 14475 71455 14517 71464
rect 15043 71504 15101 71505
rect 15043 71464 15052 71504
rect 15092 71464 15101 71504
rect 15043 71463 15101 71464
rect 15531 71499 15573 71508
rect 15531 71459 15532 71499
rect 15572 71459 15573 71499
rect 15907 71504 15965 71505
rect 15907 71464 15916 71504
rect 15956 71464 15965 71504
rect 15907 71463 15965 71464
rect 17155 71504 17213 71505
rect 17155 71464 17164 71504
rect 17204 71464 17213 71504
rect 17155 71463 17213 71464
rect 17731 71504 17789 71505
rect 17731 71464 17740 71504
rect 17780 71464 17789 71504
rect 17731 71463 17789 71464
rect 18979 71504 19037 71505
rect 18979 71464 18988 71504
rect 19028 71464 19037 71504
rect 18979 71463 19037 71464
rect 15531 71450 15573 71459
rect 13515 71441 13557 71450
rect 5163 71420 5205 71429
rect 5163 71380 5164 71420
rect 5204 71380 5205 71420
rect 5163 71371 5205 71380
rect 7083 71420 7125 71429
rect 7083 71380 7084 71420
rect 7124 71380 7125 71420
rect 7083 71371 7125 71380
rect 7179 71420 7221 71429
rect 7179 71380 7180 71420
rect 7220 71380 7221 71420
rect 7179 71371 7221 71380
rect 8515 71420 8573 71421
rect 8515 71380 8524 71420
rect 8564 71380 8573 71420
rect 8515 71379 8573 71380
rect 9483 71420 9525 71429
rect 9483 71380 9484 71420
rect 9524 71380 9525 71420
rect 9483 71371 9525 71380
rect 9579 71420 9621 71429
rect 9579 71380 9580 71420
rect 9620 71380 9621 71420
rect 9579 71371 9621 71380
rect 12459 71420 12501 71429
rect 12459 71380 12460 71420
rect 12500 71380 12501 71420
rect 12459 71371 12501 71380
rect 12555 71420 12597 71429
rect 12555 71380 12556 71420
rect 12596 71380 12597 71420
rect 12555 71371 12597 71380
rect 14571 71420 14613 71429
rect 14571 71380 14572 71420
rect 14612 71380 14613 71420
rect 14571 71371 14613 71380
rect 19363 71420 19421 71421
rect 19363 71380 19372 71420
rect 19412 71380 19421 71420
rect 19363 71379 19421 71380
rect 19939 71420 19997 71421
rect 19939 71380 19948 71420
rect 19988 71380 19997 71420
rect 19939 71379 19997 71380
rect 2955 71252 2997 71261
rect 2955 71212 2956 71252
rect 2996 71212 2997 71252
rect 2955 71203 2997 71212
rect 8715 71252 8757 71261
rect 8715 71212 8716 71252
rect 8756 71212 8757 71252
rect 8715 71203 8757 71212
rect 17355 71252 17397 71261
rect 17355 71212 17356 71252
rect 17396 71212 17397 71252
rect 17355 71203 17397 71212
rect 19179 71252 19221 71261
rect 19179 71212 19180 71252
rect 19220 71212 19221 71252
rect 19179 71203 19221 71212
rect 19563 71252 19605 71261
rect 19563 71212 19564 71252
rect 19604 71212 19605 71252
rect 19563 71203 19605 71212
rect 20139 71252 20181 71261
rect 20139 71212 20140 71252
rect 20180 71212 20181 71252
rect 20139 71203 20181 71212
rect 1152 71084 20352 71108
rect 1152 71044 3688 71084
rect 3728 71044 3770 71084
rect 3810 71044 3852 71084
rect 3892 71044 3934 71084
rect 3974 71044 4016 71084
rect 4056 71044 18808 71084
rect 18848 71044 18890 71084
rect 18930 71044 18972 71084
rect 19012 71044 19054 71084
rect 19094 71044 19136 71084
rect 19176 71044 20352 71084
rect 1152 71020 20352 71044
rect 5451 70916 5493 70925
rect 5451 70876 5452 70916
rect 5492 70876 5493 70916
rect 5451 70867 5493 70876
rect 8715 70916 8757 70925
rect 8715 70876 8716 70916
rect 8756 70876 8757 70916
rect 8715 70867 8757 70876
rect 13419 70916 13461 70925
rect 13419 70876 13420 70916
rect 13460 70876 13461 70916
rect 13419 70867 13461 70876
rect 19947 70832 19989 70841
rect 19947 70792 19948 70832
rect 19988 70792 19989 70832
rect 19947 70783 19989 70792
rect 9003 70748 9045 70757
rect 9003 70708 9004 70748
rect 9044 70708 9045 70748
rect 9003 70699 9045 70708
rect 19363 70748 19421 70749
rect 19363 70708 19372 70748
rect 19412 70708 19421 70748
rect 19363 70707 19421 70708
rect 19747 70748 19805 70749
rect 19747 70708 19756 70748
rect 19796 70708 19805 70748
rect 19747 70707 19805 70708
rect 2371 70664 2429 70665
rect 2371 70624 2380 70664
rect 2420 70624 2429 70664
rect 2371 70623 2429 70624
rect 3619 70664 3677 70665
rect 3619 70624 3628 70664
rect 3668 70624 3677 70664
rect 3619 70623 3677 70624
rect 4003 70664 4061 70665
rect 4003 70624 4012 70664
rect 4052 70624 4061 70664
rect 4003 70623 4061 70624
rect 5251 70664 5309 70665
rect 5251 70624 5260 70664
rect 5300 70624 5309 70664
rect 5251 70623 5309 70624
rect 5635 70664 5693 70665
rect 5635 70624 5644 70664
rect 5684 70624 5693 70664
rect 5635 70623 5693 70624
rect 6883 70664 6941 70665
rect 6883 70624 6892 70664
rect 6932 70624 6941 70664
rect 6883 70623 6941 70624
rect 7267 70664 7325 70665
rect 7267 70624 7276 70664
rect 7316 70624 7325 70664
rect 7267 70623 7325 70624
rect 8515 70664 8573 70665
rect 8515 70624 8524 70664
rect 8564 70624 8573 70664
rect 8515 70623 8573 70624
rect 10339 70664 10397 70665
rect 10339 70624 10348 70664
rect 10388 70624 10397 70664
rect 10339 70623 10397 70624
rect 11587 70664 11645 70665
rect 11587 70624 11596 70664
rect 11636 70624 11645 70664
rect 11587 70623 11645 70624
rect 11971 70664 12029 70665
rect 11971 70624 11980 70664
rect 12020 70624 12029 70664
rect 11971 70623 12029 70624
rect 13219 70664 13277 70665
rect 13219 70624 13228 70664
rect 13268 70624 13277 70664
rect 13219 70623 13277 70624
rect 13891 70664 13949 70665
rect 13891 70624 13900 70664
rect 13940 70624 13949 70664
rect 13891 70623 13949 70624
rect 15139 70664 15197 70665
rect 15139 70624 15148 70664
rect 15188 70624 15197 70664
rect 15139 70623 15197 70624
rect 16099 70664 16157 70665
rect 16099 70624 16108 70664
rect 16148 70624 16157 70664
rect 16099 70623 16157 70624
rect 17347 70664 17405 70665
rect 17347 70624 17356 70664
rect 17396 70624 17405 70664
rect 17347 70623 17405 70624
rect 17923 70664 17981 70665
rect 17923 70624 17932 70664
rect 17972 70624 17981 70664
rect 17923 70623 17981 70624
rect 19171 70664 19229 70665
rect 19171 70624 19180 70664
rect 19220 70624 19229 70664
rect 19171 70623 19229 70624
rect 17739 70580 17781 70589
rect 17739 70540 17740 70580
rect 17780 70540 17781 70580
rect 17739 70531 17781 70540
rect 3819 70496 3861 70505
rect 3819 70456 3820 70496
rect 3860 70456 3861 70496
rect 3819 70447 3861 70456
rect 7083 70496 7125 70505
rect 7083 70456 7084 70496
rect 7124 70456 7125 70496
rect 7083 70447 7125 70456
rect 11787 70496 11829 70505
rect 11787 70456 11788 70496
rect 11828 70456 11829 70496
rect 11787 70447 11829 70456
rect 15339 70496 15381 70505
rect 15339 70456 15340 70496
rect 15380 70456 15381 70496
rect 15339 70447 15381 70456
rect 17547 70496 17589 70505
rect 17547 70456 17548 70496
rect 17588 70456 17589 70496
rect 17547 70447 17589 70456
rect 19563 70496 19605 70505
rect 19563 70456 19564 70496
rect 19604 70456 19605 70496
rect 19563 70447 19605 70456
rect 1152 70328 20452 70352
rect 1152 70288 4928 70328
rect 4968 70288 5010 70328
rect 5050 70288 5092 70328
rect 5132 70288 5174 70328
rect 5214 70288 5256 70328
rect 5296 70288 20048 70328
rect 20088 70288 20130 70328
rect 20170 70288 20212 70328
rect 20252 70288 20294 70328
rect 20334 70288 20376 70328
rect 20416 70288 20452 70328
rect 1152 70264 20452 70288
rect 11883 70160 11925 70169
rect 11883 70120 11884 70160
rect 11924 70120 11925 70160
rect 11883 70111 11925 70120
rect 17355 70160 17397 70169
rect 17355 70120 17356 70160
rect 17396 70120 17397 70160
rect 17355 70111 17397 70120
rect 9867 70076 9909 70085
rect 9867 70036 9868 70076
rect 9908 70036 9909 70076
rect 4579 70034 4637 70035
rect 4579 69994 4588 70034
rect 4628 69994 4637 70034
rect 9867 70027 9909 70036
rect 19371 70076 19413 70085
rect 19371 70036 19372 70076
rect 19412 70036 19413 70076
rect 19371 70027 19413 70036
rect 4579 69993 4637 69994
rect 1219 69992 1277 69993
rect 1219 69952 1228 69992
rect 1268 69952 1277 69992
rect 1219 69951 1277 69952
rect 2467 69992 2525 69993
rect 2467 69952 2476 69992
rect 2516 69952 2525 69992
rect 2467 69951 2525 69952
rect 2947 69992 3005 69993
rect 2947 69952 2956 69992
rect 2996 69952 3005 69992
rect 2947 69951 3005 69952
rect 4195 69992 4253 69993
rect 4195 69952 4204 69992
rect 4244 69952 4253 69992
rect 4195 69951 4253 69952
rect 5827 69992 5885 69993
rect 5827 69952 5836 69992
rect 5876 69952 5885 69992
rect 5827 69951 5885 69952
rect 6211 69992 6269 69993
rect 6211 69952 6220 69992
rect 6260 69952 6269 69992
rect 6211 69951 6269 69952
rect 7459 69992 7517 69993
rect 7459 69952 7468 69992
rect 7508 69952 7517 69992
rect 7459 69951 7517 69952
rect 8419 69992 8477 69993
rect 8419 69952 8428 69992
rect 8468 69952 8477 69992
rect 8419 69951 8477 69952
rect 9667 69992 9725 69993
rect 9667 69952 9676 69992
rect 9716 69952 9725 69992
rect 9667 69951 9725 69952
rect 10155 69992 10197 70001
rect 10155 69952 10156 69992
rect 10196 69952 10197 69992
rect 10155 69943 10197 69952
rect 10251 69992 10293 70001
rect 10251 69952 10252 69992
rect 10292 69952 10293 69992
rect 10251 69943 10293 69952
rect 11203 69992 11261 69993
rect 11203 69952 11212 69992
rect 11252 69952 11261 69992
rect 13507 69992 13565 69993
rect 11203 69951 11261 69952
rect 11739 69982 11781 69991
rect 11739 69942 11740 69982
rect 11780 69942 11781 69982
rect 13507 69952 13516 69992
rect 13556 69952 13565 69992
rect 13507 69951 13565 69952
rect 14755 69992 14813 69993
rect 14755 69952 14764 69992
rect 14804 69952 14813 69992
rect 14755 69951 14813 69952
rect 15627 69992 15669 70001
rect 15627 69952 15628 69992
rect 15668 69952 15669 69992
rect 15627 69943 15669 69952
rect 15723 69992 15765 70001
rect 15723 69952 15724 69992
rect 15764 69952 15765 69992
rect 15723 69943 15765 69952
rect 16675 69992 16733 69993
rect 16675 69952 16684 69992
rect 16724 69952 16733 69992
rect 16675 69951 16733 69952
rect 17163 69987 17205 69996
rect 17163 69947 17164 69987
rect 17204 69947 17205 69987
rect 11739 69933 11781 69942
rect 17163 69938 17205 69947
rect 17643 69992 17685 70001
rect 17643 69952 17644 69992
rect 17684 69952 17685 69992
rect 17643 69943 17685 69952
rect 17739 69992 17781 70001
rect 17739 69952 17740 69992
rect 17780 69952 17781 69992
rect 17739 69943 17781 69952
rect 18123 69992 18165 70001
rect 18123 69952 18124 69992
rect 18164 69952 18165 69992
rect 18123 69943 18165 69952
rect 18691 69992 18749 69993
rect 18691 69952 18700 69992
rect 18740 69952 18749 69992
rect 18691 69951 18749 69952
rect 19227 69982 19269 69991
rect 19227 69942 19228 69982
rect 19268 69942 19269 69982
rect 19227 69933 19269 69942
rect 10635 69908 10677 69917
rect 10635 69868 10636 69908
rect 10676 69868 10677 69908
rect 10635 69859 10677 69868
rect 10731 69908 10773 69917
rect 10731 69868 10732 69908
rect 10772 69868 10773 69908
rect 10731 69859 10773 69868
rect 16107 69908 16149 69917
rect 16107 69868 16108 69908
rect 16148 69868 16149 69908
rect 16107 69859 16149 69868
rect 16203 69908 16245 69917
rect 16203 69868 16204 69908
rect 16244 69868 16245 69908
rect 16203 69859 16245 69868
rect 18219 69908 18261 69917
rect 18219 69868 18220 69908
rect 18260 69868 18261 69908
rect 18219 69859 18261 69868
rect 19555 69908 19613 69909
rect 19555 69868 19564 69908
rect 19604 69868 19613 69908
rect 19555 69867 19613 69868
rect 19939 69908 19997 69909
rect 19939 69868 19948 69908
rect 19988 69868 19997 69908
rect 19939 69867 19997 69868
rect 2667 69740 2709 69749
rect 2667 69700 2668 69740
rect 2708 69700 2709 69740
rect 2667 69691 2709 69700
rect 4395 69740 4437 69749
rect 4395 69700 4396 69740
rect 4436 69700 4437 69740
rect 4395 69691 4437 69700
rect 6027 69740 6069 69749
rect 6027 69700 6028 69740
rect 6068 69700 6069 69740
rect 6027 69691 6069 69700
rect 7659 69740 7701 69749
rect 7659 69700 7660 69740
rect 7700 69700 7701 69740
rect 7659 69691 7701 69700
rect 14955 69740 14997 69749
rect 14955 69700 14956 69740
rect 14996 69700 14997 69740
rect 14955 69691 14997 69700
rect 19755 69740 19797 69749
rect 19755 69700 19756 69740
rect 19796 69700 19797 69740
rect 19755 69691 19797 69700
rect 20139 69740 20181 69749
rect 20139 69700 20140 69740
rect 20180 69700 20181 69740
rect 20139 69691 20181 69700
rect 1152 69572 20352 69596
rect 1152 69532 3688 69572
rect 3728 69532 3770 69572
rect 3810 69532 3852 69572
rect 3892 69532 3934 69572
rect 3974 69532 4016 69572
rect 4056 69532 18808 69572
rect 18848 69532 18890 69572
rect 18930 69532 18972 69572
rect 19012 69532 19054 69572
rect 19094 69532 19136 69572
rect 19176 69532 20352 69572
rect 1152 69508 20352 69532
rect 11211 69320 11253 69329
rect 11211 69280 11212 69320
rect 11252 69280 11253 69320
rect 11211 69271 11253 69280
rect 17931 69320 17973 69329
rect 17931 69280 17932 69320
rect 17972 69280 17973 69320
rect 17931 69271 17973 69280
rect 17731 69236 17789 69237
rect 17731 69196 17740 69236
rect 17780 69196 17789 69236
rect 17731 69195 17789 69196
rect 19747 69236 19805 69237
rect 19747 69196 19756 69236
rect 19796 69196 19805 69236
rect 19747 69195 19805 69196
rect 16099 69194 16157 69195
rect 4395 69166 4437 69175
rect 2859 69152 2901 69161
rect 2859 69112 2860 69152
rect 2900 69112 2901 69152
rect 2859 69103 2901 69112
rect 2955 69152 2997 69161
rect 2955 69112 2956 69152
rect 2996 69112 2997 69152
rect 2955 69103 2997 69112
rect 3339 69152 3381 69161
rect 3339 69112 3340 69152
rect 3380 69112 3381 69152
rect 3339 69103 3381 69112
rect 3435 69152 3477 69161
rect 3435 69112 3436 69152
rect 3476 69112 3477 69152
rect 3435 69103 3477 69112
rect 3907 69152 3965 69153
rect 3907 69112 3916 69152
rect 3956 69112 3965 69152
rect 4395 69126 4396 69166
rect 4436 69126 4437 69166
rect 6019 69173 6077 69174
rect 4395 69117 4437 69126
rect 4771 69152 4829 69153
rect 3907 69111 3965 69112
rect 4771 69112 4780 69152
rect 4820 69112 4829 69152
rect 6019 69133 6028 69173
rect 6068 69133 6077 69173
rect 8331 69166 8373 69175
rect 6019 69132 6077 69133
rect 6795 69152 6837 69161
rect 4771 69111 4829 69112
rect 6795 69112 6796 69152
rect 6836 69112 6837 69152
rect 6795 69103 6837 69112
rect 6891 69152 6933 69161
rect 6891 69112 6892 69152
rect 6932 69112 6933 69152
rect 6891 69103 6933 69112
rect 7275 69152 7317 69161
rect 7275 69112 7276 69152
rect 7316 69112 7317 69152
rect 7275 69103 7317 69112
rect 7371 69152 7413 69161
rect 7371 69112 7372 69152
rect 7412 69112 7413 69152
rect 7371 69103 7413 69112
rect 7843 69152 7901 69153
rect 7843 69112 7852 69152
rect 7892 69112 7901 69152
rect 8331 69126 8332 69166
rect 8372 69126 8373 69166
rect 15147 69166 15189 69175
rect 8331 69117 8373 69126
rect 8899 69152 8957 69153
rect 7843 69111 7901 69112
rect 8899 69112 8908 69152
rect 8948 69112 8957 69152
rect 8899 69111 8957 69112
rect 10147 69152 10205 69153
rect 10147 69112 10156 69152
rect 10196 69112 10205 69152
rect 10147 69111 10205 69112
rect 10723 69152 10781 69153
rect 10723 69112 10732 69152
rect 10772 69112 10781 69152
rect 10723 69111 10781 69112
rect 11875 69152 11933 69153
rect 11875 69112 11884 69152
rect 11924 69112 11933 69152
rect 11875 69111 11933 69112
rect 13123 69152 13181 69153
rect 13123 69112 13132 69152
rect 13172 69112 13181 69152
rect 13123 69111 13181 69112
rect 13611 69152 13653 69161
rect 13611 69112 13612 69152
rect 13652 69112 13653 69152
rect 13611 69103 13653 69112
rect 13707 69152 13749 69161
rect 13707 69112 13708 69152
rect 13748 69112 13749 69152
rect 13707 69103 13749 69112
rect 14091 69152 14133 69161
rect 14091 69112 14092 69152
rect 14132 69112 14133 69152
rect 14091 69103 14133 69112
rect 14187 69152 14229 69161
rect 14187 69112 14188 69152
rect 14228 69112 14229 69152
rect 14187 69103 14229 69112
rect 14659 69152 14717 69153
rect 14659 69112 14668 69152
rect 14708 69112 14717 69152
rect 15147 69126 15148 69166
rect 15188 69126 15189 69166
rect 16099 69154 16108 69194
rect 16148 69154 16157 69194
rect 16099 69153 16157 69154
rect 15147 69117 15189 69126
rect 17347 69152 17405 69153
rect 14659 69111 14717 69112
rect 17347 69112 17356 69152
rect 17396 69112 17405 69152
rect 17347 69111 17405 69112
rect 18115 69152 18173 69153
rect 18115 69112 18124 69152
rect 18164 69112 18173 69152
rect 18115 69111 18173 69112
rect 19363 69152 19421 69153
rect 19363 69112 19372 69152
rect 19412 69112 19421 69152
rect 19363 69111 19421 69112
rect 8523 69068 8565 69077
rect 8523 69028 8524 69068
rect 8564 69028 8565 69068
rect 8523 69019 8565 69028
rect 13323 69068 13365 69077
rect 13323 69028 13324 69068
rect 13364 69028 13365 69068
rect 13323 69019 13365 69028
rect 15339 69068 15381 69077
rect 15339 69028 15340 69068
rect 15380 69028 15381 69068
rect 15339 69019 15381 69028
rect 4587 68984 4629 68993
rect 4587 68944 4588 68984
rect 4628 68944 4629 68984
rect 4587 68935 4629 68944
rect 6219 68984 6261 68993
rect 6219 68944 6220 68984
rect 6260 68944 6261 68984
rect 6219 68935 6261 68944
rect 10347 68984 10389 68993
rect 10347 68944 10348 68984
rect 10388 68944 10389 68984
rect 10347 68935 10389 68944
rect 17547 68984 17589 68993
rect 17547 68944 17548 68984
rect 17588 68944 17589 68984
rect 17547 68935 17589 68944
rect 19563 68984 19605 68993
rect 19563 68944 19564 68984
rect 19604 68944 19605 68984
rect 19563 68935 19605 68944
rect 19947 68984 19989 68993
rect 19947 68944 19948 68984
rect 19988 68944 19989 68984
rect 19947 68935 19989 68944
rect 1152 68816 20452 68840
rect 1152 68776 4928 68816
rect 4968 68776 5010 68816
rect 5050 68776 5092 68816
rect 5132 68776 5174 68816
rect 5214 68776 5256 68816
rect 5296 68776 20048 68816
rect 20088 68776 20130 68816
rect 20170 68776 20212 68816
rect 20252 68776 20294 68816
rect 20334 68776 20376 68816
rect 20416 68776 20452 68816
rect 1152 68752 20452 68776
rect 12363 68648 12405 68657
rect 12363 68608 12364 68648
rect 12404 68608 12405 68648
rect 12363 68599 12405 68608
rect 19371 68648 19413 68657
rect 19371 68608 19372 68648
rect 19412 68608 19413 68648
rect 19371 68599 19413 68608
rect 5163 68564 5205 68573
rect 5163 68524 5164 68564
rect 5204 68524 5205 68564
rect 5163 68515 5205 68524
rect 8043 68564 8085 68573
rect 8043 68524 8044 68564
rect 8084 68524 8085 68564
rect 8043 68515 8085 68524
rect 1507 68480 1565 68481
rect 1507 68440 1516 68480
rect 1556 68440 1565 68480
rect 1507 68439 1565 68440
rect 2755 68480 2813 68481
rect 2755 68440 2764 68480
rect 2804 68440 2813 68480
rect 2755 68439 2813 68440
rect 3435 68480 3477 68489
rect 3435 68440 3436 68480
rect 3476 68440 3477 68480
rect 3435 68431 3477 68440
rect 3531 68480 3573 68489
rect 3531 68440 3532 68480
rect 3572 68440 3573 68480
rect 3531 68431 3573 68440
rect 4011 68480 4053 68489
rect 4011 68440 4012 68480
rect 4052 68440 4053 68480
rect 4011 68431 4053 68440
rect 4483 68480 4541 68481
rect 4483 68440 4492 68480
rect 4532 68440 4541 68480
rect 4483 68439 4541 68440
rect 4971 68475 5013 68484
rect 4971 68435 4972 68475
rect 5012 68435 5013 68475
rect 4971 68426 5013 68435
rect 6315 68480 6357 68489
rect 6315 68440 6316 68480
rect 6356 68440 6357 68480
rect 6315 68431 6357 68440
rect 6411 68480 6453 68489
rect 6411 68440 6412 68480
rect 6452 68440 6453 68480
rect 6411 68431 6453 68440
rect 7363 68480 7421 68481
rect 7363 68440 7372 68480
rect 7412 68440 7421 68480
rect 7363 68439 7421 68440
rect 7851 68475 7893 68484
rect 7851 68435 7852 68475
rect 7892 68435 7893 68475
rect 8227 68480 8285 68481
rect 8227 68440 8236 68480
rect 8276 68440 8285 68480
rect 8227 68439 8285 68440
rect 9475 68480 9533 68481
rect 9475 68440 9484 68480
rect 9524 68440 9533 68480
rect 9475 68439 9533 68440
rect 10635 68480 10677 68489
rect 10635 68440 10636 68480
rect 10676 68440 10677 68480
rect 7851 68426 7893 68435
rect 10635 68431 10677 68440
rect 10731 68480 10773 68489
rect 10731 68440 10732 68480
rect 10772 68440 10773 68480
rect 10731 68431 10773 68440
rect 11211 68480 11253 68489
rect 11211 68440 11212 68480
rect 11252 68440 11253 68480
rect 11211 68431 11253 68440
rect 11683 68480 11741 68481
rect 11683 68440 11692 68480
rect 11732 68440 11741 68480
rect 14083 68480 14141 68481
rect 11683 68439 11741 68440
rect 12171 68466 12213 68475
rect 12171 68426 12172 68466
rect 12212 68426 12213 68466
rect 14083 68440 14092 68480
rect 14132 68440 14141 68480
rect 14083 68439 14141 68440
rect 15331 68480 15389 68481
rect 15331 68440 15340 68480
rect 15380 68440 15389 68480
rect 15331 68439 15389 68440
rect 15715 68480 15773 68481
rect 15715 68440 15724 68480
rect 15764 68440 15773 68480
rect 15715 68439 15773 68440
rect 16963 68480 17021 68481
rect 16963 68440 16972 68480
rect 17012 68440 17021 68480
rect 16963 68439 17021 68440
rect 17643 68480 17685 68489
rect 17643 68440 17644 68480
rect 17684 68440 17685 68480
rect 17643 68431 17685 68440
rect 17739 68480 17781 68489
rect 17739 68440 17740 68480
rect 17780 68440 17781 68480
rect 17739 68431 17781 68440
rect 18219 68480 18261 68489
rect 18219 68440 18220 68480
rect 18260 68440 18261 68480
rect 18219 68431 18261 68440
rect 18691 68480 18749 68481
rect 18691 68440 18700 68480
rect 18740 68440 18749 68480
rect 18691 68439 18749 68440
rect 19227 68470 19269 68479
rect 12171 68417 12213 68426
rect 19227 68430 19228 68470
rect 19268 68430 19269 68470
rect 19227 68421 19269 68430
rect 3915 68396 3957 68405
rect 3915 68356 3916 68396
rect 3956 68356 3957 68396
rect 3915 68347 3957 68356
rect 6795 68396 6837 68405
rect 6795 68356 6796 68396
rect 6836 68356 6837 68396
rect 6795 68347 6837 68356
rect 6891 68396 6933 68405
rect 6891 68356 6892 68396
rect 6932 68356 6933 68396
rect 6891 68347 6933 68356
rect 11115 68396 11157 68405
rect 11115 68356 11116 68396
rect 11156 68356 11157 68396
rect 11115 68347 11157 68356
rect 18123 68396 18165 68405
rect 18123 68356 18124 68396
rect 18164 68356 18165 68396
rect 18123 68347 18165 68356
rect 19555 68396 19613 68397
rect 19555 68356 19564 68396
rect 19604 68356 19613 68396
rect 19555 68355 19613 68356
rect 19939 68396 19997 68397
rect 19939 68356 19948 68396
rect 19988 68356 19997 68396
rect 19939 68355 19997 68356
rect 2955 68228 2997 68237
rect 2955 68188 2956 68228
rect 2996 68188 2997 68228
rect 2955 68179 2997 68188
rect 9675 68228 9717 68237
rect 9675 68188 9676 68228
rect 9716 68188 9717 68228
rect 9675 68179 9717 68188
rect 15531 68228 15573 68237
rect 15531 68188 15532 68228
rect 15572 68188 15573 68228
rect 15531 68179 15573 68188
rect 17163 68228 17205 68237
rect 17163 68188 17164 68228
rect 17204 68188 17205 68228
rect 17163 68179 17205 68188
rect 19755 68228 19797 68237
rect 19755 68188 19756 68228
rect 19796 68188 19797 68228
rect 19755 68179 19797 68188
rect 20139 68228 20181 68237
rect 20139 68188 20140 68228
rect 20180 68188 20181 68228
rect 20139 68179 20181 68188
rect 1152 68060 20352 68084
rect 1152 68020 3688 68060
rect 3728 68020 3770 68060
rect 3810 68020 3852 68060
rect 3892 68020 3934 68060
rect 3974 68020 4016 68060
rect 4056 68020 18808 68060
rect 18848 68020 18890 68060
rect 18930 68020 18972 68060
rect 19012 68020 19054 68060
rect 19094 68020 19136 68060
rect 19176 68020 20352 68060
rect 1152 67996 20352 68020
rect 11595 67892 11637 67901
rect 11595 67852 11596 67892
rect 11636 67852 11637 67892
rect 11595 67843 11637 67852
rect 15915 67892 15957 67901
rect 15915 67852 15916 67892
rect 15956 67852 15957 67892
rect 15915 67843 15957 67852
rect 10251 67724 10293 67733
rect 10251 67684 10252 67724
rect 10292 67684 10293 67724
rect 15715 67724 15773 67725
rect 10251 67675 10293 67684
rect 11259 67682 11301 67691
rect 15715 67684 15724 67724
rect 15764 67684 15773 67724
rect 15715 67683 15773 67684
rect 19747 67724 19805 67725
rect 19747 67684 19756 67724
rect 19796 67684 19805 67724
rect 19747 67683 19805 67684
rect 1315 67640 1373 67641
rect 1315 67600 1324 67640
rect 1364 67600 1373 67640
rect 1315 67599 1373 67600
rect 2563 67640 2621 67641
rect 2563 67600 2572 67640
rect 2612 67600 2621 67640
rect 2563 67599 2621 67600
rect 2947 67640 3005 67641
rect 2947 67600 2956 67640
rect 2996 67600 3005 67640
rect 2947 67599 3005 67600
rect 4195 67640 4253 67641
rect 4195 67600 4204 67640
rect 4244 67600 4253 67640
rect 4195 67599 4253 67600
rect 4579 67640 4637 67641
rect 4579 67600 4588 67640
rect 4628 67600 4637 67640
rect 4579 67599 4637 67600
rect 5827 67640 5885 67641
rect 5827 67600 5836 67640
rect 5876 67600 5885 67640
rect 5827 67599 5885 67600
rect 6211 67640 6269 67641
rect 6211 67600 6220 67640
rect 6260 67600 6269 67640
rect 6211 67599 6269 67600
rect 7459 67640 7517 67641
rect 7459 67600 7468 67640
rect 7508 67600 7517 67640
rect 7459 67599 7517 67600
rect 7843 67640 7901 67641
rect 7843 67600 7852 67640
rect 7892 67600 7901 67640
rect 7843 67599 7901 67600
rect 9091 67640 9149 67641
rect 9091 67600 9100 67640
rect 9140 67600 9149 67640
rect 9091 67599 9149 67600
rect 9675 67640 9717 67649
rect 9675 67600 9676 67640
rect 9716 67600 9717 67640
rect 9675 67591 9717 67600
rect 9771 67640 9813 67649
rect 9771 67600 9772 67640
rect 9812 67600 9813 67640
rect 9771 67591 9813 67600
rect 10155 67640 10197 67649
rect 11259 67642 11260 67682
rect 11300 67642 11301 67682
rect 17739 67654 17781 67663
rect 10155 67600 10156 67640
rect 10196 67600 10197 67640
rect 10155 67591 10197 67600
rect 10723 67640 10781 67641
rect 10723 67600 10732 67640
rect 10772 67600 10781 67640
rect 11259 67633 11301 67642
rect 11779 67640 11837 67641
rect 10723 67599 10781 67600
rect 11779 67600 11788 67640
rect 11828 67600 11837 67640
rect 11779 67599 11837 67600
rect 13027 67640 13085 67641
rect 13027 67600 13036 67640
rect 13076 67600 13085 67640
rect 13027 67599 13085 67600
rect 13411 67640 13469 67641
rect 13411 67600 13420 67640
rect 13460 67600 13469 67640
rect 13411 67599 13469 67600
rect 14659 67640 14717 67641
rect 14659 67600 14668 67640
rect 14708 67600 14717 67640
rect 14659 67599 14717 67600
rect 16203 67640 16245 67649
rect 16203 67600 16204 67640
rect 16244 67600 16245 67640
rect 16683 67640 16725 67649
rect 16203 67591 16245 67600
rect 16299 67620 16341 67629
rect 16299 67580 16300 67620
rect 16340 67580 16341 67620
rect 16683 67600 16684 67640
rect 16724 67600 16725 67640
rect 16683 67591 16725 67600
rect 16779 67640 16821 67649
rect 16779 67600 16780 67640
rect 16820 67600 16821 67640
rect 16779 67591 16821 67600
rect 17251 67640 17309 67641
rect 17251 67600 17260 67640
rect 17300 67600 17309 67640
rect 17739 67614 17740 67654
rect 17780 67614 17781 67654
rect 17739 67605 17781 67614
rect 18115 67640 18173 67641
rect 17251 67599 17309 67600
rect 18115 67600 18124 67640
rect 18164 67600 18173 67640
rect 18115 67599 18173 67600
rect 19363 67640 19421 67641
rect 19363 67600 19372 67640
rect 19412 67600 19421 67640
rect 19363 67599 19421 67600
rect 16299 67571 16341 67580
rect 11403 67556 11445 67565
rect 11403 67516 11404 67556
rect 11444 67516 11445 67556
rect 11403 67507 11445 67516
rect 17931 67556 17973 67565
rect 17931 67516 17932 67556
rect 17972 67516 17973 67556
rect 17931 67507 17973 67516
rect 2763 67472 2805 67481
rect 2763 67432 2764 67472
rect 2804 67432 2805 67472
rect 2763 67423 2805 67432
rect 4395 67472 4437 67481
rect 4395 67432 4396 67472
rect 4436 67432 4437 67472
rect 4395 67423 4437 67432
rect 6027 67472 6069 67481
rect 6027 67432 6028 67472
rect 6068 67432 6069 67472
rect 6027 67423 6069 67432
rect 7659 67472 7701 67481
rect 7659 67432 7660 67472
rect 7700 67432 7701 67472
rect 7659 67423 7701 67432
rect 9291 67472 9333 67481
rect 9291 67432 9292 67472
rect 9332 67432 9333 67472
rect 9291 67423 9333 67432
rect 14859 67472 14901 67481
rect 14859 67432 14860 67472
rect 14900 67432 14901 67472
rect 14859 67423 14901 67432
rect 19563 67472 19605 67481
rect 19563 67432 19564 67472
rect 19604 67432 19605 67472
rect 19563 67423 19605 67432
rect 19947 67472 19989 67481
rect 19947 67432 19948 67472
rect 19988 67432 19989 67472
rect 19947 67423 19989 67432
rect 1152 67304 20452 67328
rect 1152 67264 4928 67304
rect 4968 67264 5010 67304
rect 5050 67264 5092 67304
rect 5132 67264 5174 67304
rect 5214 67264 5256 67304
rect 5296 67264 20048 67304
rect 20088 67264 20130 67304
rect 20170 67264 20212 67304
rect 20252 67264 20294 67304
rect 20334 67264 20376 67304
rect 20416 67264 20452 67304
rect 1152 67240 20452 67264
rect 9675 67136 9717 67145
rect 9675 67096 9676 67136
rect 9716 67096 9717 67136
rect 9675 67087 9717 67096
rect 11499 67136 11541 67145
rect 11499 67096 11500 67136
rect 11540 67096 11541 67136
rect 11499 67087 11541 67096
rect 15243 67136 15285 67145
rect 15243 67096 15244 67136
rect 15284 67096 15285 67136
rect 15243 67087 15285 67096
rect 19851 67136 19893 67145
rect 19851 67096 19852 67136
rect 19892 67096 19893 67136
rect 19851 67087 19893 67096
rect 20235 67136 20277 67145
rect 20235 67096 20236 67136
rect 20276 67096 20277 67136
rect 20235 67087 20277 67096
rect 13227 67052 13269 67061
rect 13227 67012 13228 67052
rect 13268 67012 13269 67052
rect 13227 67003 13269 67012
rect 13515 66988 13557 66997
rect 1219 66968 1277 66969
rect 1219 66928 1228 66968
rect 1268 66928 1277 66968
rect 1219 66927 1277 66928
rect 2467 66968 2525 66969
rect 2467 66928 2476 66968
rect 2516 66928 2525 66968
rect 2467 66927 2525 66928
rect 3331 66968 3389 66969
rect 3331 66928 3340 66968
rect 3380 66928 3389 66968
rect 3331 66927 3389 66928
rect 4579 66968 4637 66969
rect 4579 66928 4588 66968
rect 4628 66928 4637 66968
rect 4579 66927 4637 66928
rect 4963 66968 5021 66969
rect 4963 66928 4972 66968
rect 5012 66928 5021 66968
rect 4963 66927 5021 66928
rect 6211 66968 6269 66969
rect 6211 66928 6220 66968
rect 6260 66928 6269 66968
rect 6211 66927 6269 66928
rect 7947 66968 7989 66977
rect 7947 66928 7948 66968
rect 7988 66928 7989 66968
rect 7947 66919 7989 66928
rect 8043 66968 8085 66977
rect 8043 66928 8044 66968
rect 8084 66928 8085 66968
rect 8043 66919 8085 66928
rect 8523 66968 8565 66977
rect 8523 66928 8524 66968
rect 8564 66928 8565 66968
rect 8523 66919 8565 66928
rect 8995 66968 9053 66969
rect 8995 66928 9004 66968
rect 9044 66928 9053 66968
rect 8995 66927 9053 66928
rect 9483 66963 9525 66972
rect 9483 66923 9484 66963
rect 9524 66923 9525 66963
rect 10051 66968 10109 66969
rect 10051 66928 10060 66968
rect 10100 66928 10109 66968
rect 10051 66927 10109 66928
rect 11299 66968 11357 66969
rect 11299 66928 11308 66968
rect 11348 66928 11357 66968
rect 11299 66927 11357 66928
rect 11779 66968 11837 66969
rect 11779 66928 11788 66968
rect 11828 66928 11837 66968
rect 11779 66927 11837 66928
rect 13027 66968 13085 66969
rect 13027 66928 13036 66968
rect 13076 66928 13085 66968
rect 13515 66948 13516 66988
rect 13556 66948 13557 66988
rect 13515 66939 13557 66948
rect 13611 66968 13653 66977
rect 13027 66927 13085 66928
rect 13611 66928 13612 66968
rect 13652 66928 13653 66968
rect 9483 66914 9525 66923
rect 13611 66919 13653 66928
rect 13995 66968 14037 66977
rect 13995 66928 13996 66968
rect 14036 66928 14037 66968
rect 13995 66919 14037 66928
rect 14563 66968 14621 66969
rect 14563 66928 14572 66968
rect 14612 66928 14621 66968
rect 14563 66927 14621 66928
rect 15051 66963 15093 66972
rect 15051 66923 15052 66963
rect 15092 66923 15093 66963
rect 16867 66968 16925 66969
rect 16867 66928 16876 66968
rect 16916 66928 16925 66968
rect 16867 66927 16925 66928
rect 17251 66968 17309 66969
rect 17251 66928 17260 66968
rect 17300 66928 17309 66968
rect 17251 66927 17309 66928
rect 18499 66968 18557 66969
rect 18499 66928 18508 66968
rect 18548 66928 18557 66968
rect 18499 66927 18557 66928
rect 15051 66914 15093 66923
rect 15619 66926 15677 66927
rect 8427 66884 8469 66893
rect 8427 66844 8428 66884
rect 8468 66844 8469 66884
rect 8427 66835 8469 66844
rect 14091 66884 14133 66893
rect 15619 66886 15628 66926
rect 15668 66886 15677 66926
rect 15619 66885 15677 66886
rect 14091 66844 14092 66884
rect 14132 66844 14133 66884
rect 14091 66835 14133 66844
rect 19651 66884 19709 66885
rect 19651 66844 19660 66884
rect 19700 66844 19709 66884
rect 19651 66843 19709 66844
rect 20035 66884 20093 66885
rect 20035 66844 20044 66884
rect 20084 66844 20093 66884
rect 20035 66843 20093 66844
rect 4779 66800 4821 66809
rect 4779 66760 4780 66800
rect 4820 66760 4821 66800
rect 4779 66751 4821 66760
rect 6411 66800 6453 66809
rect 6411 66760 6412 66800
rect 6452 66760 6453 66800
rect 6411 66751 6453 66760
rect 2667 66716 2709 66725
rect 2667 66676 2668 66716
rect 2708 66676 2709 66716
rect 2667 66667 2709 66676
rect 17067 66716 17109 66725
rect 17067 66676 17068 66716
rect 17108 66676 17109 66716
rect 17067 66667 17109 66676
rect 18699 66716 18741 66725
rect 18699 66676 18700 66716
rect 18740 66676 18741 66716
rect 18699 66667 18741 66676
rect 1152 66548 20352 66572
rect 1152 66508 3688 66548
rect 3728 66508 3770 66548
rect 3810 66508 3852 66548
rect 3892 66508 3934 66548
rect 3974 66508 4016 66548
rect 4056 66508 18808 66548
rect 18848 66508 18890 66548
rect 18930 66508 18972 66548
rect 19012 66508 19054 66548
rect 19094 66508 19136 66548
rect 19176 66508 20352 66548
rect 1152 66484 20352 66508
rect 17163 66296 17205 66305
rect 17163 66256 17164 66296
rect 17204 66256 17205 66296
rect 17163 66247 17205 66256
rect 19947 66296 19989 66305
rect 19947 66256 19948 66296
rect 19988 66256 19989 66296
rect 19947 66247 19989 66256
rect 4203 66212 4245 66221
rect 4203 66172 4204 66212
rect 4244 66172 4245 66212
rect 4203 66163 4245 66172
rect 6315 66212 6357 66221
rect 6315 66172 6316 66212
rect 6356 66172 6357 66212
rect 6315 66163 6357 66172
rect 6411 66212 6453 66221
rect 6411 66172 6412 66212
rect 6452 66172 6453 66212
rect 6411 66163 6453 66172
rect 18027 66212 18069 66221
rect 18027 66172 18028 66212
rect 18068 66172 18069 66212
rect 18027 66163 18069 66172
rect 19363 66212 19421 66213
rect 19363 66172 19372 66212
rect 19412 66172 19421 66212
rect 19363 66171 19421 66172
rect 19747 66212 19805 66213
rect 19747 66172 19756 66212
rect 19796 66172 19805 66212
rect 19747 66171 19805 66172
rect 5163 66142 5205 66151
rect 1411 66128 1469 66129
rect 1411 66088 1420 66128
rect 1460 66088 1469 66128
rect 1411 66087 1469 66088
rect 2659 66128 2717 66129
rect 2659 66088 2668 66128
rect 2708 66088 2717 66128
rect 2659 66087 2717 66088
rect 3627 66128 3669 66137
rect 3627 66088 3628 66128
rect 3668 66088 3669 66128
rect 3627 66079 3669 66088
rect 3723 66128 3765 66137
rect 3723 66088 3724 66128
rect 3764 66088 3765 66128
rect 3723 66079 3765 66088
rect 4107 66128 4149 66137
rect 4107 66088 4108 66128
rect 4148 66088 4149 66128
rect 4107 66079 4149 66088
rect 4675 66128 4733 66129
rect 4675 66088 4684 66128
rect 4724 66088 4733 66128
rect 5163 66102 5164 66142
rect 5204 66102 5205 66142
rect 7371 66142 7413 66151
rect 5163 66093 5205 66102
rect 5835 66128 5877 66137
rect 4675 66087 4733 66088
rect 5835 66088 5836 66128
rect 5876 66088 5877 66128
rect 5835 66079 5877 66088
rect 5931 66128 5973 66137
rect 5931 66088 5932 66128
rect 5972 66088 5973 66128
rect 5931 66079 5973 66088
rect 6883 66128 6941 66129
rect 6883 66088 6892 66128
rect 6932 66088 6941 66128
rect 7371 66102 7372 66142
rect 7412 66102 7413 66142
rect 19035 66137 19077 66146
rect 7371 66093 7413 66102
rect 9091 66128 9149 66129
rect 6883 66087 6941 66088
rect 9091 66088 9100 66128
rect 9140 66088 9149 66128
rect 9091 66087 9149 66088
rect 10339 66128 10397 66129
rect 10339 66088 10348 66128
rect 10388 66088 10397 66128
rect 10339 66087 10397 66088
rect 10723 66128 10781 66129
rect 10723 66088 10732 66128
rect 10772 66088 10781 66128
rect 10723 66087 10781 66088
rect 11971 66128 12029 66129
rect 11971 66088 11980 66128
rect 12020 66088 12029 66128
rect 11971 66087 12029 66088
rect 12355 66128 12413 66129
rect 12355 66088 12364 66128
rect 12404 66088 12413 66128
rect 12355 66087 12413 66088
rect 13603 66128 13661 66129
rect 13603 66088 13612 66128
rect 13652 66088 13661 66128
rect 13603 66087 13661 66088
rect 13987 66128 14045 66129
rect 13987 66088 13996 66128
rect 14036 66088 14045 66128
rect 13987 66087 14045 66088
rect 15235 66128 15293 66129
rect 15235 66088 15244 66128
rect 15284 66088 15293 66128
rect 15235 66087 15293 66088
rect 17451 66128 17493 66137
rect 17451 66088 17452 66128
rect 17492 66088 17493 66128
rect 17451 66079 17493 66088
rect 17547 66128 17589 66137
rect 17547 66088 17548 66128
rect 17588 66088 17589 66128
rect 17547 66079 17589 66088
rect 17931 66128 17973 66137
rect 17931 66088 17932 66128
rect 17972 66088 17973 66128
rect 17931 66079 17973 66088
rect 18499 66128 18557 66129
rect 18499 66088 18508 66128
rect 18548 66088 18557 66128
rect 19035 66097 19036 66137
rect 19076 66097 19077 66137
rect 19035 66088 19077 66097
rect 18499 66087 18557 66088
rect 7563 66044 7605 66053
rect 7563 66004 7564 66044
rect 7604 66004 7605 66044
rect 7563 65995 7605 66004
rect 2859 65960 2901 65969
rect 2859 65920 2860 65960
rect 2900 65920 2901 65960
rect 2859 65911 2901 65920
rect 5355 65960 5397 65969
rect 5355 65920 5356 65960
rect 5396 65920 5397 65960
rect 5355 65911 5397 65920
rect 10539 65960 10581 65969
rect 10539 65920 10540 65960
rect 10580 65920 10581 65960
rect 10539 65911 10581 65920
rect 12171 65960 12213 65969
rect 12171 65920 12172 65960
rect 12212 65920 12213 65960
rect 12171 65911 12213 65920
rect 13803 65960 13845 65969
rect 13803 65920 13804 65960
rect 13844 65920 13845 65960
rect 13803 65911 13845 65920
rect 15435 65960 15477 65969
rect 15435 65920 15436 65960
rect 15476 65920 15477 65960
rect 15435 65911 15477 65920
rect 19179 65960 19221 65969
rect 19179 65920 19180 65960
rect 19220 65920 19221 65960
rect 19179 65911 19221 65920
rect 19563 65960 19605 65969
rect 19563 65920 19564 65960
rect 19604 65920 19605 65960
rect 19563 65911 19605 65920
rect 1152 65792 20452 65816
rect 1152 65752 4928 65792
rect 4968 65752 5010 65792
rect 5050 65752 5092 65792
rect 5132 65752 5174 65792
rect 5214 65752 5256 65792
rect 5296 65752 20048 65792
rect 20088 65752 20130 65792
rect 20170 65752 20212 65792
rect 20252 65752 20294 65792
rect 20334 65752 20376 65792
rect 20416 65752 20452 65792
rect 1152 65728 20452 65752
rect 16299 65624 16341 65633
rect 16299 65584 16300 65624
rect 16340 65584 16341 65624
rect 16299 65575 16341 65584
rect 4491 65540 4533 65549
rect 4491 65500 4492 65540
rect 4532 65500 4533 65540
rect 4491 65491 4533 65500
rect 12555 65540 12597 65549
rect 12555 65500 12556 65540
rect 12596 65500 12597 65540
rect 12555 65491 12597 65500
rect 15435 65540 15477 65549
rect 15435 65500 15436 65540
rect 15476 65500 15477 65540
rect 15435 65491 15477 65500
rect 18315 65540 18357 65549
rect 18315 65500 18316 65540
rect 18356 65500 18357 65540
rect 18315 65491 18357 65500
rect 2763 65456 2805 65465
rect 2763 65416 2764 65456
rect 2804 65416 2805 65456
rect 2763 65407 2805 65416
rect 2859 65456 2901 65465
rect 2859 65416 2860 65456
rect 2900 65416 2901 65456
rect 2859 65407 2901 65416
rect 3243 65456 3285 65465
rect 3243 65416 3244 65456
rect 3284 65416 3285 65456
rect 3811 65456 3869 65457
rect 3243 65407 3285 65416
rect 3339 65414 3381 65423
rect 3811 65416 3820 65456
rect 3860 65416 3869 65456
rect 3811 65415 3869 65416
rect 4299 65451 4341 65460
rect 3339 65374 3340 65414
rect 3380 65374 3381 65414
rect 4299 65411 4300 65451
rect 4340 65411 4341 65451
rect 5827 65456 5885 65457
rect 5827 65416 5836 65456
rect 5876 65416 5885 65456
rect 5827 65415 5885 65416
rect 7075 65456 7133 65457
rect 7075 65416 7084 65456
rect 7124 65416 7133 65456
rect 7075 65415 7133 65416
rect 7459 65456 7517 65457
rect 7459 65416 7468 65456
rect 7508 65416 7517 65456
rect 7459 65415 7517 65416
rect 8707 65456 8765 65457
rect 8707 65416 8716 65456
rect 8756 65416 8765 65456
rect 8707 65415 8765 65416
rect 9091 65456 9149 65457
rect 9091 65416 9100 65456
rect 9140 65416 9149 65456
rect 9091 65415 9149 65416
rect 10339 65456 10397 65457
rect 10339 65416 10348 65456
rect 10388 65416 10397 65456
rect 10339 65415 10397 65416
rect 10827 65456 10869 65465
rect 10827 65416 10828 65456
rect 10868 65416 10869 65456
rect 4299 65402 4341 65411
rect 10827 65407 10869 65416
rect 10923 65456 10965 65465
rect 10923 65416 10924 65456
rect 10964 65416 10965 65456
rect 10923 65407 10965 65416
rect 11307 65456 11349 65465
rect 11307 65416 11308 65456
rect 11348 65416 11349 65456
rect 11307 65407 11349 65416
rect 11403 65456 11445 65465
rect 11403 65416 11404 65456
rect 11444 65416 11445 65456
rect 11403 65407 11445 65416
rect 11875 65456 11933 65457
rect 11875 65416 11884 65456
rect 11924 65416 11933 65456
rect 11875 65415 11933 65416
rect 12363 65451 12405 65460
rect 12363 65411 12364 65451
rect 12404 65411 12405 65451
rect 12363 65402 12405 65411
rect 13707 65456 13749 65465
rect 13707 65416 13708 65456
rect 13748 65416 13749 65456
rect 13707 65407 13749 65416
rect 13803 65456 13845 65465
rect 13803 65416 13804 65456
rect 13844 65416 13845 65456
rect 13803 65407 13845 65416
rect 14187 65456 14229 65465
rect 14187 65416 14188 65456
rect 14228 65416 14229 65456
rect 14187 65407 14229 65416
rect 14283 65456 14325 65465
rect 14283 65416 14284 65456
rect 14324 65416 14325 65456
rect 14283 65407 14325 65416
rect 14755 65456 14813 65457
rect 14755 65416 14764 65456
rect 14804 65416 14813 65456
rect 16587 65456 16629 65465
rect 14755 65415 14813 65416
rect 15291 65446 15333 65455
rect 15291 65406 15292 65446
rect 15332 65406 15333 65446
rect 16587 65416 16588 65456
rect 16628 65416 16629 65456
rect 16587 65407 16629 65416
rect 16683 65456 16725 65465
rect 16683 65416 16684 65456
rect 16724 65416 16725 65456
rect 16683 65407 16725 65416
rect 17067 65456 17109 65465
rect 17067 65416 17068 65456
rect 17108 65416 17109 65456
rect 17067 65407 17109 65416
rect 17163 65456 17205 65465
rect 17163 65416 17164 65456
rect 17204 65416 17205 65456
rect 17163 65407 17205 65416
rect 17635 65456 17693 65457
rect 17635 65416 17644 65456
rect 17684 65416 17693 65456
rect 17635 65415 17693 65416
rect 18123 65451 18165 65460
rect 18123 65411 18124 65451
rect 18164 65411 18165 65451
rect 15291 65397 15333 65406
rect 18123 65402 18165 65411
rect 3339 65365 3381 65374
rect 18979 65372 19037 65373
rect 18979 65332 18988 65372
rect 19028 65332 19037 65372
rect 18979 65331 19037 65332
rect 19363 65372 19421 65373
rect 19363 65332 19372 65372
rect 19412 65332 19421 65372
rect 19363 65331 19421 65332
rect 19747 65372 19805 65373
rect 19747 65332 19756 65372
rect 19796 65332 19805 65372
rect 19747 65331 19805 65332
rect 19563 65288 19605 65297
rect 19563 65248 19564 65288
rect 19604 65248 19605 65288
rect 19563 65239 19605 65248
rect 19947 65288 19989 65297
rect 19947 65248 19948 65288
rect 19988 65248 19989 65288
rect 19947 65239 19989 65248
rect 7275 65204 7317 65213
rect 7275 65164 7276 65204
rect 7316 65164 7317 65204
rect 7275 65155 7317 65164
rect 8907 65204 8949 65213
rect 8907 65164 8908 65204
rect 8948 65164 8949 65204
rect 8907 65155 8949 65164
rect 10539 65204 10581 65213
rect 10539 65164 10540 65204
rect 10580 65164 10581 65204
rect 10539 65155 10581 65164
rect 19179 65204 19221 65213
rect 19179 65164 19180 65204
rect 19220 65164 19221 65204
rect 19179 65155 19221 65164
rect 1152 65036 20352 65060
rect 1152 64996 3688 65036
rect 3728 64996 3770 65036
rect 3810 64996 3852 65036
rect 3892 64996 3934 65036
rect 3974 64996 4016 65036
rect 4056 64996 18808 65036
rect 18848 64996 18890 65036
rect 18930 64996 18972 65036
rect 19012 64996 19054 65036
rect 19094 64996 19136 65036
rect 19176 64996 20352 65036
rect 1152 64972 20352 64996
rect 19947 64868 19989 64877
rect 19947 64828 19948 64868
rect 19988 64828 19989 64868
rect 19947 64819 19989 64828
rect 8139 64700 8181 64709
rect 8139 64660 8140 64700
rect 8180 64660 8181 64700
rect 8139 64651 8181 64660
rect 10251 64700 10293 64709
rect 10251 64660 10252 64700
rect 10292 64660 10293 64700
rect 10251 64651 10293 64660
rect 10347 64700 10389 64709
rect 10347 64660 10348 64700
rect 10388 64660 10389 64700
rect 10347 64651 10389 64660
rect 19363 64700 19421 64701
rect 19363 64660 19372 64700
rect 19412 64660 19421 64700
rect 19363 64659 19421 64660
rect 19747 64700 19805 64701
rect 19747 64660 19756 64700
rect 19796 64660 19805 64700
rect 19747 64659 19805 64660
rect 9099 64630 9141 64639
rect 2563 64616 2621 64617
rect 2563 64576 2572 64616
rect 2612 64576 2621 64616
rect 2563 64575 2621 64576
rect 3811 64616 3869 64617
rect 3811 64576 3820 64616
rect 3860 64576 3869 64616
rect 3811 64575 3869 64576
rect 4195 64616 4253 64617
rect 4195 64576 4204 64616
rect 4244 64576 4253 64616
rect 4195 64575 4253 64576
rect 5443 64616 5501 64617
rect 5443 64576 5452 64616
rect 5492 64576 5501 64616
rect 5443 64575 5501 64576
rect 5827 64616 5885 64617
rect 5827 64576 5836 64616
rect 5876 64576 5885 64616
rect 5827 64575 5885 64576
rect 7075 64616 7133 64617
rect 7075 64576 7084 64616
rect 7124 64576 7133 64616
rect 7075 64575 7133 64576
rect 7563 64616 7605 64625
rect 7563 64576 7564 64616
rect 7604 64576 7605 64616
rect 7563 64567 7605 64576
rect 7659 64616 7701 64625
rect 7659 64576 7660 64616
rect 7700 64576 7701 64616
rect 7659 64567 7701 64576
rect 8043 64616 8085 64625
rect 8043 64576 8044 64616
rect 8084 64576 8085 64616
rect 8043 64567 8085 64576
rect 8611 64616 8669 64617
rect 8611 64576 8620 64616
rect 8660 64576 8669 64616
rect 9099 64590 9100 64630
rect 9140 64590 9141 64630
rect 11307 64630 11349 64639
rect 9099 64581 9141 64590
rect 9771 64616 9813 64625
rect 8611 64575 8669 64576
rect 9771 64576 9772 64616
rect 9812 64576 9813 64616
rect 9771 64567 9813 64576
rect 9867 64616 9909 64625
rect 9867 64576 9868 64616
rect 9908 64576 9909 64616
rect 9867 64567 9909 64576
rect 10819 64616 10877 64617
rect 10819 64576 10828 64616
rect 10868 64576 10877 64616
rect 11307 64590 11308 64630
rect 11348 64590 11349 64630
rect 11307 64581 11349 64590
rect 12355 64616 12413 64617
rect 10819 64575 10877 64576
rect 12355 64576 12364 64616
rect 12404 64576 12413 64616
rect 12355 64575 12413 64576
rect 13603 64616 13661 64617
rect 13603 64576 13612 64616
rect 13652 64576 13661 64616
rect 13603 64575 13661 64576
rect 13987 64616 14045 64617
rect 13987 64576 13996 64616
rect 14036 64576 14045 64616
rect 13987 64575 14045 64576
rect 15235 64616 15293 64617
rect 15235 64576 15244 64616
rect 15284 64576 15293 64616
rect 15235 64575 15293 64576
rect 15715 64616 15773 64617
rect 15715 64576 15724 64616
rect 15764 64576 15773 64616
rect 15715 64575 15773 64576
rect 16963 64616 17021 64617
rect 16963 64576 16972 64616
rect 17012 64576 17021 64616
rect 16963 64575 17021 64576
rect 17731 64616 17789 64617
rect 17731 64576 17740 64616
rect 17780 64576 17789 64616
rect 17731 64575 17789 64576
rect 18979 64616 19037 64617
rect 18979 64576 18988 64616
rect 19028 64576 19037 64616
rect 18979 64575 19037 64576
rect 5643 64532 5685 64541
rect 5643 64492 5644 64532
rect 5684 64492 5685 64532
rect 5643 64483 5685 64492
rect 11499 64532 11541 64541
rect 11499 64492 11500 64532
rect 11540 64492 11541 64532
rect 11499 64483 11541 64492
rect 4011 64448 4053 64457
rect 4011 64408 4012 64448
rect 4052 64408 4053 64448
rect 4011 64399 4053 64408
rect 7275 64448 7317 64457
rect 7275 64408 7276 64448
rect 7316 64408 7317 64448
rect 7275 64399 7317 64408
rect 9291 64448 9333 64457
rect 9291 64408 9292 64448
rect 9332 64408 9333 64448
rect 9291 64399 9333 64408
rect 13803 64448 13845 64457
rect 13803 64408 13804 64448
rect 13844 64408 13845 64448
rect 13803 64399 13845 64408
rect 15435 64448 15477 64457
rect 15435 64408 15436 64448
rect 15476 64408 15477 64448
rect 15435 64399 15477 64408
rect 17163 64448 17205 64457
rect 17163 64408 17164 64448
rect 17204 64408 17205 64448
rect 17163 64399 17205 64408
rect 19179 64448 19221 64457
rect 19179 64408 19180 64448
rect 19220 64408 19221 64448
rect 19179 64399 19221 64408
rect 19563 64448 19605 64457
rect 19563 64408 19564 64448
rect 19604 64408 19605 64448
rect 19563 64399 19605 64408
rect 1152 64280 20452 64304
rect 1152 64240 4928 64280
rect 4968 64240 5010 64280
rect 5050 64240 5092 64280
rect 5132 64240 5174 64280
rect 5214 64240 5256 64280
rect 5296 64240 20048 64280
rect 20088 64240 20130 64280
rect 20170 64240 20212 64280
rect 20252 64240 20294 64280
rect 20334 64240 20376 64280
rect 20416 64240 20452 64280
rect 1152 64216 20452 64240
rect 19179 64112 19221 64121
rect 19179 64072 19180 64112
rect 19220 64072 19221 64112
rect 19179 64063 19221 64072
rect 19947 64112 19989 64121
rect 19947 64072 19948 64112
rect 19988 64072 19989 64112
rect 19947 64063 19989 64072
rect 5163 64028 5205 64037
rect 5163 63988 5164 64028
rect 5204 63988 5205 64028
rect 5163 63979 5205 63988
rect 8139 64028 8181 64037
rect 8139 63988 8140 64028
rect 8180 63988 8181 64028
rect 8139 63979 8181 63988
rect 12555 64028 12597 64037
rect 12555 63988 12556 64028
rect 12596 63988 12597 64028
rect 12555 63979 12597 63988
rect 15627 64028 15669 64037
rect 15627 63988 15628 64028
rect 15668 63988 15669 64028
rect 15627 63979 15669 63988
rect 1699 63944 1757 63945
rect 1699 63904 1708 63944
rect 1748 63904 1757 63944
rect 1699 63903 1757 63904
rect 2947 63944 3005 63945
rect 2947 63904 2956 63944
rect 2996 63904 3005 63944
rect 2947 63903 3005 63904
rect 3435 63944 3477 63953
rect 3435 63904 3436 63944
rect 3476 63904 3477 63944
rect 3435 63895 3477 63904
rect 3531 63944 3573 63953
rect 3531 63904 3532 63944
rect 3572 63904 3573 63944
rect 3531 63895 3573 63904
rect 4011 63944 4053 63953
rect 4011 63904 4012 63944
rect 4052 63904 4053 63944
rect 4011 63895 4053 63904
rect 4483 63944 4541 63945
rect 4483 63904 4492 63944
rect 4532 63904 4541 63944
rect 4483 63903 4541 63904
rect 4971 63939 5013 63948
rect 4971 63899 4972 63939
rect 5012 63899 5013 63939
rect 4971 63890 5013 63899
rect 6411 63944 6453 63953
rect 6411 63904 6412 63944
rect 6452 63904 6453 63944
rect 6411 63895 6453 63904
rect 6507 63944 6549 63953
rect 6507 63904 6508 63944
rect 6548 63904 6549 63944
rect 6507 63895 6549 63904
rect 7459 63944 7517 63945
rect 7459 63904 7468 63944
rect 7508 63904 7517 63944
rect 7459 63903 7517 63904
rect 7947 63939 7989 63948
rect 7947 63899 7948 63939
rect 7988 63899 7989 63939
rect 9091 63944 9149 63945
rect 9091 63904 9100 63944
rect 9140 63904 9149 63944
rect 9091 63903 9149 63904
rect 10339 63944 10397 63945
rect 10339 63904 10348 63944
rect 10388 63904 10397 63944
rect 10339 63903 10397 63904
rect 10827 63944 10869 63953
rect 10827 63904 10828 63944
rect 10868 63904 10869 63944
rect 7947 63890 7989 63899
rect 10827 63895 10869 63904
rect 10923 63944 10965 63953
rect 10923 63904 10924 63944
rect 10964 63904 10965 63944
rect 10923 63895 10965 63904
rect 11403 63944 11445 63953
rect 11403 63904 11404 63944
rect 11444 63904 11445 63944
rect 11403 63895 11445 63904
rect 11875 63944 11933 63945
rect 11875 63904 11884 63944
rect 11924 63904 11933 63944
rect 11875 63903 11933 63904
rect 12363 63939 12405 63948
rect 12363 63899 12364 63939
rect 12404 63899 12405 63939
rect 12363 63890 12405 63899
rect 13899 63944 13941 63953
rect 13899 63904 13900 63944
rect 13940 63904 13941 63944
rect 13899 63895 13941 63904
rect 13995 63944 14037 63953
rect 13995 63904 13996 63944
rect 14036 63904 14037 63944
rect 13995 63895 14037 63904
rect 14947 63944 15005 63945
rect 14947 63904 14956 63944
rect 14996 63904 15005 63944
rect 14947 63903 15005 63904
rect 15435 63939 15477 63948
rect 15435 63899 15436 63939
rect 15476 63899 15477 63939
rect 15435 63890 15477 63899
rect 17451 63944 17493 63953
rect 17451 63904 17452 63944
rect 17492 63904 17493 63944
rect 17451 63895 17493 63904
rect 17547 63944 17589 63953
rect 17547 63904 17548 63944
rect 17588 63904 17589 63944
rect 17547 63895 17589 63904
rect 18499 63944 18557 63945
rect 18499 63904 18508 63944
rect 18548 63904 18557 63944
rect 18499 63903 18557 63904
rect 19035 63934 19077 63943
rect 19035 63894 19036 63934
rect 19076 63894 19077 63934
rect 19035 63885 19077 63894
rect 3915 63860 3957 63869
rect 3915 63820 3916 63860
rect 3956 63820 3957 63860
rect 3915 63811 3957 63820
rect 6891 63860 6933 63869
rect 6891 63820 6892 63860
rect 6932 63820 6933 63860
rect 6891 63811 6933 63820
rect 6987 63860 7029 63869
rect 6987 63820 6988 63860
rect 7028 63820 7029 63860
rect 6987 63811 7029 63820
rect 11307 63860 11349 63869
rect 11307 63820 11308 63860
rect 11348 63820 11349 63860
rect 11307 63811 11349 63820
rect 14379 63860 14421 63869
rect 14379 63820 14380 63860
rect 14420 63820 14421 63860
rect 14379 63811 14421 63820
rect 14475 63860 14517 63869
rect 14475 63820 14476 63860
rect 14516 63820 14517 63860
rect 14475 63811 14517 63820
rect 17931 63860 17973 63869
rect 17931 63820 17932 63860
rect 17972 63820 17973 63860
rect 17931 63811 17973 63820
rect 18027 63860 18069 63869
rect 18027 63820 18028 63860
rect 18068 63820 18069 63860
rect 18027 63811 18069 63820
rect 19363 63860 19421 63861
rect 19363 63820 19372 63860
rect 19412 63820 19421 63860
rect 19363 63819 19421 63820
rect 19747 63860 19805 63861
rect 19747 63820 19756 63860
rect 19796 63820 19805 63860
rect 19747 63819 19805 63820
rect 10539 63776 10581 63785
rect 10539 63736 10540 63776
rect 10580 63736 10581 63776
rect 10539 63727 10581 63736
rect 19563 63776 19605 63785
rect 19563 63736 19564 63776
rect 19604 63736 19605 63776
rect 19563 63727 19605 63736
rect 3147 63692 3189 63701
rect 3147 63652 3148 63692
rect 3188 63652 3189 63692
rect 3147 63643 3189 63652
rect 1152 63524 20352 63548
rect 1152 63484 3688 63524
rect 3728 63484 3770 63524
rect 3810 63484 3852 63524
rect 3892 63484 3934 63524
rect 3974 63484 4016 63524
rect 4056 63484 18808 63524
rect 18848 63484 18890 63524
rect 18930 63484 18972 63524
rect 19012 63484 19054 63524
rect 19094 63484 19136 63524
rect 19176 63484 20352 63524
rect 1152 63460 20352 63484
rect 10443 63356 10485 63365
rect 10443 63316 10444 63356
rect 10484 63316 10485 63356
rect 10443 63307 10485 63316
rect 8811 63272 8853 63281
rect 8811 63232 8812 63272
rect 8852 63232 8853 63272
rect 8811 63223 8853 63232
rect 17163 63272 17205 63281
rect 17163 63232 17164 63272
rect 17204 63232 17205 63272
rect 17163 63223 17205 63232
rect 19659 63272 19701 63281
rect 19659 63232 19660 63272
rect 19700 63232 19701 63272
rect 19659 63223 19701 63232
rect 3435 63188 3477 63197
rect 3435 63148 3436 63188
rect 3476 63148 3477 63188
rect 3435 63139 3477 63148
rect 19459 63188 19517 63189
rect 19459 63148 19468 63188
rect 19508 63148 19517 63188
rect 19459 63147 19517 63148
rect 4395 63118 4437 63127
rect 2859 63104 2901 63113
rect 2859 63064 2860 63104
rect 2900 63064 2901 63104
rect 2859 63055 2901 63064
rect 2955 63104 2997 63113
rect 2955 63064 2956 63104
rect 2996 63064 2997 63104
rect 2955 63055 2997 63064
rect 3339 63104 3381 63113
rect 3339 63064 3340 63104
rect 3380 63064 3381 63104
rect 3339 63055 3381 63064
rect 3907 63104 3965 63105
rect 3907 63064 3916 63104
rect 3956 63064 3965 63104
rect 4395 63078 4396 63118
rect 4436 63078 4437 63118
rect 19131 63113 19173 63122
rect 4395 63069 4437 63078
rect 5635 63104 5693 63105
rect 3907 63063 3965 63064
rect 5635 63064 5644 63104
rect 5684 63064 5693 63104
rect 5635 63063 5693 63064
rect 6883 63104 6941 63105
rect 6883 63064 6892 63104
rect 6932 63064 6941 63104
rect 6883 63063 6941 63064
rect 7363 63104 7421 63105
rect 7363 63064 7372 63104
rect 7412 63064 7421 63104
rect 7363 63063 7421 63064
rect 8611 63104 8669 63105
rect 8611 63064 8620 63104
rect 8660 63064 8669 63104
rect 8611 63063 8669 63064
rect 8995 63104 9053 63105
rect 8995 63064 9004 63104
rect 9044 63064 9053 63104
rect 8995 63063 9053 63064
rect 10243 63104 10301 63105
rect 10243 63064 10252 63104
rect 10292 63064 10301 63104
rect 10243 63063 10301 63064
rect 10627 63104 10685 63105
rect 10627 63064 10636 63104
rect 10676 63064 10685 63104
rect 10627 63063 10685 63064
rect 11875 63104 11933 63105
rect 11875 63064 11884 63104
rect 11924 63064 11933 63104
rect 11875 63063 11933 63064
rect 13795 63104 13853 63105
rect 13795 63064 13804 63104
rect 13844 63064 13853 63104
rect 13795 63063 13853 63064
rect 15043 63104 15101 63105
rect 15043 63064 15052 63104
rect 15092 63064 15101 63104
rect 15043 63063 15101 63064
rect 15523 63104 15581 63105
rect 15523 63064 15532 63104
rect 15572 63064 15581 63104
rect 15523 63063 15581 63064
rect 16771 63104 16829 63105
rect 16771 63064 16780 63104
rect 16820 63064 16829 63104
rect 16771 63063 16829 63064
rect 17547 63104 17589 63113
rect 17547 63064 17548 63104
rect 17588 63064 17589 63104
rect 17547 63055 17589 63064
rect 17643 63104 17685 63113
rect 17643 63064 17644 63104
rect 17684 63064 17685 63104
rect 17643 63055 17685 63064
rect 18027 63104 18069 63113
rect 18027 63064 18028 63104
rect 18068 63064 18069 63104
rect 18027 63055 18069 63064
rect 18123 63104 18165 63113
rect 18123 63064 18124 63104
rect 18164 63064 18165 63104
rect 18123 63055 18165 63064
rect 18595 63104 18653 63105
rect 18595 63064 18604 63104
rect 18644 63064 18653 63104
rect 19131 63073 19132 63113
rect 19172 63073 19173 63113
rect 19131 63064 19173 63073
rect 18595 63063 18653 63064
rect 4587 63020 4629 63029
rect 4587 62980 4588 63020
rect 4628 62980 4629 63020
rect 4587 62971 4629 62980
rect 7083 63020 7125 63029
rect 7083 62980 7084 63020
rect 7124 62980 7125 63020
rect 7083 62971 7125 62980
rect 16971 63020 17013 63029
rect 16971 62980 16972 63020
rect 17012 62980 17013 63020
rect 16971 62971 17013 62980
rect 19275 63020 19317 63029
rect 19275 62980 19276 63020
rect 19316 62980 19317 63020
rect 19275 62971 19317 62980
rect 12075 62936 12117 62945
rect 12075 62896 12076 62936
rect 12116 62896 12117 62936
rect 12075 62887 12117 62896
rect 15243 62936 15285 62945
rect 15243 62896 15244 62936
rect 15284 62896 15285 62936
rect 15243 62887 15285 62896
rect 17155 62936 17213 62937
rect 17155 62896 17164 62936
rect 17204 62896 17213 62936
rect 17155 62895 17213 62896
rect 1152 62768 20452 62792
rect 1152 62728 4928 62768
rect 4968 62728 5010 62768
rect 5050 62728 5092 62768
rect 5132 62728 5174 62768
rect 5214 62728 5256 62768
rect 5296 62728 20048 62768
rect 20088 62728 20130 62768
rect 20170 62728 20212 62768
rect 20252 62728 20294 62768
rect 20334 62728 20376 62768
rect 20416 62728 20452 62768
rect 1152 62704 20452 62728
rect 9291 62600 9333 62609
rect 9291 62560 9292 62600
rect 9332 62560 9333 62600
rect 9291 62551 9333 62560
rect 16779 62600 16821 62609
rect 16779 62560 16780 62600
rect 16820 62560 16821 62600
rect 16779 62551 16821 62560
rect 19467 62600 19509 62609
rect 19467 62560 19468 62600
rect 19508 62560 19509 62600
rect 19467 62551 19509 62560
rect 19851 62600 19893 62609
rect 19851 62560 19852 62600
rect 19892 62560 19893 62600
rect 19851 62551 19893 62560
rect 20235 62600 20277 62609
rect 20235 62560 20236 62600
rect 20276 62560 20277 62600
rect 20235 62551 20277 62560
rect 15627 62516 15669 62525
rect 15627 62476 15628 62516
rect 15668 62476 15669 62516
rect 15627 62467 15669 62476
rect 1219 62432 1277 62433
rect 1219 62392 1228 62432
rect 1268 62392 1277 62432
rect 1219 62391 1277 62392
rect 2467 62432 2525 62433
rect 2467 62392 2476 62432
rect 2516 62392 2525 62432
rect 2467 62391 2525 62392
rect 2947 62432 3005 62433
rect 2947 62392 2956 62432
rect 2996 62392 3005 62432
rect 2947 62391 3005 62392
rect 4195 62432 4253 62433
rect 4195 62392 4204 62432
rect 4244 62392 4253 62432
rect 4195 62391 4253 62392
rect 4579 62432 4637 62433
rect 4579 62392 4588 62432
rect 4628 62392 4637 62432
rect 4579 62391 4637 62392
rect 5827 62432 5885 62433
rect 5827 62392 5836 62432
rect 5876 62392 5885 62432
rect 5827 62391 5885 62392
rect 7563 62432 7605 62441
rect 7563 62392 7564 62432
rect 7604 62392 7605 62432
rect 7563 62383 7605 62392
rect 7659 62432 7701 62441
rect 7659 62392 7660 62432
rect 7700 62392 7701 62432
rect 7659 62383 7701 62392
rect 8611 62432 8669 62433
rect 8611 62392 8620 62432
rect 8660 62392 8669 62432
rect 8611 62391 8669 62392
rect 9099 62427 9141 62436
rect 9099 62387 9100 62427
rect 9140 62387 9141 62427
rect 10915 62432 10973 62433
rect 10915 62392 10924 62432
rect 10964 62392 10973 62432
rect 10915 62391 10973 62392
rect 12163 62432 12221 62433
rect 12163 62392 12172 62432
rect 12212 62392 12221 62432
rect 12163 62391 12221 62392
rect 13899 62432 13941 62441
rect 13899 62392 13900 62432
rect 13940 62392 13941 62432
rect 9099 62378 9141 62387
rect 13899 62383 13941 62392
rect 13995 62432 14037 62441
rect 13995 62392 13996 62432
rect 14036 62392 14037 62432
rect 13995 62383 14037 62392
rect 14947 62432 15005 62433
rect 14947 62392 14956 62432
rect 14996 62392 15005 62432
rect 14947 62391 15005 62392
rect 15435 62427 15477 62436
rect 15435 62387 15436 62427
rect 15476 62387 15477 62427
rect 18019 62432 18077 62433
rect 18019 62392 18028 62432
rect 18068 62392 18077 62432
rect 18019 62391 18077 62392
rect 19267 62432 19325 62433
rect 19267 62392 19276 62432
rect 19316 62392 19325 62432
rect 19267 62391 19325 62392
rect 15435 62378 15477 62387
rect 8043 62348 8085 62357
rect 8043 62308 8044 62348
rect 8084 62308 8085 62348
rect 8043 62299 8085 62308
rect 8139 62348 8181 62357
rect 8139 62308 8140 62348
rect 8180 62308 8181 62348
rect 8139 62299 8181 62308
rect 14379 62348 14421 62357
rect 14379 62308 14380 62348
rect 14420 62308 14421 62348
rect 14379 62299 14421 62308
rect 14475 62348 14517 62357
rect 14475 62308 14476 62348
rect 14516 62308 14517 62348
rect 14475 62299 14517 62308
rect 16579 62348 16637 62349
rect 16579 62308 16588 62348
rect 16628 62308 16637 62348
rect 16579 62307 16637 62308
rect 19651 62348 19709 62349
rect 19651 62308 19660 62348
rect 19700 62308 19709 62348
rect 19651 62307 19709 62308
rect 20035 62348 20093 62349
rect 20035 62308 20044 62348
rect 20084 62308 20093 62348
rect 20035 62307 20093 62308
rect 2667 62180 2709 62189
rect 2667 62140 2668 62180
rect 2708 62140 2709 62180
rect 2667 62131 2709 62140
rect 4395 62180 4437 62189
rect 4395 62140 4396 62180
rect 4436 62140 4437 62180
rect 4395 62131 4437 62140
rect 6027 62180 6069 62189
rect 6027 62140 6028 62180
rect 6068 62140 6069 62180
rect 6027 62131 6069 62140
rect 12363 62180 12405 62189
rect 12363 62140 12364 62180
rect 12404 62140 12405 62180
rect 12363 62131 12405 62140
rect 1152 62012 20352 62036
rect 1152 61972 3688 62012
rect 3728 61972 3770 62012
rect 3810 61972 3852 62012
rect 3892 61972 3934 62012
rect 3974 61972 4016 62012
rect 4056 61972 18808 62012
rect 18848 61972 18890 62012
rect 18930 61972 18972 62012
rect 19012 61972 19054 62012
rect 19094 61972 19136 62012
rect 19176 61972 20352 62012
rect 1152 61948 20352 61972
rect 13899 61844 13941 61853
rect 13899 61804 13900 61844
rect 13940 61804 13941 61844
rect 13899 61795 13941 61804
rect 10251 61760 10293 61769
rect 10251 61720 10252 61760
rect 10292 61720 10293 61760
rect 10251 61711 10293 61720
rect 18795 61760 18837 61769
rect 18795 61720 18796 61760
rect 18836 61720 18837 61760
rect 18795 61711 18837 61720
rect 19947 61760 19989 61769
rect 19947 61720 19948 61760
rect 19988 61720 19989 61760
rect 19947 61711 19989 61720
rect 3435 61676 3477 61685
rect 3435 61636 3436 61676
rect 3476 61636 3477 61676
rect 3435 61627 3477 61636
rect 11115 61676 11157 61685
rect 11115 61636 11116 61676
rect 11156 61636 11157 61676
rect 11115 61627 11157 61636
rect 18595 61676 18653 61677
rect 18595 61636 18604 61676
rect 18644 61636 18653 61676
rect 18595 61635 18653 61636
rect 18979 61676 19037 61677
rect 18979 61636 18988 61676
rect 19028 61636 19037 61676
rect 18979 61635 19037 61636
rect 19363 61676 19421 61677
rect 19363 61636 19372 61676
rect 19412 61636 19421 61676
rect 19363 61635 19421 61636
rect 19747 61676 19805 61677
rect 19747 61636 19756 61676
rect 19796 61636 19805 61676
rect 19747 61635 19805 61636
rect 10539 61611 10581 61620
rect 2859 61592 2901 61601
rect 2859 61552 2860 61592
rect 2900 61552 2901 61592
rect 2859 61543 2901 61552
rect 2955 61592 2997 61601
rect 2955 61552 2956 61592
rect 2996 61552 2997 61592
rect 2955 61543 2997 61552
rect 3339 61592 3381 61601
rect 4395 61597 4437 61606
rect 3339 61552 3340 61592
rect 3380 61552 3381 61592
rect 3339 61543 3381 61552
rect 3907 61592 3965 61593
rect 3907 61552 3916 61592
rect 3956 61552 3965 61592
rect 3907 61551 3965 61552
rect 4395 61557 4396 61597
rect 4436 61557 4437 61597
rect 4395 61548 4437 61557
rect 5347 61592 5405 61593
rect 5347 61552 5356 61592
rect 5396 61552 5405 61592
rect 5347 61551 5405 61552
rect 6595 61592 6653 61593
rect 6595 61552 6604 61592
rect 6644 61552 6653 61592
rect 6595 61551 6653 61552
rect 7171 61592 7229 61593
rect 7171 61552 7180 61592
rect 7220 61552 7229 61592
rect 7171 61551 7229 61552
rect 8419 61592 8477 61593
rect 8419 61552 8428 61592
rect 8468 61552 8477 61592
rect 8419 61551 8477 61552
rect 8803 61592 8861 61593
rect 8803 61552 8812 61592
rect 8852 61552 8861 61592
rect 8803 61551 8861 61552
rect 10051 61592 10109 61593
rect 10051 61552 10060 61592
rect 10100 61552 10109 61592
rect 10539 61571 10540 61611
rect 10580 61571 10581 61611
rect 12075 61606 12117 61615
rect 10539 61562 10581 61571
rect 10635 61592 10677 61601
rect 10051 61551 10109 61552
rect 10635 61552 10636 61592
rect 10676 61552 10677 61592
rect 10635 61543 10677 61552
rect 11019 61592 11061 61601
rect 11019 61552 11020 61592
rect 11060 61552 11061 61592
rect 11019 61543 11061 61552
rect 11587 61592 11645 61593
rect 11587 61552 11596 61592
rect 11636 61552 11645 61592
rect 12075 61566 12076 61606
rect 12116 61566 12117 61606
rect 12075 61557 12117 61566
rect 12451 61592 12509 61593
rect 11587 61551 11645 61552
rect 12451 61552 12460 61592
rect 12500 61552 12509 61592
rect 12451 61551 12509 61552
rect 13699 61592 13757 61593
rect 13699 61552 13708 61592
rect 13748 61552 13757 61592
rect 13699 61551 13757 61552
rect 14563 61592 14621 61593
rect 14563 61552 14572 61592
rect 14612 61552 14621 61592
rect 14563 61551 14621 61552
rect 15811 61592 15869 61593
rect 15811 61552 15820 61592
rect 15860 61552 15869 61592
rect 15811 61551 15869 61552
rect 16195 61592 16253 61593
rect 16195 61552 16204 61592
rect 16244 61552 16253 61592
rect 16195 61551 16253 61552
rect 17443 61592 17501 61593
rect 17443 61552 17452 61592
rect 17492 61552 17501 61592
rect 17443 61551 17501 61552
rect 12267 61508 12309 61517
rect 12267 61468 12268 61508
rect 12308 61468 12309 61508
rect 12267 61459 12309 61468
rect 4587 61424 4629 61433
rect 4587 61384 4588 61424
rect 4628 61384 4629 61424
rect 4587 61375 4629 61384
rect 6795 61424 6837 61433
rect 6795 61384 6796 61424
rect 6836 61384 6837 61424
rect 6795 61375 6837 61384
rect 8619 61424 8661 61433
rect 8619 61384 8620 61424
rect 8660 61384 8661 61424
rect 8619 61375 8661 61384
rect 16011 61424 16053 61433
rect 16011 61384 16012 61424
rect 16052 61384 16053 61424
rect 16011 61375 16053 61384
rect 17643 61424 17685 61433
rect 17643 61384 17644 61424
rect 17684 61384 17685 61424
rect 17643 61375 17685 61384
rect 19179 61424 19221 61433
rect 19179 61384 19180 61424
rect 19220 61384 19221 61424
rect 19179 61375 19221 61384
rect 19563 61424 19605 61433
rect 19563 61384 19564 61424
rect 19604 61384 19605 61424
rect 19563 61375 19605 61384
rect 1152 61256 20452 61280
rect 1152 61216 4928 61256
rect 4968 61216 5010 61256
rect 5050 61216 5092 61256
rect 5132 61216 5174 61256
rect 5214 61216 5256 61256
rect 5296 61216 20048 61256
rect 20088 61216 20130 61256
rect 20170 61216 20212 61256
rect 20252 61216 20294 61256
rect 20334 61216 20376 61256
rect 20416 61216 20452 61256
rect 1152 61192 20452 61216
rect 2859 61088 2901 61097
rect 2859 61048 2860 61088
rect 2900 61048 2901 61088
rect 2859 61039 2901 61048
rect 8907 61088 8949 61097
rect 8907 61048 8908 61088
rect 8948 61048 8949 61088
rect 8907 61039 8949 61048
rect 12459 61088 12501 61097
rect 12459 61048 12460 61088
rect 12500 61048 12501 61088
rect 12459 61039 12501 61048
rect 17835 61088 17877 61097
rect 17835 61048 17836 61088
rect 17876 61048 17877 61088
rect 17835 61039 17877 61048
rect 19851 61088 19893 61097
rect 19851 61048 19852 61088
rect 19892 61048 19893 61088
rect 19851 61039 19893 61048
rect 4875 61004 4917 61013
rect 4875 60964 4876 61004
rect 4916 60964 4917 61004
rect 4875 60955 4917 60964
rect 1411 60920 1469 60921
rect 1411 60880 1420 60920
rect 1460 60880 1469 60920
rect 1411 60879 1469 60880
rect 2659 60920 2717 60921
rect 2659 60880 2668 60920
rect 2708 60880 2717 60920
rect 2659 60879 2717 60880
rect 3147 60920 3189 60929
rect 3147 60880 3148 60920
rect 3188 60880 3189 60920
rect 3147 60871 3189 60880
rect 3243 60920 3285 60929
rect 3243 60880 3244 60920
rect 3284 60880 3285 60920
rect 3243 60871 3285 60880
rect 3723 60920 3765 60929
rect 3723 60880 3724 60920
rect 3764 60880 3765 60920
rect 3723 60871 3765 60880
rect 4195 60920 4253 60921
rect 4195 60880 4204 60920
rect 4244 60880 4253 60920
rect 4195 60879 4253 60880
rect 4683 60915 4725 60924
rect 4683 60875 4684 60915
rect 4724 60875 4725 60915
rect 5443 60920 5501 60921
rect 5443 60880 5452 60920
rect 5492 60880 5501 60920
rect 5443 60879 5501 60880
rect 6691 60920 6749 60921
rect 6691 60880 6700 60920
rect 6740 60880 6749 60920
rect 6691 60879 6749 60880
rect 7179 60920 7221 60929
rect 7179 60880 7180 60920
rect 7220 60880 7221 60920
rect 4683 60866 4725 60875
rect 7179 60871 7221 60880
rect 7275 60920 7317 60929
rect 7275 60880 7276 60920
rect 7316 60880 7317 60920
rect 7275 60871 7317 60880
rect 8227 60920 8285 60921
rect 8227 60880 8236 60920
rect 8276 60880 8285 60920
rect 8227 60879 8285 60880
rect 8715 60915 8757 60924
rect 8715 60875 8716 60915
rect 8756 60875 8757 60915
rect 9091 60920 9149 60921
rect 9091 60880 9100 60920
rect 9140 60880 9149 60920
rect 9091 60879 9149 60880
rect 10051 60920 10109 60921
rect 10051 60880 10060 60920
rect 10100 60880 10109 60920
rect 10051 60879 10109 60880
rect 10731 60920 10773 60929
rect 10731 60880 10732 60920
rect 10772 60880 10773 60920
rect 8715 60866 8757 60875
rect 10731 60871 10773 60880
rect 10827 60920 10869 60929
rect 10827 60880 10828 60920
rect 10868 60880 10869 60920
rect 10827 60871 10869 60880
rect 11779 60920 11837 60921
rect 11779 60880 11788 60920
rect 11828 60880 11837 60920
rect 13315 60920 13373 60921
rect 11779 60879 11837 60880
rect 12315 60910 12357 60919
rect 12315 60870 12316 60910
rect 12356 60870 12357 60910
rect 13315 60880 13324 60920
rect 13364 60880 13373 60920
rect 13315 60879 13373 60880
rect 14563 60920 14621 60921
rect 14563 60880 14572 60920
rect 14612 60880 14621 60920
rect 14563 60879 14621 60880
rect 16107 60920 16149 60929
rect 16107 60880 16108 60920
rect 16148 60880 16149 60920
rect 16107 60871 16149 60880
rect 16203 60920 16245 60929
rect 16203 60880 16204 60920
rect 16244 60880 16245 60920
rect 16203 60871 16245 60880
rect 17155 60920 17213 60921
rect 17155 60880 17164 60920
rect 17204 60880 17213 60920
rect 17155 60879 17213 60880
rect 17643 60915 17685 60924
rect 17643 60875 17644 60915
rect 17684 60875 17685 60915
rect 12315 60861 12357 60870
rect 17643 60866 17685 60875
rect 18123 60920 18165 60929
rect 18123 60880 18124 60920
rect 18164 60880 18165 60920
rect 18123 60871 18165 60880
rect 18219 60920 18261 60929
rect 18219 60880 18220 60920
rect 18260 60880 18261 60920
rect 18219 60871 18261 60880
rect 19171 60920 19229 60921
rect 19171 60880 19180 60920
rect 19220 60880 19229 60920
rect 19171 60879 19229 60880
rect 19659 60906 19701 60915
rect 19659 60866 19660 60906
rect 19700 60866 19701 60906
rect 19659 60857 19701 60866
rect 3627 60836 3669 60845
rect 3627 60796 3628 60836
rect 3668 60796 3669 60836
rect 3627 60787 3669 60796
rect 7659 60836 7701 60845
rect 7659 60796 7660 60836
rect 7700 60796 7701 60836
rect 7659 60787 7701 60796
rect 7755 60836 7797 60845
rect 7755 60796 7756 60836
rect 7796 60796 7797 60836
rect 7755 60787 7797 60796
rect 11211 60836 11253 60845
rect 11211 60796 11212 60836
rect 11252 60796 11253 60836
rect 11211 60787 11253 60796
rect 11307 60836 11349 60845
rect 11307 60796 11308 60836
rect 11348 60796 11349 60836
rect 11307 60787 11349 60796
rect 16587 60836 16629 60845
rect 16587 60796 16588 60836
rect 16628 60796 16629 60836
rect 16587 60787 16629 60796
rect 16683 60836 16725 60845
rect 16683 60796 16684 60836
rect 16724 60796 16725 60836
rect 16683 60787 16725 60796
rect 18603 60836 18645 60845
rect 18603 60796 18604 60836
rect 18644 60796 18645 60836
rect 18603 60787 18645 60796
rect 18699 60836 18741 60845
rect 18699 60796 18700 60836
rect 18740 60796 18741 60836
rect 18699 60787 18741 60796
rect 20035 60836 20093 60837
rect 20035 60796 20044 60836
rect 20084 60796 20093 60836
rect 20035 60795 20093 60796
rect 6891 60668 6933 60677
rect 6891 60628 6892 60668
rect 6932 60628 6933 60668
rect 6891 60619 6933 60628
rect 14763 60668 14805 60677
rect 14763 60628 14764 60668
rect 14804 60628 14805 60668
rect 14763 60619 14805 60628
rect 20235 60668 20277 60677
rect 20235 60628 20236 60668
rect 20276 60628 20277 60668
rect 20235 60619 20277 60628
rect 1152 60500 20352 60524
rect 1152 60460 3688 60500
rect 3728 60460 3770 60500
rect 3810 60460 3852 60500
rect 3892 60460 3934 60500
rect 3974 60460 4016 60500
rect 4056 60460 18808 60500
rect 18848 60460 18890 60500
rect 18930 60460 18972 60500
rect 19012 60460 19054 60500
rect 19094 60460 19136 60500
rect 19176 60460 20352 60500
rect 1152 60436 20352 60460
rect 2667 60332 2709 60341
rect 2667 60292 2668 60332
rect 2708 60292 2709 60332
rect 2667 60283 2709 60292
rect 10635 60332 10677 60341
rect 10635 60292 10636 60332
rect 10676 60292 10677 60332
rect 10635 60283 10677 60292
rect 17451 60332 17493 60341
rect 17451 60292 17452 60332
rect 17492 60292 17493 60332
rect 17451 60283 17493 60292
rect 19563 60332 19605 60341
rect 19563 60292 19564 60332
rect 19604 60292 19605 60332
rect 19563 60283 19605 60292
rect 6699 60164 6741 60173
rect 6699 60124 6700 60164
rect 6740 60124 6741 60164
rect 6699 60115 6741 60124
rect 13803 60164 13845 60173
rect 13803 60124 13804 60164
rect 13844 60124 13845 60164
rect 13803 60115 13845 60124
rect 19747 60164 19805 60165
rect 19747 60124 19756 60164
rect 19796 60124 19805 60164
rect 19747 60123 19805 60124
rect 7659 60094 7701 60103
rect 1219 60080 1277 60081
rect 1219 60040 1228 60080
rect 1268 60040 1277 60080
rect 1219 60039 1277 60040
rect 2467 60080 2525 60081
rect 2467 60040 2476 60080
rect 2516 60040 2525 60080
rect 2467 60039 2525 60040
rect 3043 60080 3101 60081
rect 3043 60040 3052 60080
rect 3092 60040 3101 60080
rect 3043 60039 3101 60040
rect 4291 60080 4349 60081
rect 4291 60040 4300 60080
rect 4340 60040 4349 60080
rect 4291 60039 4349 60040
rect 6123 60080 6165 60089
rect 6123 60040 6124 60080
rect 6164 60040 6165 60080
rect 6123 60031 6165 60040
rect 6219 60080 6261 60089
rect 6219 60040 6220 60080
rect 6260 60040 6261 60080
rect 6219 60031 6261 60040
rect 6603 60080 6645 60089
rect 6603 60040 6604 60080
rect 6644 60040 6645 60080
rect 6603 60031 6645 60040
rect 7171 60080 7229 60081
rect 7171 60040 7180 60080
rect 7220 60040 7229 60080
rect 7659 60054 7660 60094
rect 7700 60054 7701 60094
rect 14763 60094 14805 60103
rect 7659 60045 7701 60054
rect 9187 60080 9245 60081
rect 7171 60039 7229 60040
rect 9187 60040 9196 60080
rect 9236 60040 9245 60080
rect 9187 60039 9245 60040
rect 10435 60080 10493 60081
rect 10435 60040 10444 60080
rect 10484 60040 10493 60080
rect 10435 60039 10493 60040
rect 11491 60080 11549 60081
rect 11491 60040 11500 60080
rect 11540 60040 11549 60080
rect 11491 60039 11549 60040
rect 12739 60080 12797 60081
rect 12739 60040 12748 60080
rect 12788 60040 12797 60080
rect 12739 60039 12797 60040
rect 13227 60080 13269 60089
rect 13227 60040 13228 60080
rect 13268 60040 13269 60080
rect 13227 60031 13269 60040
rect 13323 60080 13365 60089
rect 13323 60040 13324 60080
rect 13364 60040 13365 60080
rect 13323 60031 13365 60040
rect 13707 60080 13749 60089
rect 13707 60040 13708 60080
rect 13748 60040 13749 60080
rect 13707 60031 13749 60040
rect 14275 60080 14333 60081
rect 14275 60040 14284 60080
rect 14324 60040 14333 60080
rect 14763 60054 14764 60094
rect 14804 60054 14805 60094
rect 14763 60045 14805 60054
rect 15147 60080 15189 60089
rect 14275 60039 14333 60040
rect 15147 60040 15148 60080
rect 15188 60040 15189 60080
rect 15147 60031 15189 60040
rect 15243 60080 15285 60089
rect 15243 60040 15244 60080
rect 15284 60040 15285 60080
rect 15243 60031 15285 60040
rect 15435 60080 15477 60089
rect 15435 60040 15436 60080
rect 15476 60040 15477 60080
rect 15435 60031 15477 60040
rect 16003 60080 16061 60081
rect 16003 60040 16012 60080
rect 16052 60040 16061 60080
rect 16003 60039 16061 60040
rect 17251 60080 17309 60081
rect 17251 60040 17260 60080
rect 17300 60040 17309 60080
rect 17251 60039 17309 60040
rect 18115 60080 18173 60081
rect 18115 60040 18124 60080
rect 18164 60040 18173 60080
rect 18115 60039 18173 60040
rect 19363 60080 19421 60081
rect 19363 60040 19372 60080
rect 19412 60040 19421 60080
rect 19363 60039 19421 60040
rect 12939 59996 12981 60005
rect 12939 59956 12940 59996
rect 12980 59956 12981 59996
rect 12939 59947 12981 59956
rect 14955 59996 14997 60005
rect 14955 59956 14956 59996
rect 14996 59956 14997 59996
rect 14955 59947 14997 59956
rect 4491 59912 4533 59921
rect 4491 59872 4492 59912
rect 4532 59872 4533 59912
rect 4491 59863 4533 59872
rect 7851 59912 7893 59921
rect 7851 59872 7852 59912
rect 7892 59872 7893 59912
rect 7851 59863 7893 59872
rect 15339 59912 15381 59921
rect 15339 59872 15340 59912
rect 15380 59872 15381 59912
rect 15339 59863 15381 59872
rect 19947 59912 19989 59921
rect 19947 59872 19948 59912
rect 19988 59872 19989 59912
rect 19947 59863 19989 59872
rect 1152 59744 20452 59768
rect 1152 59704 4928 59744
rect 4968 59704 5010 59744
rect 5050 59704 5092 59744
rect 5132 59704 5174 59744
rect 5214 59704 5256 59744
rect 5296 59704 20048 59744
rect 20088 59704 20130 59744
rect 20170 59704 20212 59744
rect 20252 59704 20294 59744
rect 20334 59704 20376 59744
rect 20416 59704 20452 59744
rect 1152 59680 20452 59704
rect 11307 59576 11349 59585
rect 11307 59536 11308 59576
rect 11348 59536 11349 59576
rect 11307 59527 11349 59536
rect 15435 59576 15477 59585
rect 15435 59536 15436 59576
rect 15476 59536 15477 59576
rect 15435 59527 15477 59536
rect 16875 59576 16917 59585
rect 16875 59536 16876 59576
rect 16916 59536 16917 59576
rect 16875 59527 16917 59536
rect 19179 59576 19221 59585
rect 19179 59536 19180 59576
rect 19220 59536 19221 59576
rect 19179 59527 19221 59536
rect 19947 59576 19989 59585
rect 19947 59536 19948 59576
rect 19988 59536 19989 59576
rect 19947 59527 19989 59536
rect 4875 59492 4917 59501
rect 4875 59452 4876 59492
rect 4916 59452 4917 59492
rect 4875 59443 4917 59452
rect 9291 59492 9333 59501
rect 9291 59452 9292 59492
rect 9332 59452 9333 59492
rect 9291 59443 9333 59452
rect 3147 59408 3189 59417
rect 3147 59368 3148 59408
rect 3188 59368 3189 59408
rect 3147 59359 3189 59368
rect 3243 59408 3285 59417
rect 3243 59368 3244 59408
rect 3284 59368 3285 59408
rect 3243 59359 3285 59368
rect 3723 59408 3765 59417
rect 3723 59368 3724 59408
rect 3764 59368 3765 59408
rect 3723 59359 3765 59368
rect 4195 59408 4253 59409
rect 4195 59368 4204 59408
rect 4244 59368 4253 59408
rect 4195 59367 4253 59368
rect 4683 59403 4725 59412
rect 4683 59363 4684 59403
rect 4724 59363 4725 59403
rect 6019 59408 6077 59409
rect 6019 59368 6028 59408
rect 6068 59368 6077 59408
rect 6019 59367 6077 59368
rect 7267 59408 7325 59409
rect 7267 59368 7276 59408
rect 7316 59368 7325 59408
rect 7267 59367 7325 59368
rect 7843 59408 7901 59409
rect 7843 59368 7852 59408
rect 7892 59368 7901 59408
rect 7843 59367 7901 59368
rect 9091 59408 9149 59409
rect 9091 59368 9100 59408
rect 9140 59368 9149 59408
rect 9091 59367 9149 59368
rect 9579 59408 9621 59417
rect 9579 59368 9580 59408
rect 9620 59368 9621 59408
rect 4683 59354 4725 59363
rect 9579 59359 9621 59368
rect 9675 59408 9717 59417
rect 9675 59368 9676 59408
rect 9716 59368 9717 59408
rect 9675 59359 9717 59368
rect 10627 59408 10685 59409
rect 10627 59368 10636 59408
rect 10676 59368 10685 59408
rect 13987 59408 14045 59409
rect 10627 59367 10685 59368
rect 11115 59394 11157 59403
rect 11115 59354 11116 59394
rect 11156 59354 11157 59394
rect 13987 59368 13996 59408
rect 14036 59368 14045 59408
rect 13987 59367 14045 59368
rect 15235 59408 15293 59409
rect 15235 59368 15244 59408
rect 15284 59368 15293 59408
rect 15235 59367 15293 59368
rect 15619 59408 15677 59409
rect 15619 59368 15628 59408
rect 15668 59368 15677 59408
rect 15915 59408 15957 59417
rect 15619 59367 15677 59368
rect 15723 59393 15765 59402
rect 11115 59345 11157 59354
rect 15723 59353 15724 59393
rect 15764 59353 15765 59393
rect 15915 59368 15916 59408
rect 15956 59368 15957 59408
rect 15915 59359 15957 59368
rect 16011 59408 16053 59417
rect 16011 59368 16012 59408
rect 16052 59368 16053 59408
rect 16011 59359 16053 59368
rect 16104 59408 16162 59409
rect 16104 59368 16113 59408
rect 16153 59368 16162 59408
rect 16104 59367 16162 59368
rect 17451 59408 17493 59417
rect 17451 59368 17452 59408
rect 17492 59368 17493 59408
rect 17451 59359 17493 59368
rect 17547 59408 17589 59417
rect 17547 59368 17548 59408
rect 17588 59368 17589 59408
rect 17547 59359 17589 59368
rect 17931 59408 17973 59417
rect 17931 59368 17932 59408
rect 17972 59368 17973 59408
rect 17931 59359 17973 59368
rect 18027 59408 18069 59417
rect 18027 59368 18028 59408
rect 18068 59368 18069 59408
rect 18027 59359 18069 59368
rect 18499 59408 18557 59409
rect 18499 59368 18508 59408
rect 18548 59368 18557 59408
rect 18499 59367 18557 59368
rect 19035 59398 19077 59407
rect 15723 59344 15765 59353
rect 19035 59358 19036 59398
rect 19076 59358 19077 59398
rect 19035 59349 19077 59358
rect 3627 59324 3669 59333
rect 3627 59284 3628 59324
rect 3668 59284 3669 59324
rect 3627 59275 3669 59284
rect 10059 59324 10101 59333
rect 10059 59284 10060 59324
rect 10100 59284 10101 59324
rect 10059 59275 10101 59284
rect 10155 59324 10197 59333
rect 10155 59284 10156 59324
rect 10196 59284 10197 59324
rect 10155 59275 10197 59284
rect 16675 59324 16733 59325
rect 16675 59284 16684 59324
rect 16724 59284 16733 59324
rect 16675 59283 16733 59284
rect 19363 59324 19421 59325
rect 19363 59284 19372 59324
rect 19412 59284 19421 59324
rect 19363 59283 19421 59284
rect 19747 59324 19805 59325
rect 19747 59284 19756 59324
rect 19796 59284 19805 59324
rect 19747 59283 19805 59284
rect 2763 59240 2805 59249
rect 2763 59200 2764 59240
rect 2804 59200 2805 59240
rect 2763 59191 2805 59200
rect 7467 59240 7509 59249
rect 7467 59200 7468 59240
rect 7508 59200 7509 59240
rect 7467 59191 7509 59200
rect 17067 59240 17109 59249
rect 17067 59200 17068 59240
rect 17108 59200 17109 59240
rect 17067 59191 17109 59200
rect 19563 59240 19605 59249
rect 19563 59200 19564 59240
rect 19604 59200 19605 59240
rect 19563 59191 19605 59200
rect 15627 59156 15669 59165
rect 15627 59116 15628 59156
rect 15668 59116 15669 59156
rect 15627 59107 15669 59116
rect 1152 58988 20352 59012
rect 1152 58948 3688 58988
rect 3728 58948 3770 58988
rect 3810 58948 3852 58988
rect 3892 58948 3934 58988
rect 3974 58948 4016 58988
rect 4056 58948 18808 58988
rect 18848 58948 18890 58988
rect 18930 58948 18972 58988
rect 19012 58948 19054 58988
rect 19094 58948 19136 58988
rect 19176 58948 20352 58988
rect 1152 58924 20352 58948
rect 15339 58820 15381 58829
rect 15339 58780 15340 58820
rect 15380 58780 15381 58820
rect 15339 58771 15381 58780
rect 19083 58820 19125 58829
rect 19083 58780 19084 58820
rect 19124 58780 19125 58820
rect 19083 58771 19125 58780
rect 19563 58820 19605 58829
rect 19563 58780 19564 58820
rect 19604 58780 19605 58820
rect 19563 58771 19605 58780
rect 19947 58820 19989 58829
rect 19947 58780 19948 58820
rect 19988 58780 19989 58820
rect 19947 58771 19989 58780
rect 3147 58736 3189 58745
rect 3147 58696 3148 58736
rect 3188 58696 3189 58736
rect 3147 58687 3189 58696
rect 5739 58652 5781 58661
rect 5739 58612 5740 58652
rect 5780 58612 5781 58652
rect 5739 58603 5781 58612
rect 5835 58652 5877 58661
rect 5835 58612 5836 58652
rect 5876 58612 5877 58652
rect 5835 58603 5877 58612
rect 12171 58652 12213 58661
rect 12171 58612 12172 58652
rect 12212 58612 12213 58652
rect 12171 58603 12213 58612
rect 12267 58652 12309 58661
rect 12267 58612 12268 58652
rect 12308 58612 12309 58652
rect 12267 58603 12309 58612
rect 19363 58652 19421 58653
rect 19363 58612 19372 58652
rect 19412 58612 19421 58652
rect 19363 58611 19421 58612
rect 19747 58652 19805 58653
rect 19747 58612 19756 58652
rect 19796 58612 19805 58652
rect 19747 58611 19805 58612
rect 1411 58568 1469 58569
rect 1411 58528 1420 58568
rect 1460 58528 1469 58568
rect 1411 58527 1469 58528
rect 2659 58568 2717 58569
rect 2659 58528 2668 58568
rect 2708 58528 2717 58568
rect 2659 58527 2717 58528
rect 3523 58568 3581 58569
rect 3523 58528 3532 58568
rect 3572 58528 3581 58568
rect 3523 58527 3581 58528
rect 4771 58568 4829 58569
rect 4771 58528 4780 58568
rect 4820 58528 4829 58568
rect 4771 58527 4829 58528
rect 5259 58568 5301 58577
rect 5259 58528 5260 58568
rect 5300 58528 5301 58568
rect 5259 58519 5301 58528
rect 5355 58568 5397 58577
rect 6795 58573 6837 58582
rect 5355 58528 5356 58568
rect 5396 58528 5397 58568
rect 5355 58519 5397 58528
rect 6307 58568 6365 58569
rect 6307 58528 6316 58568
rect 6356 58528 6365 58568
rect 6307 58527 6365 58528
rect 6795 58533 6796 58573
rect 6836 58533 6837 58573
rect 6795 58524 6837 58533
rect 7563 58568 7605 58577
rect 7563 58528 7564 58568
rect 7604 58528 7605 58568
rect 7563 58519 7605 58528
rect 7659 58568 7701 58577
rect 7659 58528 7660 58568
rect 7700 58528 7701 58568
rect 7659 58519 7701 58528
rect 8043 58568 8085 58577
rect 8043 58528 8044 58568
rect 8084 58528 8085 58568
rect 8043 58519 8085 58528
rect 8139 58568 8181 58577
rect 9099 58573 9141 58582
rect 13275 58577 13317 58586
rect 8139 58528 8140 58568
rect 8180 58528 8181 58568
rect 8139 58519 8181 58528
rect 8611 58568 8669 58569
rect 8611 58528 8620 58568
rect 8660 58528 8669 58568
rect 8611 58527 8669 58528
rect 9099 58533 9100 58573
rect 9140 58533 9141 58573
rect 9099 58524 9141 58533
rect 9955 58568 10013 58569
rect 9955 58528 9964 58568
rect 10004 58528 10013 58568
rect 9955 58527 10013 58528
rect 11203 58568 11261 58569
rect 11203 58528 11212 58568
rect 11252 58528 11261 58568
rect 11203 58527 11261 58528
rect 11691 58568 11733 58577
rect 11691 58528 11692 58568
rect 11732 58528 11733 58568
rect 11691 58519 11733 58528
rect 11787 58568 11829 58577
rect 11787 58528 11788 58568
rect 11828 58528 11829 58568
rect 11787 58519 11829 58528
rect 12739 58568 12797 58569
rect 12739 58528 12748 58568
rect 12788 58528 12797 58568
rect 13275 58537 13276 58577
rect 13316 58537 13317 58577
rect 13275 58528 13317 58537
rect 13699 58568 13757 58569
rect 13699 58528 13708 58568
rect 13748 58528 13757 58568
rect 12739 58527 12797 58528
rect 13699 58527 13757 58528
rect 14947 58568 15005 58569
rect 14947 58528 14956 58568
rect 14996 58528 15005 58568
rect 14947 58527 15005 58528
rect 15523 58568 15581 58569
rect 15523 58528 15532 58568
rect 15572 58528 15581 58568
rect 15523 58527 15581 58528
rect 16771 58568 16829 58569
rect 16771 58528 16780 58568
rect 16820 58528 16829 58568
rect 16771 58527 16829 58528
rect 16971 58568 17013 58577
rect 16971 58528 16972 58568
rect 17012 58528 17013 58568
rect 16971 58519 17013 58528
rect 17067 58568 17109 58577
rect 17067 58528 17068 58568
rect 17108 58528 17109 58568
rect 17067 58519 17109 58528
rect 17635 58568 17693 58569
rect 17635 58528 17644 58568
rect 17684 58528 17693 58568
rect 17635 58527 17693 58528
rect 18883 58568 18941 58569
rect 18883 58528 18892 58568
rect 18932 58528 18941 58568
rect 18883 58527 18941 58528
rect 4971 58484 5013 58493
rect 4971 58444 4972 58484
rect 5012 58444 5013 58484
rect 4971 58435 5013 58444
rect 6987 58484 7029 58493
rect 6987 58444 6988 58484
rect 7028 58444 7029 58484
rect 6987 58435 7029 58444
rect 9291 58484 9333 58493
rect 9291 58444 9292 58484
rect 9332 58444 9333 58484
rect 9291 58435 9333 58444
rect 11403 58484 11445 58493
rect 11403 58444 11404 58484
rect 11444 58444 11445 58484
rect 11403 58435 11445 58444
rect 13419 58484 13461 58493
rect 13419 58444 13420 58484
rect 13460 58444 13461 58484
rect 13419 58435 13461 58444
rect 2859 58400 2901 58409
rect 2859 58360 2860 58400
rect 2900 58360 2901 58400
rect 2859 58351 2901 58360
rect 15147 58400 15189 58409
rect 15147 58360 15148 58400
rect 15188 58360 15189 58400
rect 15147 58351 15189 58360
rect 17251 58400 17309 58401
rect 17251 58360 17260 58400
rect 17300 58360 17309 58400
rect 17251 58359 17309 58360
rect 1152 58232 20452 58256
rect 1152 58192 4928 58232
rect 4968 58192 5010 58232
rect 5050 58192 5092 58232
rect 5132 58192 5174 58232
rect 5214 58192 5256 58232
rect 5296 58192 20048 58232
rect 20088 58192 20130 58232
rect 20170 58192 20212 58232
rect 20252 58192 20294 58232
rect 20334 58192 20376 58232
rect 20416 58192 20452 58232
rect 1152 58168 20452 58192
rect 4099 58064 4157 58065
rect 4099 58024 4108 58064
rect 4148 58024 4157 58064
rect 4099 58023 4157 58024
rect 6795 58064 6837 58073
rect 6795 58024 6796 58064
rect 6836 58024 6837 58064
rect 6795 58015 6837 58024
rect 9003 58064 9045 58073
rect 9003 58024 9004 58064
rect 9044 58024 9045 58064
rect 9003 58015 9045 58024
rect 13323 58064 13365 58073
rect 13323 58024 13324 58064
rect 13364 58024 13365 58064
rect 13323 58015 13365 58024
rect 11211 57980 11253 57989
rect 11211 57940 11212 57980
rect 11252 57940 11253 57980
rect 11211 57931 11253 57940
rect 15627 57980 15669 57989
rect 15627 57940 15628 57980
rect 15668 57940 15669 57980
rect 15627 57931 15669 57940
rect 17355 57980 17397 57989
rect 17355 57940 17356 57980
rect 17396 57940 17397 57980
rect 17355 57931 17397 57940
rect 18507 57938 18549 57947
rect 1315 57896 1373 57897
rect 1315 57856 1324 57896
rect 1364 57856 1373 57896
rect 1315 57855 1373 57856
rect 2563 57896 2621 57897
rect 2563 57856 2572 57896
rect 2612 57856 2621 57896
rect 2563 57855 2621 57856
rect 3147 57896 3189 57905
rect 3147 57856 3148 57896
rect 3188 57856 3189 57896
rect 3147 57847 3189 57856
rect 3339 57896 3381 57905
rect 3339 57856 3340 57896
rect 3380 57856 3381 57896
rect 3339 57847 3381 57856
rect 3435 57896 3477 57905
rect 3435 57856 3436 57896
rect 3476 57856 3477 57896
rect 3435 57847 3477 57856
rect 3619 57896 3677 57897
rect 3619 57856 3628 57896
rect 3668 57856 3677 57896
rect 3619 57855 3677 57856
rect 3715 57896 3773 57897
rect 3715 57856 3724 57896
rect 3764 57856 3773 57896
rect 3715 57855 3773 57856
rect 3915 57896 3957 57905
rect 3915 57856 3916 57896
rect 3956 57856 3957 57896
rect 3915 57847 3957 57856
rect 4011 57896 4053 57905
rect 4011 57856 4012 57896
rect 4052 57856 4053 57896
rect 4011 57847 4053 57856
rect 4104 57896 4162 57897
rect 4104 57856 4113 57896
rect 4153 57856 4162 57896
rect 4104 57855 4162 57856
rect 5347 57896 5405 57897
rect 5347 57856 5356 57896
rect 5396 57856 5405 57896
rect 5347 57855 5405 57856
rect 6595 57896 6653 57897
rect 6595 57856 6604 57896
rect 6644 57856 6653 57896
rect 6595 57855 6653 57856
rect 7555 57896 7613 57897
rect 7555 57856 7564 57896
rect 7604 57856 7613 57896
rect 7555 57855 7613 57856
rect 8803 57896 8861 57897
rect 8803 57856 8812 57896
rect 8852 57856 8861 57896
rect 8803 57855 8861 57856
rect 11011 57896 11069 57897
rect 11011 57856 11020 57896
rect 11060 57856 11069 57896
rect 11011 57855 11069 57856
rect 11875 57896 11933 57897
rect 11875 57856 11884 57896
rect 11924 57856 11933 57896
rect 11875 57855 11933 57856
rect 13123 57896 13181 57897
rect 13123 57856 13132 57896
rect 13172 57856 13181 57896
rect 13123 57855 13181 57856
rect 13987 57896 14045 57897
rect 13987 57856 13996 57896
rect 14036 57856 14045 57896
rect 13987 57855 14045 57856
rect 15235 57896 15293 57897
rect 15235 57856 15244 57896
rect 15284 57856 15293 57896
rect 15235 57855 15293 57856
rect 15715 57896 15773 57897
rect 15715 57856 15724 57896
rect 15764 57856 15773 57896
rect 15715 57855 15773 57856
rect 15907 57896 15965 57897
rect 15907 57856 15916 57896
rect 15956 57856 15965 57896
rect 15907 57855 15965 57856
rect 17155 57896 17213 57897
rect 17155 57856 17164 57896
rect 17204 57856 17213 57896
rect 17155 57855 17213 57856
rect 17547 57896 17589 57905
rect 17547 57856 17548 57896
rect 17588 57856 17589 57896
rect 9763 57854 9821 57855
rect 9763 57814 9772 57854
rect 9812 57814 9821 57854
rect 17547 57847 17589 57856
rect 17643 57896 17685 57905
rect 17643 57856 17644 57896
rect 17684 57856 17685 57896
rect 17643 57847 17685 57856
rect 17739 57896 17781 57905
rect 17739 57856 17740 57896
rect 17780 57856 17781 57896
rect 17739 57847 17781 57856
rect 17835 57896 17877 57905
rect 17835 57856 17836 57896
rect 17876 57856 17877 57896
rect 17835 57847 17877 57856
rect 18115 57896 18173 57897
rect 18115 57856 18124 57896
rect 18164 57856 18173 57896
rect 18115 57855 18173 57856
rect 18411 57896 18453 57905
rect 18411 57856 18412 57896
rect 18452 57856 18453 57896
rect 18507 57898 18508 57938
rect 18548 57898 18549 57938
rect 18507 57889 18549 57898
rect 18987 57896 19029 57905
rect 18411 57847 18453 57856
rect 18987 57856 18988 57896
rect 19028 57856 19029 57896
rect 18987 57847 19029 57856
rect 19083 57896 19125 57905
rect 19083 57856 19084 57896
rect 19124 57856 19125 57896
rect 19083 57847 19125 57856
rect 19179 57896 19221 57905
rect 19179 57856 19180 57896
rect 19220 57856 19221 57896
rect 19179 57847 19221 57856
rect 19275 57896 19317 57905
rect 19275 57856 19276 57896
rect 19316 57856 19317 57896
rect 19275 57847 19317 57856
rect 19467 57896 19509 57905
rect 19467 57856 19468 57896
rect 19508 57856 19509 57896
rect 19467 57847 19509 57856
rect 19659 57896 19701 57905
rect 19659 57856 19660 57896
rect 19700 57856 19701 57896
rect 19659 57847 19701 57856
rect 9763 57813 9821 57814
rect 19843 57812 19901 57813
rect 19843 57772 19852 57812
rect 19892 57772 19901 57812
rect 19843 57771 19901 57772
rect 3427 57728 3485 57729
rect 3427 57688 3436 57728
rect 3476 57688 3485 57728
rect 3427 57687 3485 57688
rect 20043 57728 20085 57737
rect 20043 57688 20044 57728
rect 20084 57688 20085 57728
rect 20043 57679 20085 57688
rect 2763 57644 2805 57653
rect 2763 57604 2764 57644
rect 2804 57604 2805 57644
rect 2763 57595 2805 57604
rect 15435 57644 15477 57653
rect 15435 57604 15436 57644
rect 15476 57604 15477 57644
rect 15435 57595 15477 57604
rect 19659 57644 19701 57653
rect 19659 57604 19660 57644
rect 19700 57604 19701 57644
rect 18787 57602 18845 57603
rect 18787 57562 18796 57602
rect 18836 57562 18845 57602
rect 19659 57595 19701 57604
rect 18787 57561 18845 57562
rect 1152 57476 20352 57500
rect 1152 57436 3688 57476
rect 3728 57436 3770 57476
rect 3810 57436 3852 57476
rect 3892 57436 3934 57476
rect 3974 57436 4016 57476
rect 4056 57436 18808 57476
rect 18848 57436 18890 57476
rect 18930 57436 18972 57476
rect 19012 57436 19054 57476
rect 19094 57436 19136 57476
rect 19176 57436 20352 57476
rect 1152 57412 20352 57436
rect 2763 57308 2805 57317
rect 2763 57268 2764 57308
rect 2804 57268 2805 57308
rect 2763 57259 2805 57268
rect 7179 57308 7221 57317
rect 7179 57268 7180 57308
rect 7220 57268 7221 57308
rect 7179 57259 7221 57268
rect 17739 57308 17781 57317
rect 17739 57268 17740 57308
rect 17780 57268 17781 57308
rect 17739 57259 17781 57268
rect 19947 57224 19989 57233
rect 19947 57184 19948 57224
rect 19988 57184 19989 57224
rect 19947 57175 19989 57184
rect 3627 57140 3669 57149
rect 3627 57100 3628 57140
rect 3668 57100 3669 57140
rect 3627 57091 3669 57100
rect 10059 57140 10101 57149
rect 10059 57100 10060 57140
rect 10100 57100 10101 57140
rect 10059 57091 10101 57100
rect 10155 57140 10197 57149
rect 10155 57100 10156 57140
rect 10196 57100 10197 57140
rect 10155 57091 10197 57100
rect 18027 57140 18069 57149
rect 18027 57100 18028 57140
rect 18068 57100 18069 57140
rect 18027 57091 18069 57100
rect 4635 57065 4677 57074
rect 15243 57070 15285 57079
rect 1315 57056 1373 57057
rect 1315 57016 1324 57056
rect 1364 57016 1373 57056
rect 1315 57015 1373 57016
rect 2563 57056 2621 57057
rect 2563 57016 2572 57056
rect 2612 57016 2621 57056
rect 2563 57015 2621 57016
rect 3051 57056 3093 57065
rect 3051 57016 3052 57056
rect 3092 57016 3093 57056
rect 3051 57007 3093 57016
rect 3147 57056 3189 57065
rect 3147 57016 3148 57056
rect 3188 57016 3189 57056
rect 3147 57007 3189 57016
rect 3531 57056 3573 57065
rect 3531 57016 3532 57056
rect 3572 57016 3573 57056
rect 3531 57007 3573 57016
rect 4099 57056 4157 57057
rect 4099 57016 4108 57056
rect 4148 57016 4157 57056
rect 4635 57025 4636 57065
rect 4676 57025 4677 57065
rect 4635 57016 4677 57025
rect 4971 57056 5013 57065
rect 4971 57016 4972 57056
rect 5012 57016 5013 57056
rect 4099 57015 4157 57016
rect 4971 57007 5013 57016
rect 5067 57056 5109 57065
rect 5067 57016 5068 57056
rect 5108 57016 5109 57056
rect 5067 57007 5109 57016
rect 6987 57056 7029 57065
rect 6987 57016 6988 57056
rect 7028 57016 7029 57056
rect 6987 57007 7029 57016
rect 7179 57056 7221 57065
rect 7179 57016 7180 57056
rect 7220 57016 7221 57056
rect 7179 57007 7221 57016
rect 7371 57056 7413 57065
rect 7371 57016 7372 57056
rect 7412 57016 7413 57056
rect 7371 57007 7413 57016
rect 7467 57056 7509 57065
rect 7467 57016 7468 57056
rect 7508 57016 7509 57056
rect 7467 57007 7509 57016
rect 7563 57056 7605 57065
rect 7563 57016 7564 57056
rect 7604 57016 7605 57056
rect 7563 57007 7605 57016
rect 7843 57056 7901 57057
rect 7843 57016 7852 57056
rect 7892 57016 7901 57056
rect 7843 57015 7901 57016
rect 9091 57056 9149 57057
rect 9091 57016 9100 57056
rect 9140 57016 9149 57056
rect 9091 57015 9149 57016
rect 9579 57056 9621 57065
rect 9579 57016 9580 57056
rect 9620 57016 9621 57056
rect 9579 57007 9621 57016
rect 9675 57056 9717 57065
rect 11115 57061 11157 57070
rect 9675 57016 9676 57056
rect 9716 57016 9717 57056
rect 9675 57007 9717 57016
rect 10627 57056 10685 57057
rect 10627 57016 10636 57056
rect 10676 57016 10685 57056
rect 10627 57015 10685 57016
rect 11115 57021 11116 57061
rect 11156 57021 11157 57061
rect 11115 57012 11157 57021
rect 11971 57056 12029 57057
rect 11971 57016 11980 57056
rect 12020 57016 12029 57056
rect 11971 57015 12029 57016
rect 13219 57056 13277 57057
rect 13219 57016 13228 57056
rect 13268 57016 13277 57056
rect 13219 57015 13277 57016
rect 13707 57056 13749 57065
rect 13707 57016 13708 57056
rect 13748 57016 13749 57056
rect 13707 57007 13749 57016
rect 13803 57056 13845 57065
rect 13803 57016 13804 57056
rect 13844 57016 13845 57056
rect 13803 57007 13845 57016
rect 14187 57056 14229 57065
rect 14187 57016 14188 57056
rect 14228 57016 14229 57056
rect 14187 57007 14229 57016
rect 14283 57056 14325 57065
rect 14283 57016 14284 57056
rect 14324 57016 14325 57056
rect 14283 57007 14325 57016
rect 14755 57056 14813 57057
rect 14755 57016 14764 57056
rect 14804 57016 14813 57056
rect 15243 57030 15244 57070
rect 15284 57030 15285 57070
rect 20131 57070 20189 57071
rect 15243 57021 15285 57030
rect 16291 57056 16349 57057
rect 14755 57015 14813 57016
rect 16291 57016 16300 57056
rect 16340 57016 16349 57056
rect 16291 57015 16349 57016
rect 17539 57056 17597 57057
rect 17539 57016 17548 57056
rect 17588 57016 17597 57056
rect 17539 57015 17597 57016
rect 17931 57056 17973 57065
rect 17931 57016 17932 57056
rect 17972 57016 17973 57056
rect 17931 57007 17973 57016
rect 18123 57056 18165 57065
rect 18123 57016 18124 57056
rect 18164 57016 18165 57056
rect 18123 57007 18165 57016
rect 18307 57056 18365 57057
rect 18307 57016 18316 57056
rect 18356 57016 18365 57056
rect 18307 57015 18365 57016
rect 19555 57056 19613 57057
rect 19555 57016 19564 57056
rect 19604 57016 19613 57056
rect 19555 57015 19613 57016
rect 19947 57056 19989 57065
rect 19947 57016 19948 57056
rect 19988 57016 19989 57056
rect 20131 57030 20140 57070
rect 20180 57030 20189 57070
rect 20131 57029 20189 57030
rect 20227 57056 20285 57057
rect 19947 57007 19989 57016
rect 20227 57016 20236 57056
rect 20276 57016 20285 57056
rect 20227 57015 20285 57016
rect 4779 56972 4821 56981
rect 4779 56932 4780 56972
rect 4820 56932 4821 56972
rect 4779 56923 4821 56932
rect 9291 56972 9333 56981
rect 9291 56932 9292 56972
rect 9332 56932 9333 56972
rect 9291 56923 9333 56932
rect 11307 56972 11349 56981
rect 11307 56932 11308 56972
rect 11348 56932 11349 56972
rect 11307 56923 11349 56932
rect 13419 56972 13461 56981
rect 13419 56932 13420 56972
rect 13460 56932 13461 56972
rect 13419 56923 13461 56932
rect 19755 56972 19797 56981
rect 19755 56932 19756 56972
rect 19796 56932 19797 56972
rect 19755 56923 19797 56932
rect 5251 56888 5309 56889
rect 5251 56848 5260 56888
rect 5300 56848 5309 56888
rect 5251 56847 5309 56848
rect 7651 56888 7709 56889
rect 7651 56848 7660 56888
rect 7700 56848 7709 56888
rect 7651 56847 7709 56848
rect 15435 56888 15477 56897
rect 15435 56848 15436 56888
rect 15476 56848 15477 56888
rect 15435 56839 15477 56848
rect 17739 56888 17781 56897
rect 17739 56848 17740 56888
rect 17780 56848 17781 56888
rect 17739 56839 17781 56848
rect 1152 56720 20452 56744
rect 1152 56680 4928 56720
rect 4968 56680 5010 56720
rect 5050 56680 5092 56720
rect 5132 56680 5174 56720
rect 5214 56680 5256 56720
rect 5296 56680 20048 56720
rect 20088 56680 20130 56720
rect 20170 56680 20212 56720
rect 20252 56680 20294 56720
rect 20334 56680 20376 56720
rect 20416 56680 20452 56720
rect 1152 56656 20452 56680
rect 3051 56552 3093 56561
rect 3051 56512 3052 56552
rect 3092 56512 3093 56552
rect 3051 56503 3093 56512
rect 4875 56552 4917 56561
rect 4875 56512 4876 56552
rect 4916 56512 4917 56552
rect 4875 56503 4917 56512
rect 5067 56552 5109 56561
rect 5067 56512 5068 56552
rect 5108 56512 5109 56552
rect 5067 56503 5109 56512
rect 11115 56552 11157 56561
rect 11115 56512 11116 56552
rect 11156 56512 11157 56552
rect 11115 56503 11157 56512
rect 16683 56552 16725 56561
rect 16683 56512 16684 56552
rect 16724 56512 16725 56552
rect 16683 56503 16725 56512
rect 17155 56552 17213 56553
rect 17155 56512 17164 56552
rect 17204 56512 17213 56552
rect 17155 56511 17213 56512
rect 17635 56552 17693 56553
rect 17635 56512 17644 56552
rect 17684 56512 17693 56552
rect 17635 56511 17693 56512
rect 19659 56552 19701 56561
rect 19659 56512 19660 56552
rect 19700 56512 19701 56552
rect 19659 56503 19701 56512
rect 7947 56468 7989 56477
rect 7947 56428 7948 56468
rect 7988 56428 7989 56468
rect 7947 56419 7989 56428
rect 13419 56468 13461 56477
rect 13419 56428 13420 56468
rect 13460 56428 13461 56468
rect 13419 56419 13461 56428
rect 15531 56468 15573 56477
rect 15531 56428 15532 56468
rect 15572 56428 15573 56468
rect 15531 56419 15573 56428
rect 1603 56384 1661 56385
rect 1603 56344 1612 56384
rect 1652 56344 1661 56384
rect 1603 56343 1661 56344
rect 2851 56384 2909 56385
rect 2851 56344 2860 56384
rect 2900 56344 2909 56384
rect 2851 56343 2909 56344
rect 3427 56384 3485 56385
rect 3427 56344 3436 56384
rect 3476 56344 3485 56384
rect 3427 56343 3485 56344
rect 4675 56384 4733 56385
rect 4675 56344 4684 56384
rect 4724 56344 4733 56384
rect 4675 56343 4733 56344
rect 5155 56384 5213 56385
rect 5155 56344 5164 56384
rect 5204 56344 5213 56384
rect 5155 56343 5213 56344
rect 5827 56384 5885 56385
rect 5827 56344 5836 56384
rect 5876 56344 5885 56384
rect 5827 56343 5885 56344
rect 7075 56384 7133 56385
rect 7075 56344 7084 56384
rect 7124 56344 7133 56384
rect 7075 56343 7133 56344
rect 7555 56384 7613 56385
rect 7555 56344 7564 56384
rect 7604 56344 7613 56384
rect 7555 56343 7613 56344
rect 7851 56384 7893 56393
rect 7851 56344 7852 56384
rect 7892 56344 7893 56384
rect 7851 56335 7893 56344
rect 8427 56384 8469 56393
rect 8427 56344 8428 56384
rect 8468 56344 8469 56384
rect 8427 56335 8469 56344
rect 8619 56384 8661 56393
rect 8619 56344 8620 56384
rect 8660 56344 8661 56384
rect 8619 56335 8661 56344
rect 8707 56384 8765 56385
rect 8707 56344 8716 56384
rect 8756 56344 8765 56384
rect 8707 56343 8765 56344
rect 8907 56384 8949 56393
rect 8907 56344 8908 56384
rect 8948 56344 8949 56384
rect 8907 56335 8949 56344
rect 9099 56384 9141 56393
rect 9099 56344 9100 56384
rect 9140 56344 9141 56384
rect 9099 56335 9141 56344
rect 9667 56384 9725 56385
rect 9667 56344 9676 56384
rect 9716 56344 9725 56384
rect 9667 56343 9725 56344
rect 10915 56384 10973 56385
rect 10915 56344 10924 56384
rect 10964 56344 10973 56384
rect 10915 56343 10973 56344
rect 11971 56384 12029 56385
rect 11971 56344 11980 56384
rect 12020 56344 12029 56384
rect 11971 56343 12029 56344
rect 13219 56384 13277 56385
rect 13219 56344 13228 56384
rect 13268 56344 13277 56384
rect 13219 56343 13277 56344
rect 13803 56384 13845 56393
rect 13803 56344 13804 56384
rect 13844 56344 13845 56384
rect 13803 56335 13845 56344
rect 13899 56384 13941 56393
rect 13899 56344 13900 56384
rect 13940 56344 13941 56384
rect 13899 56335 13941 56344
rect 14283 56384 14325 56393
rect 14283 56344 14284 56384
rect 14324 56344 14325 56384
rect 14283 56335 14325 56344
rect 14379 56384 14421 56393
rect 14379 56344 14380 56384
rect 14420 56344 14421 56384
rect 14379 56335 14421 56344
rect 14851 56384 14909 56385
rect 14851 56344 14860 56384
rect 14900 56344 14909 56384
rect 14851 56343 14909 56344
rect 15339 56379 15381 56388
rect 15339 56339 15340 56379
rect 15380 56339 15381 56379
rect 15339 56330 15381 56339
rect 16875 56384 16917 56393
rect 16875 56344 16876 56384
rect 16916 56344 16917 56384
rect 16875 56335 16917 56344
rect 16971 56384 17013 56393
rect 16971 56344 16972 56384
rect 17012 56344 17013 56384
rect 16971 56335 17013 56344
rect 17355 56384 17397 56393
rect 17355 56344 17356 56384
rect 17396 56344 17397 56384
rect 17355 56335 17397 56344
rect 17451 56384 17493 56393
rect 17451 56344 17452 56384
rect 17492 56344 17493 56384
rect 17451 56335 17493 56344
rect 17931 56384 17973 56393
rect 17931 56344 17932 56384
rect 17972 56344 17973 56384
rect 17931 56335 17973 56344
rect 18027 56384 18069 56393
rect 18027 56344 18028 56384
rect 18068 56344 18069 56384
rect 18027 56335 18069 56344
rect 18507 56384 18549 56393
rect 18507 56344 18508 56384
rect 18548 56344 18549 56384
rect 18507 56335 18549 56344
rect 18979 56384 19037 56385
rect 18979 56344 18988 56384
rect 19028 56344 19037 56384
rect 19851 56384 19893 56393
rect 18979 56343 19037 56344
rect 19467 56370 19509 56379
rect 19467 56330 19468 56370
rect 19508 56330 19509 56370
rect 19851 56344 19852 56384
rect 19892 56344 19893 56384
rect 19851 56335 19893 56344
rect 20043 56384 20085 56393
rect 20043 56344 20044 56384
rect 20084 56344 20085 56384
rect 20043 56335 20085 56344
rect 20131 56384 20189 56385
rect 20131 56344 20140 56384
rect 20180 56344 20189 56384
rect 20131 56343 20189 56344
rect 19467 56321 19509 56330
rect 16483 56300 16541 56301
rect 16483 56260 16492 56300
rect 16532 56260 16541 56300
rect 16483 56259 16541 56260
rect 18411 56300 18453 56309
rect 18411 56260 18412 56300
rect 18452 56260 18453 56300
rect 18411 56251 18453 56260
rect 7275 56216 7317 56225
rect 7275 56176 7276 56216
rect 7316 56176 7317 56216
rect 7275 56167 7317 56176
rect 8227 56216 8285 56217
rect 8227 56176 8236 56216
rect 8276 56176 8285 56216
rect 8227 56175 8285 56176
rect 8427 56216 8469 56225
rect 8427 56176 8428 56216
rect 8468 56176 8469 56216
rect 8427 56167 8469 56176
rect 8907 56216 8949 56225
rect 8907 56176 8908 56216
rect 8948 56176 8949 56216
rect 8907 56167 8949 56176
rect 19851 56132 19893 56141
rect 19851 56092 19852 56132
rect 19892 56092 19893 56132
rect 19851 56083 19893 56092
rect 1152 55964 20352 55988
rect 1152 55924 3688 55964
rect 3728 55924 3770 55964
rect 3810 55924 3852 55964
rect 3892 55924 3934 55964
rect 3974 55924 4016 55964
rect 4056 55924 18808 55964
rect 18848 55924 18890 55964
rect 18930 55924 18972 55964
rect 19012 55924 19054 55964
rect 19094 55924 19136 55964
rect 19176 55924 20352 55964
rect 1152 55900 20352 55924
rect 5931 55796 5973 55805
rect 5931 55756 5932 55796
rect 5972 55756 5973 55796
rect 5931 55747 5973 55756
rect 17163 55796 17205 55805
rect 17163 55756 17164 55796
rect 17204 55756 17205 55796
rect 17163 55747 17205 55756
rect 19851 55796 19893 55805
rect 19851 55756 19852 55796
rect 19892 55756 19893 55796
rect 19851 55747 19893 55756
rect 2763 55712 2805 55721
rect 2763 55672 2764 55712
rect 2804 55672 2805 55712
rect 2763 55663 2805 55672
rect 10059 55712 10101 55721
rect 10059 55672 10060 55712
rect 10100 55672 10101 55712
rect 10059 55663 10101 55672
rect 10923 55628 10965 55637
rect 10923 55588 10924 55628
rect 10964 55588 10965 55628
rect 10923 55579 10965 55588
rect 1315 55544 1373 55545
rect 1315 55504 1324 55544
rect 1364 55504 1373 55544
rect 1315 55503 1373 55504
rect 2563 55544 2621 55545
rect 2563 55504 2572 55544
rect 2612 55504 2621 55544
rect 2563 55503 2621 55504
rect 3139 55544 3197 55545
rect 3139 55504 3148 55544
rect 3188 55504 3197 55544
rect 3139 55503 3197 55504
rect 3235 55544 3293 55545
rect 3235 55504 3244 55544
rect 3284 55504 3293 55544
rect 3235 55503 3293 55504
rect 3435 55544 3477 55553
rect 3435 55504 3436 55544
rect 3476 55504 3477 55544
rect 3435 55495 3477 55504
rect 3531 55544 3573 55553
rect 3531 55504 3532 55544
rect 3572 55504 3573 55544
rect 3531 55495 3573 55504
rect 3624 55544 3682 55545
rect 3624 55504 3633 55544
rect 3673 55504 3682 55544
rect 3624 55503 3682 55504
rect 3915 55544 3957 55553
rect 3915 55504 3916 55544
rect 3956 55504 3957 55544
rect 3915 55495 3957 55504
rect 4011 55544 4053 55553
rect 4011 55504 4012 55544
rect 4052 55504 4053 55544
rect 4011 55495 4053 55504
rect 4483 55544 4541 55545
rect 4483 55504 4492 55544
rect 4532 55504 4541 55544
rect 4483 55503 4541 55504
rect 5731 55544 5789 55545
rect 5731 55504 5740 55544
rect 5780 55504 5789 55544
rect 5731 55503 5789 55504
rect 6219 55544 6261 55553
rect 6219 55504 6220 55544
rect 6260 55504 6261 55544
rect 6219 55495 6261 55504
rect 6315 55544 6357 55553
rect 6315 55504 6316 55544
rect 6356 55504 6357 55544
rect 6315 55495 6357 55504
rect 6699 55544 6741 55553
rect 6699 55504 6700 55544
rect 6740 55504 6741 55544
rect 6699 55495 6741 55504
rect 6795 55544 6837 55553
rect 7755 55549 7797 55558
rect 11931 55553 11973 55562
rect 6795 55504 6796 55544
rect 6836 55504 6837 55544
rect 6795 55495 6837 55504
rect 7267 55544 7325 55545
rect 7267 55504 7276 55544
rect 7316 55504 7325 55544
rect 7267 55503 7325 55504
rect 7755 55509 7756 55549
rect 7796 55509 7797 55549
rect 7755 55500 7797 55509
rect 8139 55544 8181 55553
rect 8139 55504 8140 55544
rect 8180 55504 8181 55544
rect 8139 55495 8181 55504
rect 8235 55544 8277 55553
rect 8235 55504 8236 55544
rect 8276 55504 8277 55544
rect 8235 55495 8277 55504
rect 8331 55544 8373 55553
rect 8331 55504 8332 55544
rect 8372 55504 8373 55544
rect 8331 55495 8373 55504
rect 8427 55544 8469 55553
rect 8427 55504 8428 55544
rect 8468 55504 8469 55544
rect 8427 55495 8469 55504
rect 8611 55544 8669 55545
rect 8611 55504 8620 55544
rect 8660 55504 8669 55544
rect 8611 55503 8669 55504
rect 9859 55544 9917 55545
rect 9859 55504 9868 55544
rect 9908 55504 9917 55544
rect 9859 55503 9917 55504
rect 10347 55544 10389 55553
rect 10347 55504 10348 55544
rect 10388 55504 10389 55544
rect 10347 55495 10389 55504
rect 10443 55544 10485 55553
rect 10443 55504 10444 55544
rect 10484 55504 10485 55544
rect 10443 55495 10485 55504
rect 10827 55544 10869 55553
rect 10827 55504 10828 55544
rect 10868 55504 10869 55544
rect 10827 55495 10869 55504
rect 11395 55544 11453 55545
rect 11395 55504 11404 55544
rect 11444 55504 11453 55544
rect 11931 55513 11932 55553
rect 11972 55513 11973 55553
rect 11931 55504 11973 55513
rect 13219 55544 13277 55545
rect 13219 55504 13228 55544
rect 13268 55504 13277 55544
rect 11395 55503 11453 55504
rect 13219 55503 13277 55504
rect 14467 55544 14525 55545
rect 14467 55504 14476 55544
rect 14516 55504 14525 55544
rect 14467 55503 14525 55504
rect 15715 55544 15773 55545
rect 15715 55504 15724 55544
rect 15764 55504 15773 55544
rect 15715 55503 15773 55504
rect 16963 55544 17021 55545
rect 16963 55504 16972 55544
rect 17012 55504 17021 55544
rect 16963 55503 17021 55504
rect 17643 55544 17685 55553
rect 17643 55504 17644 55544
rect 17684 55504 17685 55544
rect 17643 55495 17685 55504
rect 17739 55544 17781 55553
rect 17739 55504 17740 55544
rect 17780 55504 17781 55544
rect 17739 55495 17781 55504
rect 18403 55544 18461 55545
rect 18403 55504 18412 55544
rect 18452 55504 18461 55544
rect 18403 55503 18461 55504
rect 19651 55544 19709 55545
rect 19651 55504 19660 55544
rect 19700 55504 19709 55544
rect 19651 55503 19709 55504
rect 7947 55460 7989 55469
rect 7947 55420 7948 55460
rect 7988 55420 7989 55460
rect 7947 55411 7989 55420
rect 12075 55460 12117 55469
rect 12075 55420 12076 55460
rect 12116 55420 12117 55460
rect 12075 55411 12117 55420
rect 3523 55376 3581 55377
rect 3523 55336 3532 55376
rect 3572 55336 3581 55376
rect 3523 55335 3581 55336
rect 4195 55376 4253 55377
rect 4195 55336 4204 55376
rect 4244 55336 4253 55376
rect 4195 55335 4253 55336
rect 14667 55376 14709 55385
rect 14667 55336 14668 55376
rect 14708 55336 14709 55376
rect 14667 55327 14709 55336
rect 17923 55376 17981 55377
rect 17923 55336 17932 55376
rect 17972 55336 17981 55376
rect 17923 55335 17981 55336
rect 1152 55208 20452 55232
rect 1152 55168 4928 55208
rect 4968 55168 5010 55208
rect 5050 55168 5092 55208
rect 5132 55168 5174 55208
rect 5214 55168 5256 55208
rect 5296 55168 20048 55208
rect 20088 55168 20130 55208
rect 20170 55168 20212 55208
rect 20252 55168 20294 55208
rect 20334 55168 20376 55208
rect 20416 55168 20452 55208
rect 1152 55144 20452 55168
rect 2859 55040 2901 55049
rect 2859 55000 2860 55040
rect 2900 55000 2901 55040
rect 2859 54991 2901 55000
rect 3051 55040 3093 55049
rect 3051 55000 3052 55040
rect 3092 55000 3093 55040
rect 3051 54991 3093 55000
rect 6987 55040 7029 55049
rect 6987 55000 6988 55040
rect 7028 55000 7029 55040
rect 6987 54991 7029 55000
rect 7651 55040 7709 55041
rect 7651 55000 7660 55040
rect 7700 55000 7709 55040
rect 7651 54999 7709 55000
rect 11979 55040 12021 55049
rect 11979 55000 11980 55040
rect 12020 55000 12021 55040
rect 11979 54991 12021 55000
rect 16299 55040 16341 55049
rect 16299 55000 16300 55040
rect 16340 55000 16341 55040
rect 16299 54991 16341 55000
rect 17827 55040 17885 55041
rect 17827 55000 17836 55040
rect 17876 55000 17885 55040
rect 17827 54999 17885 55000
rect 18115 55040 18173 55041
rect 18115 55000 18124 55040
rect 18164 55000 18173 55040
rect 18115 54999 18173 55000
rect 18507 55040 18549 55049
rect 18507 55000 18508 55040
rect 18548 55000 18549 55040
rect 18507 54991 18549 55000
rect 1411 54872 1469 54873
rect 1411 54832 1420 54872
rect 1460 54832 1469 54872
rect 1411 54831 1469 54832
rect 2659 54872 2717 54873
rect 2659 54832 2668 54872
rect 2708 54832 2717 54872
rect 2659 54831 2717 54832
rect 3139 54872 3197 54873
rect 3139 54832 3148 54872
rect 3188 54832 3197 54872
rect 3139 54831 3197 54832
rect 3331 54872 3389 54873
rect 3331 54832 3340 54872
rect 3380 54832 3389 54872
rect 3331 54831 3389 54832
rect 4579 54872 4637 54873
rect 4579 54832 4588 54872
rect 4628 54832 4637 54872
rect 4579 54831 4637 54832
rect 5539 54872 5597 54873
rect 5539 54832 5548 54872
rect 5588 54832 5597 54872
rect 5539 54831 5597 54832
rect 6787 54872 6845 54873
rect 6787 54832 6796 54872
rect 6836 54832 6845 54872
rect 6787 54831 6845 54832
rect 7371 54872 7413 54881
rect 7371 54832 7372 54872
rect 7412 54832 7413 54872
rect 7371 54823 7413 54832
rect 7467 54872 7509 54881
rect 7467 54832 7468 54872
rect 7508 54832 7509 54872
rect 7467 54823 7509 54832
rect 8227 54872 8285 54873
rect 8227 54832 8236 54872
rect 8276 54832 8285 54872
rect 8227 54831 8285 54832
rect 9475 54872 9533 54873
rect 9475 54832 9484 54872
rect 9524 54832 9533 54872
rect 9475 54831 9533 54832
rect 10059 54872 10101 54881
rect 10059 54832 10060 54872
rect 10100 54832 10101 54872
rect 10059 54823 10101 54832
rect 10155 54872 10197 54881
rect 10155 54832 10156 54872
rect 10196 54832 10197 54872
rect 10155 54823 10197 54832
rect 10251 54872 10293 54881
rect 10251 54832 10252 54872
rect 10292 54832 10293 54872
rect 10251 54823 10293 54832
rect 10347 54872 10389 54881
rect 10347 54832 10348 54872
rect 10388 54832 10389 54872
rect 10347 54823 10389 54832
rect 10531 54872 10589 54873
rect 10531 54832 10540 54872
rect 10580 54832 10589 54872
rect 10531 54831 10589 54832
rect 11779 54872 11837 54873
rect 11779 54832 11788 54872
rect 11828 54832 11837 54872
rect 11779 54831 11837 54832
rect 12931 54872 12989 54873
rect 12931 54832 12940 54872
rect 12980 54832 12989 54872
rect 12931 54831 12989 54832
rect 14179 54872 14237 54873
rect 14179 54832 14188 54872
rect 14228 54832 14237 54872
rect 14179 54831 14237 54832
rect 14851 54872 14909 54873
rect 14851 54832 14860 54872
rect 14900 54832 14909 54872
rect 14851 54831 14909 54832
rect 16099 54872 16157 54873
rect 16099 54832 16108 54872
rect 16148 54832 16157 54872
rect 16099 54831 16157 54832
rect 16683 54872 16725 54881
rect 16683 54832 16684 54872
rect 16724 54832 16725 54872
rect 16683 54823 16725 54832
rect 16875 54872 16917 54881
rect 16875 54832 16876 54872
rect 16916 54832 16917 54872
rect 16875 54823 16917 54832
rect 16963 54872 17021 54873
rect 16963 54832 16972 54872
rect 17012 54832 17021 54872
rect 16963 54831 17021 54832
rect 17355 54872 17397 54881
rect 17355 54832 17356 54872
rect 17396 54832 17397 54872
rect 17355 54823 17397 54832
rect 17451 54872 17493 54881
rect 17451 54832 17452 54872
rect 17492 54832 17493 54872
rect 17451 54823 17493 54832
rect 17547 54872 17589 54881
rect 17547 54832 17548 54872
rect 17588 54832 17589 54872
rect 17547 54823 17589 54832
rect 17643 54872 17685 54881
rect 17643 54832 17644 54872
rect 17684 54832 17685 54872
rect 17643 54823 17685 54832
rect 17923 54872 17981 54873
rect 17923 54832 17932 54872
rect 17972 54832 17981 54872
rect 17923 54831 17981 54832
rect 18691 54872 18749 54873
rect 18691 54832 18700 54872
rect 18740 54832 18749 54872
rect 18691 54831 18749 54832
rect 19939 54872 19997 54873
rect 19939 54832 19948 54872
rect 19988 54832 19997 54872
rect 19939 54831 19997 54832
rect 4779 54620 4821 54629
rect 4779 54580 4780 54620
rect 4820 54580 4821 54620
rect 4779 54571 4821 54580
rect 9675 54620 9717 54629
rect 9675 54580 9676 54620
rect 9716 54580 9717 54620
rect 9675 54571 9717 54580
rect 14379 54620 14421 54629
rect 14379 54580 14380 54620
rect 14420 54580 14421 54620
rect 14379 54571 14421 54580
rect 16683 54620 16725 54629
rect 16683 54580 16684 54620
rect 16724 54580 16725 54620
rect 16683 54571 16725 54580
rect 18507 54620 18549 54629
rect 18507 54580 18508 54620
rect 18548 54580 18549 54620
rect 18507 54571 18549 54580
rect 1152 54452 20352 54476
rect 1152 54412 3688 54452
rect 3728 54412 3770 54452
rect 3810 54412 3852 54452
rect 3892 54412 3934 54452
rect 3974 54412 4016 54452
rect 4056 54412 18808 54452
rect 18848 54412 18890 54452
rect 18930 54412 18972 54452
rect 19012 54412 19054 54452
rect 19094 54412 19136 54452
rect 19176 54412 20352 54452
rect 1152 54388 20352 54412
rect 15339 54200 15381 54209
rect 15339 54160 15340 54200
rect 15380 54160 15381 54200
rect 15339 54151 15381 54160
rect 3723 54116 3765 54125
rect 3723 54076 3724 54116
rect 3764 54076 3765 54116
rect 3723 54067 3765 54076
rect 17259 54116 17301 54125
rect 17259 54076 17260 54116
rect 17300 54076 17301 54116
rect 17259 54067 17301 54076
rect 19371 54116 19413 54125
rect 19371 54076 19372 54116
rect 19412 54076 19413 54116
rect 19371 54067 19413 54076
rect 4683 54046 4725 54055
rect 12939 54051 12981 54060
rect 1411 54032 1469 54033
rect 1411 53992 1420 54032
rect 1460 53992 1469 54032
rect 1411 53991 1469 53992
rect 2659 54032 2717 54033
rect 2659 53992 2668 54032
rect 2708 53992 2717 54032
rect 2659 53991 2717 53992
rect 3147 54032 3189 54041
rect 3147 53992 3148 54032
rect 3188 53992 3189 54032
rect 3147 53983 3189 53992
rect 3243 54032 3285 54041
rect 3243 53992 3244 54032
rect 3284 53992 3285 54032
rect 3243 53983 3285 53992
rect 3627 54032 3669 54041
rect 3627 53992 3628 54032
rect 3668 53992 3669 54032
rect 3627 53983 3669 53992
rect 4195 54032 4253 54033
rect 4195 53992 4204 54032
rect 4244 53992 4253 54032
rect 4683 54006 4684 54046
rect 4724 54006 4725 54046
rect 4683 53997 4725 54006
rect 5067 54032 5109 54041
rect 4195 53991 4253 53992
rect 5067 53992 5068 54032
rect 5108 53992 5109 54032
rect 5067 53983 5109 53992
rect 5163 54032 5205 54041
rect 5163 53992 5164 54032
rect 5204 53992 5205 54032
rect 5163 53983 5205 53992
rect 5259 54032 5301 54041
rect 5259 53992 5260 54032
rect 5300 53992 5301 54032
rect 5259 53983 5301 53992
rect 5731 54032 5789 54033
rect 5731 53992 5740 54032
rect 5780 53992 5789 54032
rect 5731 53991 5789 53992
rect 6979 54032 7037 54033
rect 6979 53992 6988 54032
rect 7028 53992 7037 54032
rect 6979 53991 7037 53992
rect 7267 54032 7325 54033
rect 7267 53992 7276 54032
rect 7316 53992 7325 54032
rect 7267 53991 7325 53992
rect 8515 54032 8573 54033
rect 8515 53992 8524 54032
rect 8564 53992 8573 54032
rect 8515 53991 8573 53992
rect 9003 54032 9045 54041
rect 9003 53992 9004 54032
rect 9044 53992 9045 54032
rect 9003 53983 9045 53992
rect 9099 54032 9141 54041
rect 9099 53992 9100 54032
rect 9140 53992 9141 54032
rect 9099 53983 9141 53992
rect 9483 54032 9525 54041
rect 9483 53992 9484 54032
rect 9524 53992 9525 54032
rect 9483 53983 9525 53992
rect 9579 54032 9621 54041
rect 10539 54037 10581 54046
rect 9579 53992 9580 54032
rect 9620 53992 9621 54032
rect 9579 53983 9621 53992
rect 10051 54032 10109 54033
rect 10051 53992 10060 54032
rect 10100 53992 10109 54032
rect 10051 53991 10109 53992
rect 10539 53997 10540 54037
rect 10580 53997 10581 54037
rect 10539 53988 10581 53997
rect 10915 54032 10973 54033
rect 10915 53992 10924 54032
rect 10964 53992 10973 54032
rect 10915 53991 10973 53992
rect 11203 54032 11261 54033
rect 11203 53992 11212 54032
rect 11252 53992 11261 54032
rect 11203 53991 11261 53992
rect 12451 54032 12509 54033
rect 12451 53992 12460 54032
rect 12500 53992 12509 54032
rect 12939 54011 12940 54051
rect 12980 54011 12981 54051
rect 14475 54046 14517 54055
rect 18411 54046 18453 54055
rect 12939 54002 12981 54011
rect 13035 54032 13077 54041
rect 12451 53991 12509 53992
rect 13035 53992 13036 54032
rect 13076 53992 13077 54032
rect 13035 53983 13077 53992
rect 13419 54032 13461 54041
rect 13419 53992 13420 54032
rect 13460 53992 13461 54032
rect 13419 53983 13461 53992
rect 13515 54032 13557 54041
rect 13515 53992 13516 54032
rect 13556 53992 13557 54032
rect 13515 53983 13557 53992
rect 13987 54032 14045 54033
rect 13987 53992 13996 54032
rect 14036 53992 14045 54032
rect 14475 54006 14476 54046
rect 14516 54006 14517 54046
rect 14475 53997 14517 54006
rect 15147 54032 15189 54041
rect 13987 53991 14045 53992
rect 15147 53992 15148 54032
rect 15188 53992 15189 54032
rect 15147 53983 15189 53992
rect 15339 54032 15381 54041
rect 15339 53992 15340 54032
rect 15380 53992 15381 54032
rect 15339 53983 15381 53992
rect 15531 54032 15573 54041
rect 15531 53992 15532 54032
rect 15572 53992 15573 54032
rect 15531 53983 15573 53992
rect 15627 54032 15669 54041
rect 15627 53992 15628 54032
rect 15668 53992 15669 54032
rect 15627 53983 15669 53992
rect 15723 54032 15765 54041
rect 15723 53992 15724 54032
rect 15764 53992 15765 54032
rect 15723 53983 15765 53992
rect 16203 54037 16245 54046
rect 16203 53997 16204 54037
rect 16244 53997 16245 54037
rect 16203 53988 16245 53997
rect 16675 54032 16733 54033
rect 16675 53992 16684 54032
rect 16724 53992 16733 54032
rect 16675 53991 16733 53992
rect 17163 54032 17205 54041
rect 17163 53992 17164 54032
rect 17204 53992 17205 54032
rect 17163 53983 17205 53992
rect 17643 54032 17685 54041
rect 17643 53992 17644 54032
rect 17684 53992 17685 54032
rect 17643 53983 17685 53992
rect 17739 54032 17781 54041
rect 17739 53992 17740 54032
rect 17780 53992 17781 54032
rect 18411 54006 18412 54046
rect 18452 54006 18453 54046
rect 18411 53997 18453 54006
rect 18883 54032 18941 54033
rect 17739 53983 17781 53992
rect 18883 53992 18892 54032
rect 18932 53992 18941 54032
rect 18883 53991 18941 53992
rect 19467 54032 19509 54041
rect 19467 53992 19468 54032
rect 19508 53992 19509 54032
rect 19467 53983 19509 53992
rect 19851 54032 19893 54041
rect 19851 53992 19852 54032
rect 19892 53992 19893 54032
rect 19851 53983 19893 53992
rect 19947 54032 19989 54041
rect 19947 53992 19948 54032
rect 19988 53992 19989 54032
rect 19947 53983 19989 53992
rect 2859 53948 2901 53957
rect 2859 53908 2860 53948
rect 2900 53908 2901 53948
rect 2859 53899 2901 53908
rect 8715 53948 8757 53957
rect 8715 53908 8716 53948
rect 8756 53908 8757 53948
rect 8715 53899 8757 53908
rect 14667 53948 14709 53957
rect 14667 53908 14668 53948
rect 14708 53908 14709 53948
rect 14667 53899 14709 53908
rect 16011 53948 16053 53957
rect 16011 53908 16012 53948
rect 16052 53908 16053 53948
rect 16011 53899 16053 53908
rect 4875 53864 4917 53873
rect 4875 53824 4876 53864
rect 4916 53824 4917 53864
rect 4875 53815 4917 53824
rect 5347 53864 5405 53865
rect 5347 53824 5356 53864
rect 5396 53824 5405 53864
rect 5347 53823 5405 53824
rect 5547 53864 5589 53873
rect 5547 53824 5548 53864
rect 5588 53824 5589 53864
rect 5547 53815 5589 53824
rect 10731 53864 10773 53873
rect 10731 53824 10732 53864
rect 10772 53824 10773 53864
rect 10731 53815 10773 53824
rect 11019 53864 11061 53873
rect 11019 53824 11020 53864
rect 11060 53824 11061 53864
rect 11019 53815 11061 53824
rect 12651 53864 12693 53873
rect 12651 53824 12652 53864
rect 12692 53824 12693 53864
rect 12651 53815 12693 53824
rect 15811 53864 15869 53865
rect 15811 53824 15820 53864
rect 15860 53824 15869 53864
rect 15811 53823 15869 53824
rect 18219 53864 18261 53873
rect 18219 53824 18220 53864
rect 18260 53824 18261 53864
rect 18219 53815 18261 53824
rect 1152 53696 20452 53720
rect 1152 53656 4928 53696
rect 4968 53656 5010 53696
rect 5050 53656 5092 53696
rect 5132 53656 5174 53696
rect 5214 53656 5256 53696
rect 5296 53656 20048 53696
rect 20088 53656 20130 53696
rect 20170 53656 20212 53696
rect 20252 53656 20294 53696
rect 20334 53656 20376 53696
rect 20416 53656 20452 53696
rect 1152 53632 20452 53656
rect 3051 53528 3093 53537
rect 3051 53488 3052 53528
rect 3092 53488 3093 53528
rect 3051 53479 3093 53488
rect 5835 53528 5877 53537
rect 5835 53488 5836 53528
rect 5876 53488 5877 53528
rect 5835 53479 5877 53488
rect 8035 53528 8093 53529
rect 8035 53488 8044 53528
rect 8084 53488 8093 53528
rect 8035 53487 8093 53488
rect 8803 53528 8861 53529
rect 8803 53488 8812 53528
rect 8852 53488 8861 53528
rect 8803 53487 8861 53488
rect 12747 53528 12789 53537
rect 12747 53488 12748 53528
rect 12788 53488 12789 53528
rect 12747 53479 12789 53488
rect 15243 53528 15285 53537
rect 15243 53488 15244 53528
rect 15284 53488 15285 53528
rect 15243 53479 15285 53488
rect 20139 53528 20181 53537
rect 20139 53488 20140 53528
rect 20180 53488 20181 53528
rect 20139 53479 20181 53488
rect 6027 53444 6069 53453
rect 6027 53404 6028 53444
rect 6068 53404 6069 53444
rect 6027 53395 6069 53404
rect 14859 53444 14901 53453
rect 14859 53404 14860 53444
rect 14900 53404 14901 53444
rect 14859 53395 14901 53404
rect 1219 53360 1277 53361
rect 1219 53320 1228 53360
rect 1268 53320 1277 53360
rect 1219 53319 1277 53320
rect 2467 53360 2525 53361
rect 2467 53320 2476 53360
rect 2516 53320 2525 53360
rect 2467 53319 2525 53320
rect 2955 53360 2997 53369
rect 2955 53320 2956 53360
rect 2996 53320 2997 53360
rect 2955 53311 2997 53320
rect 3147 53360 3189 53369
rect 3147 53320 3148 53360
rect 3188 53320 3189 53360
rect 3147 53311 3189 53320
rect 3243 53360 3285 53369
rect 3243 53320 3244 53360
rect 3284 53320 3285 53360
rect 3243 53311 3285 53320
rect 4387 53360 4445 53361
rect 4387 53320 4396 53360
rect 4436 53320 4445 53360
rect 4387 53319 4445 53320
rect 5635 53360 5693 53361
rect 5635 53320 5644 53360
rect 5684 53320 5693 53360
rect 5635 53319 5693 53320
rect 6219 53355 6261 53364
rect 6219 53315 6220 53355
rect 6260 53315 6261 53355
rect 6691 53360 6749 53361
rect 6691 53320 6700 53360
rect 6740 53320 6749 53360
rect 6691 53319 6749 53320
rect 7179 53360 7221 53369
rect 7179 53320 7180 53360
rect 7220 53320 7221 53360
rect 6219 53306 6261 53315
rect 7179 53311 7221 53320
rect 7659 53360 7701 53369
rect 7659 53320 7660 53360
rect 7700 53320 7701 53360
rect 7659 53311 7701 53320
rect 7755 53360 7797 53369
rect 7755 53320 7756 53360
rect 7796 53320 7797 53360
rect 7755 53311 7797 53320
rect 8235 53360 8277 53369
rect 8235 53320 8236 53360
rect 8276 53320 8277 53360
rect 8235 53311 8277 53320
rect 8331 53360 8373 53369
rect 8331 53320 8332 53360
rect 8372 53320 8373 53360
rect 8331 53311 8373 53320
rect 8523 53360 8565 53369
rect 8523 53320 8524 53360
rect 8564 53320 8565 53360
rect 8523 53311 8565 53320
rect 8619 53360 8661 53369
rect 8619 53320 8620 53360
rect 8660 53320 8661 53360
rect 8619 53311 8661 53320
rect 8995 53360 9053 53361
rect 8995 53320 9004 53360
rect 9044 53320 9053 53360
rect 8995 53319 9053 53320
rect 10243 53360 10301 53361
rect 10243 53320 10252 53360
rect 10292 53320 10301 53360
rect 10243 53319 10301 53320
rect 10819 53360 10877 53361
rect 10819 53320 10828 53360
rect 10868 53320 10877 53360
rect 10819 53319 10877 53320
rect 10923 53360 10965 53369
rect 10923 53320 10924 53360
rect 10964 53320 10965 53360
rect 10923 53311 10965 53320
rect 11115 53360 11157 53369
rect 11115 53320 11116 53360
rect 11156 53320 11157 53360
rect 11115 53311 11157 53320
rect 11299 53360 11357 53361
rect 11299 53320 11308 53360
rect 11348 53320 11357 53360
rect 11299 53319 11357 53320
rect 12547 53360 12605 53361
rect 12547 53320 12556 53360
rect 12596 53320 12605 53360
rect 12547 53319 12605 53320
rect 13131 53360 13173 53369
rect 13131 53320 13132 53360
rect 13172 53320 13173 53360
rect 13131 53311 13173 53320
rect 13227 53360 13269 53369
rect 13227 53320 13228 53360
rect 13268 53320 13269 53360
rect 13227 53311 13269 53320
rect 13611 53360 13653 53369
rect 13611 53320 13612 53360
rect 13652 53320 13653 53360
rect 13611 53311 13653 53320
rect 13707 53360 13749 53369
rect 13707 53320 13708 53360
rect 13748 53320 13749 53360
rect 13707 53311 13749 53320
rect 14179 53360 14237 53361
rect 14179 53320 14188 53360
rect 14228 53320 14237 53360
rect 15427 53360 15485 53361
rect 14179 53319 14237 53320
rect 14715 53350 14757 53359
rect 14715 53310 14716 53350
rect 14756 53310 14757 53350
rect 15427 53320 15436 53360
rect 15476 53320 15485 53360
rect 15427 53319 15485 53320
rect 16875 53360 16917 53369
rect 16875 53320 16876 53360
rect 16916 53320 16917 53360
rect 14715 53301 14757 53310
rect 16675 53318 16733 53319
rect 7275 53276 7317 53285
rect 16675 53278 16684 53318
rect 16724 53278 16733 53318
rect 16875 53311 16917 53320
rect 16971 53360 17013 53369
rect 16971 53320 16972 53360
rect 17012 53320 17013 53360
rect 16971 53311 17013 53320
rect 17067 53360 17109 53369
rect 17067 53320 17068 53360
rect 17108 53320 17109 53360
rect 17067 53311 17109 53320
rect 17163 53360 17205 53369
rect 17163 53320 17164 53360
rect 17204 53320 17205 53360
rect 17163 53311 17205 53320
rect 17547 53360 17589 53369
rect 17547 53320 17548 53360
rect 17588 53320 17589 53360
rect 17547 53311 17589 53320
rect 17643 53360 17685 53369
rect 17643 53320 17644 53360
rect 17684 53320 17685 53360
rect 17643 53311 17685 53320
rect 17739 53360 17781 53369
rect 17739 53320 17740 53360
rect 17780 53320 17781 53360
rect 17739 53311 17781 53320
rect 17835 53360 17877 53369
rect 17835 53320 17836 53360
rect 17876 53320 17877 53360
rect 17835 53311 17877 53320
rect 18019 53360 18077 53361
rect 18019 53320 18028 53360
rect 18068 53320 18077 53360
rect 18019 53319 18077 53320
rect 19267 53360 19325 53361
rect 19267 53320 19276 53360
rect 19316 53320 19325 53360
rect 19267 53319 19325 53320
rect 19659 53360 19701 53369
rect 19659 53320 19660 53360
rect 19700 53320 19701 53360
rect 19659 53311 19701 53320
rect 19851 53360 19893 53369
rect 19851 53320 19852 53360
rect 19892 53320 19893 53360
rect 19851 53311 19893 53320
rect 19939 53360 19997 53361
rect 19939 53320 19948 53360
rect 19988 53320 19997 53360
rect 19939 53319 19997 53320
rect 20227 53360 20285 53361
rect 20227 53320 20236 53360
rect 20276 53320 20285 53360
rect 20227 53319 20285 53320
rect 16675 53277 16733 53278
rect 7275 53236 7276 53276
rect 7316 53236 7317 53276
rect 7275 53227 7317 53236
rect 19467 53192 19509 53201
rect 19467 53152 19468 53192
rect 19508 53152 19509 53192
rect 19467 53143 19509 53152
rect 2667 53108 2709 53117
rect 2667 53068 2668 53108
rect 2708 53068 2709 53108
rect 2667 53059 2709 53068
rect 10443 53108 10485 53117
rect 10443 53068 10444 53108
rect 10484 53068 10485 53108
rect 10443 53059 10485 53068
rect 11115 53108 11157 53117
rect 11115 53068 11116 53108
rect 11156 53068 11157 53108
rect 11115 53059 11157 53068
rect 19659 53108 19701 53117
rect 19659 53068 19660 53108
rect 19700 53068 19701 53108
rect 19659 53059 19701 53068
rect 1152 52940 20352 52964
rect 1152 52900 3688 52940
rect 3728 52900 3770 52940
rect 3810 52900 3852 52940
rect 3892 52900 3934 52940
rect 3974 52900 4016 52940
rect 4056 52900 18808 52940
rect 18848 52900 18890 52940
rect 18930 52900 18972 52940
rect 19012 52900 19054 52940
rect 19094 52900 19136 52940
rect 19176 52900 20352 52940
rect 1152 52876 20352 52900
rect 11395 52772 11453 52773
rect 11395 52732 11404 52772
rect 11444 52732 11453 52772
rect 11395 52731 11453 52732
rect 16107 52772 16149 52781
rect 16107 52732 16108 52772
rect 16148 52732 16149 52772
rect 16107 52723 16149 52732
rect 18219 52772 18261 52781
rect 18219 52732 18220 52772
rect 18260 52732 18261 52772
rect 18219 52723 18261 52732
rect 3715 52688 3773 52689
rect 3715 52648 3724 52688
rect 3764 52648 3773 52688
rect 3715 52647 3773 52648
rect 12931 52688 12989 52689
rect 12931 52648 12940 52688
rect 12980 52648 12989 52688
rect 12931 52647 12989 52648
rect 17163 52688 17205 52697
rect 17163 52648 17164 52688
rect 17204 52648 17205 52688
rect 17163 52639 17205 52648
rect 11691 52604 11733 52613
rect 11691 52564 11692 52604
rect 11732 52564 11733 52604
rect 10339 52562 10397 52563
rect 6027 52533 6069 52542
rect 1411 52520 1469 52521
rect 1411 52480 1420 52520
rect 1460 52480 1469 52520
rect 1411 52479 1469 52480
rect 2659 52520 2717 52521
rect 2659 52480 2668 52520
rect 2708 52480 2717 52520
rect 2659 52479 2717 52480
rect 3051 52520 3093 52529
rect 3051 52480 3052 52520
rect 3092 52480 3093 52520
rect 3051 52471 3093 52480
rect 3339 52520 3381 52529
rect 3339 52480 3340 52520
rect 3380 52480 3381 52520
rect 3339 52471 3381 52480
rect 3531 52520 3573 52529
rect 3531 52480 3532 52520
rect 3572 52480 3573 52520
rect 3531 52471 3573 52480
rect 3723 52520 3765 52529
rect 3723 52480 3724 52520
rect 3764 52480 3765 52520
rect 3723 52471 3765 52480
rect 3819 52520 3861 52529
rect 3819 52480 3820 52520
rect 3860 52480 3861 52520
rect 3819 52471 3861 52480
rect 4195 52520 4253 52521
rect 4195 52480 4204 52520
rect 4244 52480 4253 52520
rect 4195 52479 4253 52480
rect 5443 52520 5501 52521
rect 5443 52480 5452 52520
rect 5492 52480 5501 52520
rect 5443 52479 5501 52480
rect 5835 52520 5877 52529
rect 5835 52480 5836 52520
rect 5876 52480 5877 52520
rect 6027 52493 6028 52533
rect 6068 52493 6069 52533
rect 6027 52484 6069 52493
rect 6219 52520 6261 52529
rect 5835 52471 5877 52480
rect 6219 52480 6220 52520
rect 6260 52480 6261 52520
rect 6219 52471 6261 52480
rect 6411 52520 6453 52529
rect 6411 52480 6412 52520
rect 6452 52480 6453 52520
rect 6411 52471 6453 52480
rect 6499 52520 6557 52521
rect 6499 52480 6508 52520
rect 6548 52480 6557 52520
rect 6499 52479 6557 52480
rect 6883 52520 6941 52521
rect 6883 52480 6892 52520
rect 6932 52480 6941 52520
rect 6883 52479 6941 52480
rect 8131 52520 8189 52521
rect 8131 52480 8140 52520
rect 8180 52480 8189 52520
rect 8131 52479 8189 52480
rect 8323 52520 8381 52521
rect 8323 52480 8332 52520
rect 8372 52480 8381 52520
rect 8323 52479 8381 52480
rect 9571 52520 9629 52521
rect 9571 52480 9580 52520
rect 9620 52480 9629 52520
rect 9571 52479 9629 52480
rect 10155 52520 10197 52529
rect 10155 52480 10156 52520
rect 10196 52480 10197 52520
rect 10155 52471 10197 52480
rect 10251 52520 10293 52529
rect 10339 52522 10348 52562
rect 10388 52522 10397 52562
rect 11691 52555 11733 52564
rect 16587 52604 16629 52613
rect 16587 52564 16588 52604
rect 16628 52564 16629 52604
rect 16587 52555 16629 52564
rect 20139 52565 20181 52574
rect 10339 52521 10397 52522
rect 10251 52480 10252 52520
rect 10292 52480 10293 52520
rect 10251 52471 10293 52480
rect 10731 52520 10773 52529
rect 10731 52480 10732 52520
rect 10772 52480 10773 52520
rect 10731 52471 10773 52480
rect 10827 52520 10869 52529
rect 10827 52480 10828 52520
rect 10868 52480 10869 52520
rect 10827 52471 10869 52480
rect 10923 52520 10965 52529
rect 10923 52480 10924 52520
rect 10964 52480 10965 52520
rect 10923 52471 10965 52480
rect 11203 52520 11261 52521
rect 11203 52480 11212 52520
rect 11252 52480 11261 52520
rect 11203 52479 11261 52480
rect 11595 52520 11637 52529
rect 11595 52480 11596 52520
rect 11636 52480 11637 52520
rect 11595 52471 11637 52480
rect 11787 52520 11829 52529
rect 11787 52480 11788 52520
rect 11828 52480 11829 52520
rect 11787 52471 11829 52480
rect 12459 52520 12501 52529
rect 12459 52480 12460 52520
rect 12500 52480 12501 52520
rect 12459 52471 12501 52480
rect 12555 52520 12597 52529
rect 12555 52480 12556 52520
rect 12596 52480 12597 52520
rect 12555 52471 12597 52480
rect 12747 52520 12789 52529
rect 12747 52480 12748 52520
rect 12788 52480 12789 52520
rect 12747 52471 12789 52480
rect 12939 52520 12981 52529
rect 12939 52480 12940 52520
rect 12980 52480 12981 52520
rect 12939 52471 12981 52480
rect 13035 52520 13077 52529
rect 13035 52480 13036 52520
rect 13076 52480 13077 52520
rect 13035 52471 13077 52480
rect 13219 52520 13277 52521
rect 13219 52480 13228 52520
rect 13268 52480 13277 52520
rect 13219 52479 13277 52480
rect 13315 52520 13373 52521
rect 13315 52480 13324 52520
rect 13364 52480 13373 52520
rect 13315 52479 13373 52480
rect 13515 52520 13557 52529
rect 13515 52480 13516 52520
rect 13556 52480 13557 52520
rect 13515 52471 13557 52480
rect 13611 52520 13653 52529
rect 13611 52480 13612 52520
rect 13652 52480 13653 52520
rect 13611 52471 13653 52480
rect 13704 52520 13762 52521
rect 13704 52480 13713 52520
rect 13753 52480 13762 52520
rect 13704 52479 13762 52480
rect 14187 52520 14229 52529
rect 14187 52480 14188 52520
rect 14228 52480 14229 52520
rect 14187 52471 14229 52480
rect 14275 52520 14333 52521
rect 14275 52480 14284 52520
rect 14324 52480 14333 52520
rect 14275 52479 14333 52480
rect 14659 52520 14717 52521
rect 14659 52480 14668 52520
rect 14708 52480 14717 52520
rect 14659 52479 14717 52480
rect 15907 52520 15965 52521
rect 15907 52480 15916 52520
rect 15956 52480 15965 52520
rect 15907 52479 15965 52480
rect 16491 52520 16533 52529
rect 16491 52480 16492 52520
rect 16532 52480 16533 52520
rect 16491 52471 16533 52480
rect 16683 52520 16725 52529
rect 16683 52480 16684 52520
rect 16724 52480 16725 52520
rect 16683 52471 16725 52480
rect 16875 52520 16917 52529
rect 16875 52480 16876 52520
rect 16916 52480 16917 52520
rect 16875 52471 16917 52480
rect 17163 52520 17205 52529
rect 17163 52480 17164 52520
rect 17204 52480 17205 52520
rect 17163 52471 17205 52480
rect 17355 52520 17397 52529
rect 17355 52480 17356 52520
rect 17396 52480 17397 52520
rect 17355 52471 17397 52480
rect 17547 52520 17589 52529
rect 17547 52480 17548 52520
rect 17588 52480 17589 52520
rect 17547 52471 17589 52480
rect 17643 52520 17685 52529
rect 17643 52480 17644 52520
rect 17684 52480 17685 52520
rect 17643 52471 17685 52480
rect 17835 52520 17877 52529
rect 17835 52480 17836 52520
rect 17876 52480 17877 52520
rect 17835 52471 17877 52480
rect 18027 52520 18069 52529
rect 18027 52480 18028 52520
rect 18068 52480 18069 52520
rect 18027 52471 18069 52480
rect 18403 52520 18461 52521
rect 18403 52480 18412 52520
rect 18452 52480 18461 52520
rect 18403 52479 18461 52480
rect 19651 52520 19709 52521
rect 19651 52480 19660 52520
rect 19700 52480 19709 52520
rect 19651 52479 19709 52480
rect 19851 52520 19893 52529
rect 19851 52480 19852 52520
rect 19892 52480 19893 52520
rect 19851 52471 19893 52480
rect 19947 52520 19989 52529
rect 19947 52480 19948 52520
rect 19988 52480 19989 52520
rect 19947 52471 19989 52480
rect 20043 52520 20085 52529
rect 20043 52480 20044 52520
rect 20084 52480 20085 52520
rect 20139 52525 20140 52565
rect 20180 52525 20181 52565
rect 20139 52516 20181 52525
rect 20043 52471 20085 52480
rect 5643 52436 5685 52445
rect 5643 52396 5644 52436
rect 5684 52396 5685 52436
rect 5643 52387 5685 52396
rect 6315 52436 6357 52445
rect 6315 52396 6316 52436
rect 6356 52396 6357 52436
rect 6315 52387 6357 52396
rect 17451 52436 17493 52445
rect 17451 52396 17452 52436
rect 17492 52396 17493 52436
rect 17451 52387 17493 52396
rect 2859 52352 2901 52361
rect 2859 52312 2860 52352
rect 2900 52312 2901 52352
rect 2859 52303 2901 52312
rect 3243 52352 3285 52361
rect 3243 52312 3244 52352
rect 3284 52312 3285 52352
rect 3243 52303 3285 52312
rect 5931 52352 5973 52361
rect 5931 52312 5932 52352
rect 5972 52312 5973 52352
rect 5931 52303 5973 52312
rect 6699 52352 6741 52361
rect 6699 52312 6700 52352
rect 6740 52312 6741 52352
rect 6699 52303 6741 52312
rect 9771 52352 9813 52361
rect 9771 52312 9772 52352
rect 9812 52312 9813 52352
rect 9771 52303 9813 52312
rect 10435 52352 10493 52353
rect 10435 52312 10444 52352
rect 10484 52312 10493 52352
rect 10435 52311 10493 52312
rect 10627 52352 10685 52353
rect 10627 52312 10636 52352
rect 10676 52312 10685 52352
rect 10627 52311 10685 52312
rect 11107 52352 11165 52353
rect 11107 52312 11116 52352
rect 11156 52312 11165 52352
rect 11107 52311 11165 52312
rect 12259 52352 12317 52353
rect 12259 52312 12268 52352
rect 12308 52312 12317 52352
rect 12259 52311 12317 52312
rect 13699 52352 13757 52353
rect 13699 52312 13708 52352
rect 13748 52312 13757 52352
rect 13699 52311 13757 52312
rect 17931 52352 17973 52361
rect 17931 52312 17932 52352
rect 17972 52312 17973 52352
rect 17931 52303 17973 52312
rect 1152 52184 20452 52208
rect 1152 52144 4928 52184
rect 4968 52144 5010 52184
rect 5050 52144 5092 52184
rect 5132 52144 5174 52184
rect 5214 52144 5256 52184
rect 5296 52144 20048 52184
rect 20088 52144 20130 52184
rect 20170 52144 20212 52184
rect 20252 52144 20294 52184
rect 20334 52144 20376 52184
rect 20416 52144 20452 52184
rect 1152 52120 20452 52144
rect 3051 52016 3093 52025
rect 3051 51976 3052 52016
rect 3092 51976 3093 52016
rect 3051 51967 3093 51976
rect 5451 52016 5493 52025
rect 5451 51976 5452 52016
rect 5492 51976 5493 52016
rect 5451 51967 5493 51976
rect 6603 52016 6645 52025
rect 6603 51976 6604 52016
rect 6644 51976 6645 52016
rect 6603 51967 6645 51976
rect 12939 52016 12981 52025
rect 12939 51976 12940 52016
rect 12980 51976 12981 52016
rect 12939 51967 12981 51976
rect 15819 52016 15861 52025
rect 15819 51976 15820 52016
rect 15860 51976 15861 52016
rect 15819 51967 15861 51976
rect 17931 52016 17973 52025
rect 17931 51976 17932 52016
rect 17972 51976 17973 52016
rect 17931 51967 17973 51976
rect 18404 51863 18462 51864
rect 1411 51848 1469 51849
rect 1411 51808 1420 51848
rect 1460 51808 1469 51848
rect 1411 51807 1469 51808
rect 2659 51848 2717 51849
rect 2659 51808 2668 51848
rect 2708 51808 2717 51848
rect 2659 51807 2717 51808
rect 3243 51843 3285 51852
rect 3243 51803 3244 51843
rect 3284 51803 3285 51843
rect 3715 51848 3773 51849
rect 3715 51808 3724 51848
rect 3764 51808 3773 51848
rect 3715 51807 3773 51808
rect 4203 51848 4245 51857
rect 4203 51808 4204 51848
rect 4244 51808 4245 51848
rect 3243 51794 3285 51803
rect 4203 51799 4245 51808
rect 4299 51848 4341 51857
rect 4299 51808 4300 51848
rect 4340 51808 4341 51848
rect 4299 51799 4341 51808
rect 4683 51848 4725 51857
rect 4683 51808 4684 51848
rect 4724 51808 4725 51848
rect 4683 51799 4725 51808
rect 4779 51848 4821 51857
rect 4779 51808 4780 51848
rect 4820 51808 4821 51848
rect 4779 51799 4821 51808
rect 5347 51848 5405 51849
rect 5347 51808 5356 51848
rect 5396 51808 5405 51848
rect 5347 51807 5405 51808
rect 5635 51848 5693 51849
rect 5635 51808 5644 51848
rect 5684 51808 5693 51848
rect 5635 51807 5693 51808
rect 5739 51848 5781 51857
rect 5739 51808 5740 51848
rect 5780 51808 5781 51848
rect 5739 51799 5781 51808
rect 5931 51848 5973 51857
rect 5931 51808 5932 51848
rect 5972 51808 5973 51848
rect 5931 51799 5973 51808
rect 6115 51848 6173 51849
rect 6115 51808 6124 51848
rect 6164 51808 6173 51848
rect 6115 51807 6173 51808
rect 6219 51848 6261 51857
rect 6219 51808 6220 51848
rect 6260 51808 6261 51848
rect 6219 51799 6261 51808
rect 6411 51848 6453 51857
rect 6411 51808 6412 51848
rect 6452 51808 6453 51848
rect 7267 51848 7325 51849
rect 6411 51799 6453 51808
rect 6747 51838 6789 51847
rect 6747 51798 6748 51838
rect 6788 51798 6789 51838
rect 7267 51808 7276 51848
rect 7316 51808 7325 51848
rect 7267 51807 7325 51808
rect 7755 51848 7797 51857
rect 7755 51808 7756 51848
rect 7796 51808 7797 51848
rect 7755 51799 7797 51808
rect 8235 51848 8277 51857
rect 8235 51808 8236 51848
rect 8276 51808 8277 51848
rect 8235 51799 8277 51808
rect 8331 51848 8373 51857
rect 8331 51808 8332 51848
rect 8372 51808 8373 51848
rect 8331 51799 8373 51808
rect 9859 51848 9917 51849
rect 9859 51808 9868 51848
rect 9908 51808 9917 51848
rect 9859 51807 9917 51808
rect 11107 51848 11165 51849
rect 11107 51808 11116 51848
rect 11156 51808 11165 51848
rect 11107 51807 11165 51808
rect 11491 51848 11549 51849
rect 11491 51808 11500 51848
rect 11540 51808 11549 51848
rect 11491 51807 11549 51808
rect 12739 51848 12797 51849
rect 12739 51808 12748 51848
rect 12788 51808 12797 51848
rect 12739 51807 12797 51808
rect 13507 51848 13565 51849
rect 13507 51808 13516 51848
rect 13556 51808 13565 51848
rect 13507 51807 13565 51808
rect 14755 51848 14813 51849
rect 14755 51808 14764 51848
rect 14804 51808 14813 51848
rect 14755 51807 14813 51808
rect 15907 51848 15965 51849
rect 15907 51808 15916 51848
rect 15956 51808 15965 51848
rect 15907 51807 15965 51808
rect 16203 51848 16245 51857
rect 16203 51808 16204 51848
rect 16244 51808 16245 51848
rect 16203 51799 16245 51808
rect 16299 51848 16341 51857
rect 16299 51808 16300 51848
rect 16340 51808 16341 51848
rect 16299 51799 16341 51808
rect 16683 51848 16725 51857
rect 16683 51808 16684 51848
rect 16724 51808 16725 51848
rect 16683 51799 16725 51808
rect 17251 51848 17309 51849
rect 17251 51808 17260 51848
rect 17300 51808 17309 51848
rect 18123 51848 18165 51857
rect 17251 51807 17309 51808
rect 17739 51834 17781 51843
rect 6747 51789 6789 51798
rect 17739 51794 17740 51834
rect 17780 51794 17781 51834
rect 18123 51808 18124 51848
rect 18164 51808 18165 51848
rect 18404 51823 18413 51863
rect 18453 51823 18462 51863
rect 18404 51822 18462 51823
rect 18691 51848 18749 51849
rect 18123 51799 18165 51808
rect 18691 51808 18700 51848
rect 18740 51808 18749 51848
rect 18691 51807 18749 51808
rect 19939 51848 19997 51849
rect 19939 51808 19948 51848
rect 19988 51808 19997 51848
rect 19939 51807 19997 51808
rect 17739 51785 17781 51794
rect 7851 51764 7893 51773
rect 7851 51724 7852 51764
rect 7892 51724 7893 51764
rect 7851 51715 7893 51724
rect 16779 51764 16821 51773
rect 16779 51724 16780 51764
rect 16820 51724 16821 51764
rect 16779 51715 16821 51724
rect 2859 51680 2901 51689
rect 2859 51640 2860 51680
rect 2900 51640 2901 51680
rect 2859 51631 2901 51640
rect 5931 51680 5973 51689
rect 5931 51640 5932 51680
rect 5972 51640 5973 51680
rect 5931 51631 5973 51640
rect 6411 51596 6453 51605
rect 6411 51556 6412 51596
rect 6452 51556 6453 51596
rect 6411 51547 6453 51556
rect 11307 51596 11349 51605
rect 11307 51556 11308 51596
rect 11348 51556 11349 51596
rect 11307 51547 11349 51556
rect 13323 51596 13365 51605
rect 13323 51556 13324 51596
rect 13364 51556 13365 51596
rect 13323 51547 13365 51556
rect 18123 51596 18165 51605
rect 18123 51556 18124 51596
rect 18164 51556 18165 51596
rect 18123 51547 18165 51556
rect 20139 51596 20181 51605
rect 20139 51556 20140 51596
rect 20180 51556 20181 51596
rect 20139 51547 20181 51556
rect 1152 51428 20352 51452
rect 1152 51388 3688 51428
rect 3728 51388 3770 51428
rect 3810 51388 3852 51428
rect 3892 51388 3934 51428
rect 3974 51388 4016 51428
rect 4056 51388 18808 51428
rect 18848 51388 18890 51428
rect 18930 51388 18972 51428
rect 19012 51388 19054 51428
rect 19094 51388 19136 51428
rect 19176 51388 20352 51428
rect 1152 51364 20352 51388
rect 6123 51260 6165 51269
rect 6123 51220 6124 51260
rect 6164 51220 6165 51260
rect 6123 51211 6165 51220
rect 12747 51260 12789 51269
rect 12747 51220 12748 51260
rect 12788 51220 12789 51260
rect 12747 51211 12789 51220
rect 3051 51176 3093 51185
rect 3051 51136 3052 51176
rect 3092 51136 3093 51176
rect 3051 51127 3093 51136
rect 18027 51176 18069 51185
rect 18027 51136 18028 51176
rect 18068 51136 18069 51176
rect 18027 51127 18069 51136
rect 3531 51092 3573 51101
rect 3531 51052 3532 51092
rect 3572 51052 3573 51092
rect 3531 51043 3573 51052
rect 8619 51092 8661 51101
rect 8619 51052 8620 51092
rect 8660 51052 8661 51092
rect 8619 51043 8661 51052
rect 14187 51092 14229 51101
rect 14187 51052 14188 51092
rect 14228 51052 14229 51092
rect 14187 51043 14229 51052
rect 19563 51092 19605 51101
rect 19563 51052 19564 51092
rect 19604 51052 19605 51092
rect 19563 51043 19605 51052
rect 9627 51017 9669 51026
rect 1219 51008 1277 51009
rect 1219 50968 1228 51008
rect 1268 50968 1277 51008
rect 1219 50967 1277 50968
rect 2467 51008 2525 51009
rect 2467 50968 2476 51008
rect 2516 50968 2525 51008
rect 2467 50967 2525 50968
rect 3051 51008 3093 51017
rect 3051 50968 3052 51008
rect 3092 50968 3093 51008
rect 3051 50959 3093 50968
rect 3339 51008 3381 51017
rect 3339 50968 3340 51008
rect 3380 50968 3381 51008
rect 3339 50959 3381 50968
rect 3627 51008 3669 51017
rect 3627 50968 3628 51008
rect 3668 50968 3669 51008
rect 3627 50959 3669 50968
rect 3819 51008 3861 51017
rect 3819 50968 3820 51008
rect 3860 50968 3861 51008
rect 3819 50959 3861 50968
rect 3915 51008 3957 51017
rect 3915 50968 3916 51008
rect 3956 50968 3957 51008
rect 3915 50959 3957 50968
rect 4011 51008 4053 51017
rect 4011 50968 4012 51008
rect 4052 50968 4053 51008
rect 4011 50959 4053 50968
rect 4107 51008 4149 51017
rect 4107 50968 4108 51008
rect 4148 50968 4149 51008
rect 4107 50959 4149 50968
rect 4675 51008 4733 51009
rect 4675 50968 4684 51008
rect 4724 50968 4733 51008
rect 4675 50967 4733 50968
rect 5923 51008 5981 51009
rect 5923 50968 5932 51008
rect 5972 50968 5981 51008
rect 5923 50967 5981 50968
rect 6307 51008 6365 51009
rect 6307 50968 6316 51008
rect 6356 50968 6365 51008
rect 6307 50967 6365 50968
rect 7555 51008 7613 51009
rect 7555 50968 7564 51008
rect 7604 50968 7613 51008
rect 7555 50967 7613 50968
rect 8043 51008 8085 51017
rect 8043 50968 8044 51008
rect 8084 50968 8085 51008
rect 8043 50959 8085 50968
rect 8139 51008 8181 51017
rect 8139 50968 8140 51008
rect 8180 50968 8181 51008
rect 8139 50959 8181 50968
rect 8523 51008 8565 51017
rect 8523 50968 8524 51008
rect 8564 50968 8565 51008
rect 8523 50959 8565 50968
rect 9091 51008 9149 51009
rect 9091 50968 9100 51008
rect 9140 50968 9149 51008
rect 9627 50977 9628 51017
rect 9668 50977 9669 51017
rect 13227 51022 13269 51031
rect 9627 50968 9669 50977
rect 11299 51008 11357 51009
rect 11299 50968 11308 51008
rect 11348 50968 11357 51008
rect 9091 50967 9149 50968
rect 11299 50967 11357 50968
rect 12547 51008 12605 51009
rect 12547 50968 12556 51008
rect 12596 50968 12605 51008
rect 13227 50982 13228 51022
rect 13268 50982 13269 51022
rect 18603 51022 18645 51031
rect 13227 50973 13269 50982
rect 13699 51008 13757 51009
rect 12547 50967 12605 50968
rect 13699 50968 13708 51008
rect 13748 50968 13757 51008
rect 13699 50967 13757 50968
rect 14283 51008 14325 51017
rect 14283 50968 14284 51008
rect 14324 50968 14325 51008
rect 14283 50959 14325 50968
rect 14667 51008 14709 51017
rect 14667 50968 14668 51008
rect 14708 50968 14709 51008
rect 14667 50959 14709 50968
rect 14763 51008 14805 51017
rect 14763 50968 14764 51008
rect 14804 50968 14805 51008
rect 14763 50959 14805 50968
rect 15523 51008 15581 51009
rect 15523 50968 15532 51008
rect 15572 50968 15581 51008
rect 15523 50967 15581 50968
rect 16771 51008 16829 51009
rect 16771 50968 16780 51008
rect 16820 50968 16829 51008
rect 16771 50967 16829 50968
rect 17355 51008 17397 51017
rect 17355 50968 17356 51008
rect 17396 50968 17397 51008
rect 17355 50959 17397 50968
rect 17547 51008 17589 51017
rect 17547 50968 17548 51008
rect 17588 50968 17589 51008
rect 17547 50959 17589 50968
rect 17635 51008 17693 51009
rect 17635 50968 17644 51008
rect 17684 50968 17693 51008
rect 17635 50967 17693 50968
rect 18027 51008 18069 51017
rect 18027 50968 18028 51008
rect 18068 50968 18069 51008
rect 18603 50982 18604 51022
rect 18644 50982 18645 51022
rect 18603 50973 18645 50982
rect 19075 51008 19133 51009
rect 18027 50959 18069 50968
rect 19075 50968 19084 51008
rect 19124 50968 19133 51008
rect 19075 50967 19133 50968
rect 19659 51008 19701 51017
rect 19659 50968 19660 51008
rect 19700 50968 19701 51008
rect 19659 50959 19701 50968
rect 20043 51008 20085 51017
rect 20043 50968 20044 51008
rect 20084 50968 20085 51008
rect 20043 50959 20085 50968
rect 20139 50988 20181 50997
rect 20139 50948 20140 50988
rect 20180 50948 20181 50988
rect 20139 50939 20181 50948
rect 7755 50924 7797 50933
rect 7755 50884 7756 50924
rect 7796 50884 7797 50924
rect 7755 50875 7797 50884
rect 13035 50924 13077 50933
rect 13035 50884 13036 50924
rect 13076 50884 13077 50924
rect 13035 50875 13077 50884
rect 18411 50924 18453 50933
rect 18411 50884 18412 50924
rect 18452 50884 18453 50924
rect 18411 50875 18453 50884
rect 2667 50840 2709 50849
rect 2667 50800 2668 50840
rect 2708 50800 2709 50840
rect 2667 50791 2709 50800
rect 2859 50840 2901 50849
rect 2859 50800 2860 50840
rect 2900 50800 2901 50840
rect 2859 50791 2901 50800
rect 9771 50840 9813 50849
rect 9771 50800 9772 50840
rect 9812 50800 9813 50840
rect 9771 50791 9813 50800
rect 16971 50840 17013 50849
rect 16971 50800 16972 50840
rect 17012 50800 17013 50840
rect 16971 50791 17013 50800
rect 17443 50840 17501 50841
rect 17443 50800 17452 50840
rect 17492 50800 17501 50840
rect 17443 50799 17501 50800
rect 17835 50840 17877 50849
rect 17835 50800 17836 50840
rect 17876 50800 17877 50840
rect 17835 50791 17877 50800
rect 1152 50672 20452 50696
rect 1152 50632 4928 50672
rect 4968 50632 5010 50672
rect 5050 50632 5092 50672
rect 5132 50632 5174 50672
rect 5214 50632 5256 50672
rect 5296 50632 20048 50672
rect 20088 50632 20130 50672
rect 20170 50632 20212 50672
rect 20252 50632 20294 50672
rect 20334 50632 20376 50672
rect 20416 50632 20452 50672
rect 1152 50608 20452 50632
rect 16971 50504 17013 50513
rect 16971 50464 16972 50504
rect 17012 50464 17013 50504
rect 16971 50455 17013 50464
rect 7947 50420 7989 50429
rect 7947 50380 7948 50420
rect 7988 50380 7989 50420
rect 7947 50371 7989 50380
rect 12651 50420 12693 50429
rect 12651 50380 12652 50420
rect 12692 50380 12693 50420
rect 12651 50371 12693 50380
rect 18987 50420 19029 50429
rect 18987 50380 18988 50420
rect 19028 50380 19029 50420
rect 18987 50371 19029 50380
rect 19275 50420 19317 50429
rect 19275 50380 19276 50420
rect 19316 50380 19317 50420
rect 19275 50371 19317 50380
rect 2563 50336 2621 50337
rect 2563 50296 2572 50336
rect 2612 50296 2621 50336
rect 2563 50295 2621 50296
rect 3811 50336 3869 50337
rect 3811 50296 3820 50336
rect 3860 50296 3869 50336
rect 3811 50295 3869 50296
rect 4099 50336 4157 50337
rect 4099 50296 4108 50336
rect 4148 50296 4157 50336
rect 4099 50295 4157 50296
rect 4579 50336 4637 50337
rect 4579 50296 4588 50336
rect 4628 50296 4637 50336
rect 4579 50295 4637 50296
rect 5827 50336 5885 50337
rect 5827 50296 5836 50336
rect 5876 50296 5885 50336
rect 5827 50295 5885 50296
rect 6403 50336 6461 50337
rect 6403 50296 6412 50336
rect 6452 50296 6461 50336
rect 6403 50295 6461 50296
rect 7363 50336 7421 50337
rect 7363 50296 7372 50336
rect 7412 50296 7421 50336
rect 7755 50336 7797 50345
rect 7363 50295 7421 50296
rect 7659 50291 7701 50300
rect 7659 50251 7660 50291
rect 7700 50251 7701 50291
rect 7755 50296 7756 50336
rect 7796 50296 7797 50336
rect 7755 50287 7797 50296
rect 7851 50336 7893 50345
rect 7851 50296 7852 50336
rect 7892 50296 7893 50336
rect 7851 50287 7893 50296
rect 8227 50336 8285 50337
rect 8227 50296 8236 50336
rect 8276 50296 8285 50336
rect 8227 50295 8285 50296
rect 9475 50336 9533 50337
rect 9475 50296 9484 50336
rect 9524 50296 9533 50336
rect 9475 50295 9533 50296
rect 11203 50336 11261 50337
rect 11203 50296 11212 50336
rect 11252 50296 11261 50336
rect 11203 50295 11261 50296
rect 12451 50336 12509 50337
rect 12451 50296 12460 50336
rect 12500 50296 12509 50336
rect 12451 50295 12509 50296
rect 13027 50336 13085 50337
rect 13027 50296 13036 50336
rect 13076 50296 13085 50336
rect 13027 50295 13085 50296
rect 14275 50336 14333 50337
rect 14275 50296 14284 50336
rect 14324 50296 14333 50336
rect 14275 50295 14333 50296
rect 15523 50336 15581 50337
rect 15523 50296 15532 50336
rect 15572 50296 15581 50336
rect 15523 50295 15581 50296
rect 16771 50336 16829 50337
rect 16771 50296 16780 50336
rect 16820 50296 16829 50336
rect 17355 50336 17397 50345
rect 16771 50295 16829 50296
rect 17163 50323 17205 50332
rect 17163 50283 17164 50323
rect 17204 50283 17205 50323
rect 17355 50296 17356 50336
rect 17396 50296 17397 50336
rect 17355 50287 17397 50296
rect 17539 50336 17597 50337
rect 17539 50296 17548 50336
rect 17588 50296 17597 50336
rect 17539 50295 17597 50296
rect 18787 50336 18845 50337
rect 18787 50296 18796 50336
rect 18836 50296 18845 50336
rect 18787 50295 18845 50296
rect 19179 50336 19221 50345
rect 19179 50296 19180 50336
rect 19220 50296 19221 50336
rect 19179 50287 19221 50296
rect 19371 50336 19413 50345
rect 19371 50296 19372 50336
rect 19412 50296 19413 50336
rect 19371 50287 19413 50296
rect 19459 50336 19517 50337
rect 19459 50296 19468 50336
rect 19508 50296 19517 50336
rect 19755 50336 19797 50345
rect 19459 50295 19517 50296
rect 19659 50291 19701 50300
rect 17163 50274 17205 50283
rect 7659 50242 7701 50251
rect 19659 50251 19660 50291
rect 19700 50251 19701 50291
rect 19755 50296 19756 50336
rect 19796 50296 19797 50336
rect 19755 50287 19797 50296
rect 19947 50336 19989 50345
rect 19947 50296 19948 50336
rect 19988 50296 19989 50336
rect 19843 50294 19901 50295
rect 19843 50254 19852 50294
rect 19892 50254 19901 50294
rect 19947 50287 19989 50296
rect 20139 50336 20181 50345
rect 20139 50296 20140 50336
rect 20180 50296 20181 50336
rect 20139 50287 20181 50296
rect 20227 50336 20285 50337
rect 20227 50296 20236 50336
rect 20276 50296 20285 50336
rect 20227 50295 20285 50296
rect 19843 50253 19901 50254
rect 19659 50242 19701 50251
rect 2379 50084 2421 50093
rect 2379 50044 2380 50084
rect 2420 50044 2421 50084
rect 2379 50035 2421 50044
rect 4011 50084 4053 50093
rect 4011 50044 4012 50084
rect 4052 50044 4053 50084
rect 4011 50035 4053 50044
rect 6027 50084 6069 50093
rect 6027 50044 6028 50084
rect 6068 50044 6069 50084
rect 6027 50035 6069 50044
rect 9675 50084 9717 50093
rect 9675 50044 9676 50084
rect 9716 50044 9717 50084
rect 9675 50035 9717 50044
rect 12843 50084 12885 50093
rect 12843 50044 12844 50084
rect 12884 50044 12885 50084
rect 12843 50035 12885 50044
rect 17163 50084 17205 50093
rect 17163 50044 17164 50084
rect 17204 50044 17205 50084
rect 17163 50035 17205 50044
rect 1152 49916 20352 49940
rect 1152 49876 3688 49916
rect 3728 49876 3770 49916
rect 3810 49876 3852 49916
rect 3892 49876 3934 49916
rect 3974 49876 4016 49916
rect 4056 49876 18808 49916
rect 18848 49876 18890 49916
rect 18930 49876 18972 49916
rect 19012 49876 19054 49916
rect 19094 49876 19136 49916
rect 19176 49876 20352 49916
rect 1152 49852 20352 49876
rect 7083 49748 7125 49757
rect 7083 49708 7084 49748
rect 7124 49708 7125 49748
rect 7083 49699 7125 49708
rect 7267 49748 7325 49749
rect 7267 49708 7276 49748
rect 7316 49708 7325 49748
rect 7267 49707 7325 49708
rect 8235 49748 8277 49757
rect 8235 49708 8236 49748
rect 8276 49708 8277 49748
rect 8235 49699 8277 49708
rect 15243 49748 15285 49757
rect 15243 49708 15244 49748
rect 15284 49708 15285 49748
rect 15243 49699 15285 49708
rect 16675 49748 16733 49749
rect 16675 49708 16684 49748
rect 16724 49708 16733 49748
rect 16675 49707 16733 49708
rect 18411 49748 18453 49757
rect 18411 49708 18412 49748
rect 18452 49708 18453 49748
rect 18411 49699 18453 49708
rect 3819 49580 3861 49589
rect 3819 49540 3820 49580
rect 3860 49540 3861 49580
rect 3819 49531 3861 49540
rect 3915 49580 3957 49589
rect 3915 49540 3916 49580
rect 3956 49540 3957 49580
rect 3915 49531 3957 49540
rect 10155 49580 10197 49589
rect 10155 49540 10156 49580
rect 10196 49540 10197 49580
rect 10155 49531 10197 49540
rect 13899 49580 13941 49589
rect 13899 49540 13900 49580
rect 13940 49540 13941 49580
rect 13899 49531 13941 49540
rect 2859 49510 2901 49519
rect 2859 49470 2860 49510
rect 2900 49470 2901 49510
rect 2859 49461 2901 49470
rect 3331 49496 3389 49497
rect 3331 49456 3340 49496
rect 3380 49456 3389 49496
rect 3331 49455 3389 49456
rect 4299 49496 4341 49505
rect 4299 49456 4300 49496
rect 4340 49456 4341 49496
rect 4299 49447 4341 49456
rect 4395 49496 4437 49505
rect 4395 49456 4396 49496
rect 4436 49456 4437 49496
rect 4395 49447 4437 49456
rect 4779 49496 4821 49505
rect 4779 49456 4780 49496
rect 4820 49456 4821 49496
rect 4779 49447 4821 49456
rect 4875 49496 4917 49505
rect 4875 49456 4876 49496
rect 4916 49456 4917 49496
rect 4875 49447 4917 49456
rect 4971 49496 5013 49505
rect 4971 49456 4972 49496
rect 5012 49456 5013 49496
rect 4971 49447 5013 49456
rect 5635 49496 5693 49497
rect 5635 49456 5644 49496
rect 5684 49456 5693 49496
rect 5635 49455 5693 49456
rect 6883 49496 6941 49497
rect 6883 49456 6892 49496
rect 6932 49456 6941 49496
rect 6883 49455 6941 49456
rect 7563 49496 7605 49505
rect 7563 49456 7564 49496
rect 7604 49456 7605 49496
rect 7563 49447 7605 49456
rect 7659 49496 7701 49505
rect 7659 49456 7660 49496
rect 7700 49456 7701 49496
rect 7659 49447 7701 49456
rect 7939 49496 7997 49497
rect 7939 49456 7948 49496
rect 7988 49456 7997 49496
rect 7939 49455 7997 49456
rect 8235 49496 8277 49505
rect 8235 49456 8236 49496
rect 8276 49456 8277 49496
rect 8235 49447 8277 49456
rect 8427 49496 8469 49505
rect 8427 49456 8428 49496
rect 8468 49456 8469 49496
rect 8427 49447 8469 49456
rect 9579 49496 9621 49505
rect 9579 49456 9580 49496
rect 9620 49456 9621 49496
rect 9579 49447 9621 49456
rect 9675 49496 9717 49505
rect 9675 49456 9676 49496
rect 9716 49456 9717 49496
rect 9675 49447 9717 49456
rect 10059 49496 10101 49505
rect 11115 49501 11157 49510
rect 10059 49456 10060 49496
rect 10100 49456 10101 49496
rect 10059 49447 10101 49456
rect 10627 49496 10685 49497
rect 10627 49456 10636 49496
rect 10676 49456 10685 49496
rect 10627 49455 10685 49456
rect 11115 49461 11116 49501
rect 11156 49461 11157 49501
rect 11115 49452 11157 49461
rect 12939 49501 12981 49510
rect 12939 49461 12940 49501
rect 12980 49461 12981 49501
rect 12939 49452 12981 49461
rect 13411 49496 13469 49497
rect 13411 49456 13420 49496
rect 13460 49456 13469 49496
rect 13411 49455 13469 49456
rect 13995 49496 14037 49505
rect 13995 49456 13996 49496
rect 14036 49456 14037 49496
rect 13995 49447 14037 49456
rect 14379 49496 14421 49505
rect 14379 49456 14380 49496
rect 14420 49456 14421 49496
rect 14379 49447 14421 49456
rect 14475 49496 14517 49505
rect 14475 49456 14476 49496
rect 14516 49456 14517 49496
rect 14475 49447 14517 49456
rect 15051 49496 15093 49505
rect 15051 49456 15052 49496
rect 15092 49456 15093 49496
rect 15051 49447 15093 49456
rect 15243 49496 15285 49505
rect 15243 49456 15244 49496
rect 15284 49456 15285 49496
rect 15243 49447 15285 49456
rect 15435 49496 15477 49505
rect 15435 49456 15436 49496
rect 15476 49456 15477 49496
rect 15435 49447 15477 49456
rect 15531 49496 15573 49505
rect 15531 49456 15532 49496
rect 15572 49456 15573 49496
rect 15531 49447 15573 49456
rect 15627 49496 15669 49505
rect 15627 49456 15628 49496
rect 15668 49456 15669 49496
rect 15627 49447 15669 49456
rect 15723 49496 15765 49505
rect 15723 49456 15724 49496
rect 15764 49456 15765 49496
rect 15723 49447 15765 49456
rect 16003 49496 16061 49497
rect 16003 49456 16012 49496
rect 16052 49456 16061 49496
rect 16003 49455 16061 49456
rect 16299 49496 16341 49505
rect 16299 49456 16300 49496
rect 16340 49456 16341 49496
rect 16299 49447 16341 49456
rect 16395 49496 16437 49505
rect 16395 49456 16396 49496
rect 16436 49456 16437 49496
rect 16395 49447 16437 49456
rect 16963 49496 17021 49497
rect 16963 49456 16972 49496
rect 17012 49456 17021 49496
rect 16963 49455 17021 49456
rect 18211 49496 18269 49497
rect 18211 49456 18220 49496
rect 18260 49456 18269 49496
rect 18211 49455 18269 49456
rect 18595 49496 18653 49497
rect 18595 49456 18604 49496
rect 18644 49456 18653 49496
rect 18595 49455 18653 49456
rect 19843 49496 19901 49497
rect 19843 49456 19852 49496
rect 19892 49456 19901 49496
rect 19843 49455 19901 49456
rect 2667 49412 2709 49421
rect 2667 49372 2668 49412
rect 2708 49372 2709 49412
rect 2667 49363 2709 49372
rect 11307 49412 11349 49421
rect 11307 49372 11308 49412
rect 11348 49372 11349 49412
rect 11307 49363 11349 49372
rect 4675 49328 4733 49329
rect 4675 49288 4684 49328
rect 4724 49288 4733 49328
rect 4675 49287 4733 49288
rect 12747 49328 12789 49337
rect 12747 49288 12748 49328
rect 12788 49288 12789 49328
rect 12747 49279 12789 49288
rect 18411 49328 18453 49337
rect 18411 49288 18412 49328
rect 18452 49288 18453 49328
rect 18411 49279 18453 49288
rect 20043 49328 20085 49337
rect 20043 49288 20044 49328
rect 20084 49288 20085 49328
rect 20043 49279 20085 49288
rect 1152 49160 20452 49184
rect 1152 49120 4928 49160
rect 4968 49120 5010 49160
rect 5050 49120 5092 49160
rect 5132 49120 5174 49160
rect 5214 49120 5256 49160
rect 5296 49120 20048 49160
rect 20088 49120 20130 49160
rect 20170 49120 20212 49160
rect 20252 49120 20294 49160
rect 20334 49120 20376 49160
rect 20416 49120 20452 49160
rect 1152 49096 20452 49120
rect 3627 48992 3669 49001
rect 3627 48952 3628 48992
rect 3668 48952 3669 48992
rect 3627 48943 3669 48952
rect 9483 48992 9525 49001
rect 9483 48952 9484 48992
rect 9524 48952 9525 48992
rect 9483 48943 9525 48952
rect 13131 48992 13173 49001
rect 13131 48952 13132 48992
rect 13172 48952 13173 48992
rect 13131 48943 13173 48952
rect 17163 48992 17205 49001
rect 17163 48952 17164 48992
rect 17204 48952 17205 48992
rect 17163 48943 17205 48952
rect 17347 48992 17405 48993
rect 17347 48952 17356 48992
rect 17396 48952 17405 48992
rect 17347 48951 17405 48952
rect 17835 48992 17877 49001
rect 17835 48952 17836 48992
rect 17876 48952 17877 48992
rect 17835 48943 17877 48952
rect 7467 48908 7509 48917
rect 7467 48868 7468 48908
rect 7508 48868 7509 48908
rect 7467 48859 7509 48868
rect 11499 48908 11541 48917
rect 11499 48868 11500 48908
rect 11540 48868 11541 48908
rect 11499 48859 11541 48868
rect 15147 48908 15189 48917
rect 15147 48868 15148 48908
rect 15188 48868 15189 48908
rect 15147 48859 15189 48868
rect 1315 48824 1373 48825
rect 1315 48784 1324 48824
rect 1364 48784 1373 48824
rect 1315 48783 1373 48784
rect 2563 48824 2621 48825
rect 2563 48784 2572 48824
rect 2612 48784 2621 48824
rect 2563 48783 2621 48784
rect 3139 48824 3197 48825
rect 3139 48784 3148 48824
rect 3188 48784 3197 48824
rect 3139 48783 3197 48784
rect 3243 48824 3285 48833
rect 3243 48784 3244 48824
rect 3284 48784 3285 48824
rect 3243 48775 3285 48784
rect 3435 48824 3477 48833
rect 3435 48784 3436 48824
rect 3476 48784 3477 48824
rect 4291 48824 4349 48825
rect 3435 48775 3477 48784
rect 3771 48814 3813 48823
rect 3771 48774 3772 48814
rect 3812 48774 3813 48814
rect 4291 48784 4300 48824
rect 4340 48784 4349 48824
rect 4291 48783 4349 48784
rect 4779 48824 4821 48833
rect 4779 48784 4780 48824
rect 4820 48784 4821 48824
rect 4779 48775 4821 48784
rect 4875 48824 4917 48833
rect 4875 48784 4876 48824
rect 4916 48784 4917 48824
rect 4875 48775 4917 48784
rect 5259 48824 5301 48833
rect 5259 48784 5260 48824
rect 5300 48784 5301 48824
rect 5259 48775 5301 48784
rect 5355 48824 5397 48833
rect 5355 48784 5356 48824
rect 5396 48784 5397 48824
rect 5355 48775 5397 48784
rect 5739 48824 5781 48833
rect 5739 48784 5740 48824
rect 5780 48784 5781 48824
rect 5739 48775 5781 48784
rect 5835 48824 5877 48833
rect 5835 48784 5836 48824
rect 5876 48784 5877 48824
rect 5835 48775 5877 48784
rect 6219 48824 6261 48833
rect 6219 48784 6220 48824
rect 6260 48784 6261 48824
rect 6219 48775 6261 48784
rect 6315 48824 6357 48833
rect 6315 48784 6316 48824
rect 6356 48784 6357 48824
rect 6315 48775 6357 48784
rect 6787 48824 6845 48825
rect 6787 48784 6796 48824
rect 6836 48784 6845 48824
rect 6787 48783 6845 48784
rect 7275 48819 7317 48828
rect 7275 48779 7276 48819
rect 7316 48779 7317 48819
rect 3771 48765 3813 48774
rect 7275 48770 7317 48779
rect 7659 48824 7701 48833
rect 7659 48784 7660 48824
rect 7700 48784 7701 48824
rect 7659 48775 7701 48784
rect 7851 48824 7893 48833
rect 7851 48784 7852 48824
rect 7892 48784 7893 48824
rect 7851 48775 7893 48784
rect 8035 48824 8093 48825
rect 8035 48784 8044 48824
rect 8084 48784 8093 48824
rect 8035 48783 8093 48784
rect 9283 48824 9341 48825
rect 9283 48784 9292 48824
rect 9332 48784 9341 48824
rect 9283 48783 9341 48784
rect 9771 48824 9813 48833
rect 9771 48784 9772 48824
rect 9812 48784 9813 48824
rect 9771 48775 9813 48784
rect 9867 48824 9909 48833
rect 9867 48784 9868 48824
rect 9908 48784 9909 48824
rect 9867 48775 9909 48784
rect 10251 48824 10293 48833
rect 10251 48784 10252 48824
rect 10292 48784 10293 48824
rect 10251 48775 10293 48784
rect 10347 48824 10389 48833
rect 10347 48784 10348 48824
rect 10388 48784 10389 48824
rect 10347 48775 10389 48784
rect 10819 48824 10877 48825
rect 10819 48784 10828 48824
rect 10868 48784 10877 48824
rect 11683 48824 11741 48825
rect 10819 48783 10877 48784
rect 11355 48814 11397 48823
rect 11355 48774 11356 48814
rect 11396 48774 11397 48814
rect 11683 48784 11692 48824
rect 11732 48784 11741 48824
rect 11683 48783 11741 48784
rect 12931 48824 12989 48825
rect 12931 48784 12940 48824
rect 12980 48784 12989 48824
rect 12931 48783 12989 48784
rect 13699 48824 13757 48825
rect 13699 48784 13708 48824
rect 13748 48784 13757 48824
rect 13699 48783 13757 48784
rect 14947 48824 15005 48825
rect 14947 48784 14956 48824
rect 14996 48784 15005 48824
rect 14947 48783 15005 48784
rect 15435 48824 15477 48833
rect 15435 48784 15436 48824
rect 15476 48784 15477 48824
rect 15435 48775 15477 48784
rect 15531 48824 15573 48833
rect 15531 48784 15532 48824
rect 15572 48784 15573 48824
rect 15531 48775 15573 48784
rect 16483 48824 16541 48825
rect 16483 48784 16492 48824
rect 16532 48784 16541 48824
rect 16483 48783 16541 48784
rect 16971 48819 17013 48828
rect 16971 48779 16972 48819
rect 17012 48779 17013 48819
rect 11355 48765 11397 48774
rect 16971 48770 17013 48779
rect 17451 48824 17493 48833
rect 17451 48784 17452 48824
rect 17492 48784 17493 48824
rect 17451 48775 17493 48784
rect 17547 48824 17589 48833
rect 17547 48784 17548 48824
rect 17588 48784 17589 48824
rect 17547 48775 17589 48784
rect 17643 48824 17685 48833
rect 17643 48784 17644 48824
rect 17684 48784 17685 48824
rect 17643 48775 17685 48784
rect 18027 48819 18069 48828
rect 18027 48779 18028 48819
rect 18068 48779 18069 48819
rect 18499 48824 18557 48825
rect 18499 48784 18508 48824
rect 18548 48784 18557 48824
rect 18499 48783 18557 48784
rect 18987 48824 19029 48833
rect 18987 48784 18988 48824
rect 19028 48784 19029 48824
rect 18027 48770 18069 48779
rect 18987 48775 19029 48784
rect 19083 48824 19125 48833
rect 19083 48784 19084 48824
rect 19124 48784 19125 48824
rect 19083 48775 19125 48784
rect 19467 48824 19509 48833
rect 19467 48784 19468 48824
rect 19508 48784 19509 48824
rect 19467 48775 19509 48784
rect 19563 48824 19605 48833
rect 19563 48784 19564 48824
rect 19604 48784 19605 48824
rect 19563 48775 19605 48784
rect 19851 48824 19893 48833
rect 19851 48784 19852 48824
rect 19892 48784 19893 48824
rect 19851 48775 19893 48784
rect 20043 48824 20085 48833
rect 20043 48784 20044 48824
rect 20084 48784 20085 48824
rect 20043 48775 20085 48784
rect 20131 48824 20189 48825
rect 20131 48784 20140 48824
rect 20180 48784 20189 48824
rect 20131 48783 20189 48784
rect 15915 48740 15957 48749
rect 15915 48700 15916 48740
rect 15956 48700 15957 48740
rect 15915 48691 15957 48700
rect 16011 48740 16053 48749
rect 16011 48700 16012 48740
rect 16052 48700 16053 48740
rect 16011 48691 16053 48700
rect 3435 48656 3477 48665
rect 3435 48616 3436 48656
rect 3476 48616 3477 48656
rect 3435 48607 3477 48616
rect 7659 48656 7701 48665
rect 7659 48616 7660 48656
rect 7700 48616 7701 48656
rect 7659 48607 7701 48616
rect 2763 48572 2805 48581
rect 2763 48532 2764 48572
rect 2804 48532 2805 48572
rect 2763 48523 2805 48532
rect 19851 48572 19893 48581
rect 19851 48532 19852 48572
rect 19892 48532 19893 48572
rect 19851 48523 19893 48532
rect 1152 48404 20352 48428
rect 1152 48364 3688 48404
rect 3728 48364 3770 48404
rect 3810 48364 3852 48404
rect 3892 48364 3934 48404
rect 3974 48364 4016 48404
rect 4056 48364 18808 48404
rect 18848 48364 18890 48404
rect 18930 48364 18972 48404
rect 19012 48364 19054 48404
rect 19094 48364 19136 48404
rect 19176 48364 20352 48404
rect 1152 48340 20352 48364
rect 3243 48236 3285 48245
rect 3243 48196 3244 48236
rect 3284 48196 3285 48236
rect 3243 48187 3285 48196
rect 11691 48236 11733 48245
rect 11691 48196 11692 48236
rect 11732 48196 11733 48236
rect 11691 48187 11733 48196
rect 16203 48236 16245 48245
rect 16203 48196 16204 48236
rect 16244 48196 16245 48236
rect 16203 48187 16245 48196
rect 18411 48236 18453 48245
rect 18411 48196 18412 48236
rect 18452 48196 18453 48236
rect 18411 48187 18453 48196
rect 20043 48236 20085 48245
rect 20043 48196 20044 48236
rect 20084 48196 20085 48236
rect 20043 48187 20085 48196
rect 6795 48152 6837 48161
rect 6795 48112 6796 48152
rect 6836 48112 6837 48152
rect 6795 48103 6837 48112
rect 13035 48068 13077 48077
rect 13035 48028 13036 48068
rect 13076 48028 13077 48068
rect 13035 48019 13077 48028
rect 13131 48068 13173 48077
rect 13131 48028 13132 48068
rect 13172 48028 13173 48068
rect 13131 48019 13173 48028
rect 1219 47984 1277 47985
rect 1219 47944 1228 47984
rect 1268 47944 1277 47984
rect 1219 47943 1277 47944
rect 2467 47984 2525 47985
rect 2467 47944 2476 47984
rect 2516 47944 2525 47984
rect 2467 47943 2525 47944
rect 2859 47984 2901 47993
rect 2859 47944 2860 47984
rect 2900 47944 2901 47984
rect 2859 47935 2901 47944
rect 3051 47984 3093 47993
rect 3051 47944 3052 47984
rect 3092 47944 3093 47984
rect 3051 47935 3093 47944
rect 3427 47984 3485 47985
rect 3427 47944 3436 47984
rect 3476 47944 3485 47984
rect 3427 47943 3485 47944
rect 4675 47984 4733 47985
rect 4675 47944 4684 47984
rect 4724 47944 4733 47984
rect 4675 47943 4733 47944
rect 5347 47984 5405 47985
rect 5347 47944 5356 47984
rect 5396 47944 5405 47984
rect 5347 47943 5405 47944
rect 6595 47984 6653 47985
rect 6595 47944 6604 47984
rect 6644 47944 6653 47984
rect 6595 47943 6653 47944
rect 6987 47984 7029 47993
rect 6987 47944 6988 47984
rect 7028 47944 7029 47984
rect 6987 47935 7029 47944
rect 7083 47984 7125 47993
rect 7083 47944 7084 47984
rect 7124 47944 7125 47984
rect 7083 47935 7125 47944
rect 7467 47984 7509 47993
rect 7467 47944 7468 47984
rect 7508 47944 7509 47984
rect 7467 47935 7509 47944
rect 7563 47984 7605 47993
rect 7563 47944 7564 47984
rect 7604 47944 7605 47984
rect 7563 47935 7605 47944
rect 7659 47984 7701 47993
rect 7659 47944 7660 47984
rect 7700 47944 7701 47984
rect 7659 47935 7701 47944
rect 7755 47984 7797 47993
rect 7755 47944 7756 47984
rect 7796 47944 7797 47984
rect 7755 47935 7797 47944
rect 8611 47984 8669 47985
rect 8611 47944 8620 47984
rect 8660 47944 8669 47984
rect 8611 47943 8669 47944
rect 9859 47984 9917 47985
rect 9859 47944 9868 47984
rect 9908 47944 9917 47984
rect 9859 47943 9917 47944
rect 10243 47984 10301 47985
rect 10243 47944 10252 47984
rect 10292 47944 10301 47984
rect 10243 47943 10301 47944
rect 11491 47984 11549 47985
rect 11491 47944 11500 47984
rect 11540 47944 11549 47984
rect 11491 47943 11549 47944
rect 12555 47984 12597 47993
rect 12555 47944 12556 47984
rect 12596 47944 12597 47984
rect 12555 47935 12597 47944
rect 12651 47984 12693 47993
rect 14091 47989 14133 47998
rect 12651 47944 12652 47984
rect 12692 47944 12693 47984
rect 12651 47935 12693 47944
rect 13603 47984 13661 47985
rect 13603 47944 13612 47984
rect 13652 47944 13661 47984
rect 13603 47943 13661 47944
rect 14091 47949 14092 47989
rect 14132 47949 14133 47989
rect 14091 47940 14133 47949
rect 14755 47984 14813 47985
rect 14755 47944 14764 47984
rect 14804 47944 14813 47984
rect 14755 47943 14813 47944
rect 16003 47984 16061 47985
rect 16003 47944 16012 47984
rect 16052 47944 16061 47984
rect 16003 47943 16061 47944
rect 16395 47984 16437 47993
rect 16395 47944 16396 47984
rect 16436 47944 16437 47984
rect 16395 47935 16437 47944
rect 16491 47984 16533 47993
rect 16491 47944 16492 47984
rect 16532 47944 16533 47984
rect 16491 47935 16533 47944
rect 16963 47984 17021 47985
rect 16963 47944 16972 47984
rect 17012 47944 17021 47984
rect 16963 47943 17021 47944
rect 18211 47984 18269 47985
rect 18211 47944 18220 47984
rect 18260 47944 18269 47984
rect 18211 47943 18269 47944
rect 18595 47984 18653 47985
rect 18595 47944 18604 47984
rect 18644 47944 18653 47984
rect 18595 47943 18653 47944
rect 19843 47984 19901 47985
rect 19843 47944 19852 47984
rect 19892 47944 19901 47984
rect 19843 47943 19901 47944
rect 14283 47900 14325 47909
rect 14283 47860 14284 47900
rect 14324 47860 14325 47900
rect 14283 47851 14325 47860
rect 2667 47816 2709 47825
rect 2667 47776 2668 47816
rect 2708 47776 2709 47816
rect 2667 47767 2709 47776
rect 2955 47816 2997 47825
rect 2955 47776 2956 47816
rect 2996 47776 2997 47816
rect 2955 47767 2997 47776
rect 7267 47816 7325 47817
rect 7267 47776 7276 47816
rect 7316 47776 7325 47816
rect 7267 47775 7325 47776
rect 10059 47816 10101 47825
rect 10059 47776 10060 47816
rect 10100 47776 10101 47816
rect 10059 47767 10101 47776
rect 16675 47816 16733 47817
rect 16675 47776 16684 47816
rect 16724 47776 16733 47816
rect 16675 47775 16733 47776
rect 1152 47648 20452 47672
rect 1152 47608 4928 47648
rect 4968 47608 5010 47648
rect 5050 47608 5092 47648
rect 5132 47608 5174 47648
rect 5214 47608 5256 47648
rect 5296 47608 20048 47648
rect 20088 47608 20130 47648
rect 20170 47608 20212 47648
rect 20252 47608 20294 47648
rect 20334 47608 20376 47648
rect 20416 47608 20452 47648
rect 1152 47584 20452 47608
rect 6403 47480 6461 47481
rect 6403 47440 6412 47480
rect 6452 47440 6461 47480
rect 6403 47439 6461 47440
rect 12363 47480 12405 47489
rect 12363 47440 12364 47480
rect 12404 47440 12405 47480
rect 12363 47431 12405 47440
rect 13995 47480 14037 47489
rect 13995 47440 13996 47480
rect 14036 47440 14037 47480
rect 13995 47431 14037 47440
rect 16395 47480 16437 47489
rect 16395 47440 16396 47480
rect 16436 47440 16437 47480
rect 16395 47431 16437 47440
rect 2571 47396 2613 47405
rect 2571 47356 2572 47396
rect 2612 47356 2613 47396
rect 2571 47347 2613 47356
rect 10347 47396 10389 47405
rect 10347 47356 10348 47396
rect 10388 47356 10389 47396
rect 10347 47347 10389 47356
rect 2475 47312 2517 47321
rect 2475 47272 2476 47312
rect 2516 47272 2517 47312
rect 2475 47263 2517 47272
rect 2667 47312 2709 47321
rect 2667 47272 2668 47312
rect 2708 47272 2709 47312
rect 2667 47263 2709 47272
rect 2755 47312 2813 47313
rect 2755 47272 2764 47312
rect 2804 47272 2813 47312
rect 2755 47271 2813 47272
rect 2947 47312 3005 47313
rect 2947 47272 2956 47312
rect 2996 47272 3005 47312
rect 2947 47271 3005 47272
rect 4195 47312 4253 47313
rect 4195 47272 4204 47312
rect 4244 47272 4253 47312
rect 4195 47271 4253 47272
rect 4587 47312 4629 47321
rect 4587 47272 4588 47312
rect 4628 47272 4629 47312
rect 4587 47263 4629 47272
rect 4875 47312 4917 47321
rect 4875 47272 4876 47312
rect 4916 47272 4917 47312
rect 4875 47263 4917 47272
rect 6603 47312 6645 47321
rect 6603 47272 6604 47312
rect 6644 47272 6645 47312
rect 6603 47263 6645 47272
rect 6699 47312 6741 47321
rect 6699 47272 6700 47312
rect 6740 47272 6741 47312
rect 6699 47263 6741 47272
rect 6883 47312 6941 47313
rect 6883 47272 6892 47312
rect 6932 47272 6941 47312
rect 6883 47271 6941 47272
rect 8131 47312 8189 47313
rect 8131 47272 8140 47312
rect 8180 47272 8189 47312
rect 8131 47271 8189 47272
rect 8619 47312 8661 47321
rect 8619 47272 8620 47312
rect 8660 47272 8661 47312
rect 8619 47263 8661 47272
rect 8715 47312 8757 47321
rect 8715 47272 8716 47312
rect 8756 47272 8757 47312
rect 8715 47263 8757 47272
rect 9667 47312 9725 47313
rect 9667 47272 9676 47312
rect 9716 47272 9725 47312
rect 9667 47271 9725 47272
rect 10155 47307 10197 47316
rect 10155 47267 10156 47307
rect 10196 47267 10197 47307
rect 10915 47312 10973 47313
rect 10915 47272 10924 47312
rect 10964 47272 10973 47312
rect 10915 47271 10973 47272
rect 12163 47312 12221 47313
rect 12163 47272 12172 47312
rect 12212 47272 12221 47312
rect 12163 47271 12221 47272
rect 12547 47312 12605 47313
rect 12547 47272 12556 47312
rect 12596 47272 12605 47312
rect 12547 47271 12605 47272
rect 13795 47312 13853 47313
rect 13795 47272 13804 47312
rect 13844 47272 13853 47312
rect 13795 47271 13853 47272
rect 14947 47312 15005 47313
rect 14947 47272 14956 47312
rect 14996 47272 15005 47312
rect 14947 47271 15005 47272
rect 16195 47312 16253 47313
rect 16195 47272 16204 47312
rect 16244 47272 16253 47312
rect 16195 47271 16253 47272
rect 16771 47312 16829 47313
rect 16771 47272 16780 47312
rect 16820 47272 16829 47312
rect 16771 47271 16829 47272
rect 18019 47312 18077 47313
rect 18019 47272 18028 47312
rect 18068 47272 18077 47312
rect 18019 47271 18077 47272
rect 18595 47312 18653 47313
rect 18595 47272 18604 47312
rect 18644 47272 18653 47312
rect 18595 47271 18653 47272
rect 19843 47312 19901 47313
rect 19843 47272 19852 47312
rect 19892 47272 19901 47312
rect 19843 47271 19901 47272
rect 10155 47258 10197 47267
rect 9099 47228 9141 47237
rect 9099 47188 9100 47228
rect 9140 47188 9141 47228
rect 9099 47179 9141 47188
rect 9195 47228 9237 47237
rect 9195 47188 9196 47228
rect 9236 47188 9237 47228
rect 9195 47179 9237 47188
rect 8331 47144 8373 47153
rect 8331 47104 8332 47144
rect 8372 47104 8373 47144
rect 8331 47095 8373 47104
rect 4395 47060 4437 47069
rect 4395 47020 4396 47060
rect 4436 47020 4437 47060
rect 4395 47011 4437 47020
rect 4587 47060 4629 47069
rect 4587 47020 4588 47060
rect 4628 47020 4629 47060
rect 4587 47011 4629 47020
rect 18219 47060 18261 47069
rect 18219 47020 18220 47060
rect 18260 47020 18261 47060
rect 18219 47011 18261 47020
rect 20043 47060 20085 47069
rect 20043 47020 20044 47060
rect 20084 47020 20085 47060
rect 20043 47011 20085 47020
rect 1152 46892 20352 46916
rect 1152 46852 3688 46892
rect 3728 46852 3770 46892
rect 3810 46852 3852 46892
rect 3892 46852 3934 46892
rect 3974 46852 4016 46892
rect 4056 46852 18808 46892
rect 18848 46852 18890 46892
rect 18930 46852 18972 46892
rect 19012 46852 19054 46892
rect 19094 46852 19136 46892
rect 19176 46852 20352 46892
rect 1152 46828 20352 46852
rect 3435 46556 3477 46565
rect 3435 46516 3436 46556
rect 3476 46516 3477 46556
rect 10731 46556 10773 46565
rect 3435 46507 3477 46516
rect 6123 46514 6165 46523
rect 10731 46516 10732 46556
rect 10772 46516 10773 46556
rect 4491 46486 4533 46495
rect 1219 46472 1277 46473
rect 1219 46432 1228 46472
rect 1268 46432 1277 46472
rect 1219 46431 1277 46432
rect 2467 46472 2525 46473
rect 2467 46432 2476 46472
rect 2516 46432 2525 46472
rect 2467 46431 2525 46432
rect 2955 46472 2997 46481
rect 2955 46432 2956 46472
rect 2996 46432 2997 46472
rect 2955 46423 2997 46432
rect 3051 46472 3093 46481
rect 3051 46432 3052 46472
rect 3092 46432 3093 46472
rect 3051 46423 3093 46432
rect 3531 46472 3573 46481
rect 3531 46432 3532 46472
rect 3572 46432 3573 46472
rect 3531 46423 3573 46432
rect 4003 46472 4061 46473
rect 4003 46432 4012 46472
rect 4052 46432 4061 46472
rect 4491 46446 4492 46486
rect 4532 46446 4533 46486
rect 4491 46437 4533 46446
rect 4971 46472 5013 46481
rect 4003 46431 4061 46432
rect 4971 46432 4972 46472
rect 5012 46432 5013 46472
rect 4971 46423 5013 46432
rect 5067 46472 5109 46481
rect 5067 46432 5068 46472
rect 5108 46432 5109 46472
rect 5067 46423 5109 46432
rect 5163 46472 5205 46481
rect 5163 46432 5164 46472
rect 5204 46432 5205 46472
rect 6123 46474 6124 46514
rect 6164 46474 6165 46514
rect 6123 46465 6165 46474
rect 6211 46514 6269 46515
rect 6211 46474 6220 46514
rect 6260 46474 6269 46514
rect 7267 46514 7325 46515
rect 6211 46473 6269 46474
rect 6315 46472 6357 46481
rect 5163 46423 5205 46432
rect 6315 46432 6316 46472
rect 6356 46432 6357 46472
rect 6315 46423 6357 46432
rect 6411 46472 6453 46481
rect 6411 46432 6412 46472
rect 6452 46432 6453 46472
rect 6411 46423 6453 46432
rect 6691 46472 6749 46473
rect 6691 46432 6700 46472
rect 6740 46432 6749 46472
rect 6691 46431 6749 46432
rect 7083 46472 7125 46481
rect 7083 46432 7084 46472
rect 7124 46432 7125 46472
rect 7083 46423 7125 46432
rect 7179 46472 7221 46481
rect 7267 46474 7276 46514
rect 7316 46474 7325 46514
rect 10731 46507 10773 46516
rect 13419 46556 13461 46565
rect 13419 46516 13420 46556
rect 13460 46516 13461 46556
rect 13419 46507 13461 46516
rect 19083 46556 19125 46565
rect 19083 46516 19084 46556
rect 19124 46516 19125 46556
rect 19083 46507 19125 46516
rect 7267 46473 7325 46474
rect 7179 46432 7180 46472
rect 7220 46432 7221 46472
rect 7179 46423 7221 46432
rect 7755 46472 7797 46481
rect 7755 46432 7756 46472
rect 7796 46432 7797 46472
rect 7755 46423 7797 46432
rect 7851 46472 7893 46481
rect 7851 46432 7852 46472
rect 7892 46432 7893 46472
rect 7851 46423 7893 46432
rect 8043 46472 8085 46481
rect 8043 46432 8044 46472
rect 8084 46432 8085 46472
rect 8043 46423 8085 46432
rect 8235 46472 8277 46481
rect 8235 46432 8236 46472
rect 8276 46432 8277 46472
rect 8235 46423 8277 46432
rect 8419 46472 8477 46473
rect 8419 46432 8428 46472
rect 8468 46432 8477 46472
rect 8419 46431 8477 46432
rect 9667 46472 9725 46473
rect 9667 46432 9676 46472
rect 9716 46432 9725 46472
rect 9667 46431 9725 46432
rect 10155 46472 10197 46481
rect 10155 46432 10156 46472
rect 10196 46432 10197 46472
rect 10155 46423 10197 46432
rect 10251 46472 10293 46481
rect 10251 46432 10252 46472
rect 10292 46432 10293 46472
rect 10251 46423 10293 46432
rect 10635 46472 10677 46481
rect 11691 46477 11733 46486
rect 10635 46432 10636 46472
rect 10676 46432 10677 46472
rect 10635 46423 10677 46432
rect 11203 46472 11261 46473
rect 11203 46432 11212 46472
rect 11252 46432 11261 46472
rect 11203 46431 11261 46432
rect 11691 46437 11692 46477
rect 11732 46437 11733 46477
rect 11691 46428 11733 46437
rect 12843 46472 12885 46481
rect 12843 46432 12844 46472
rect 12884 46432 12885 46472
rect 12843 46423 12885 46432
rect 12939 46472 12981 46481
rect 12939 46432 12940 46472
rect 12980 46432 12981 46472
rect 12939 46423 12981 46432
rect 13323 46472 13365 46481
rect 14379 46477 14421 46486
rect 13323 46432 13324 46472
rect 13364 46432 13365 46472
rect 13323 46423 13365 46432
rect 13891 46472 13949 46473
rect 13891 46432 13900 46472
rect 13940 46432 13949 46472
rect 13891 46431 13949 46432
rect 14379 46437 14380 46477
rect 14420 46437 14421 46477
rect 14379 46428 14421 46437
rect 15331 46472 15389 46473
rect 15331 46432 15340 46472
rect 15380 46432 15389 46472
rect 15331 46431 15389 46432
rect 16579 46472 16637 46473
rect 16579 46432 16588 46472
rect 16628 46432 16637 46472
rect 16579 46431 16637 46432
rect 16971 46472 17013 46481
rect 16971 46432 16972 46472
rect 17012 46432 17013 46472
rect 16971 46423 17013 46432
rect 17067 46472 17109 46481
rect 17067 46432 17068 46472
rect 17108 46432 17109 46472
rect 17067 46423 17109 46432
rect 17163 46472 17205 46481
rect 17163 46432 17164 46472
rect 17204 46432 17205 46472
rect 17163 46423 17205 46432
rect 18507 46472 18549 46481
rect 18507 46432 18508 46472
rect 18548 46432 18549 46472
rect 18507 46423 18549 46432
rect 18603 46472 18645 46481
rect 18603 46432 18604 46472
rect 18644 46432 18645 46472
rect 18603 46423 18645 46432
rect 18987 46472 19029 46481
rect 20043 46477 20085 46486
rect 18987 46432 18988 46472
rect 19028 46432 19029 46472
rect 18987 46423 19029 46432
rect 19555 46472 19613 46473
rect 19555 46432 19564 46472
rect 19604 46432 19613 46472
rect 19555 46431 19613 46432
rect 20043 46437 20044 46477
rect 20084 46437 20085 46477
rect 20043 46428 20085 46437
rect 2667 46388 2709 46397
rect 2667 46348 2668 46388
rect 2708 46348 2709 46388
rect 2667 46339 2709 46348
rect 9867 46388 9909 46397
rect 9867 46348 9868 46388
rect 9908 46348 9909 46388
rect 9867 46339 9909 46348
rect 14571 46388 14613 46397
rect 14571 46348 14572 46388
rect 14612 46348 14613 46388
rect 14571 46339 14613 46348
rect 20235 46388 20277 46397
rect 20235 46348 20236 46388
rect 20276 46348 20277 46388
rect 20235 46339 20277 46348
rect 4683 46304 4725 46313
rect 4683 46264 4684 46304
rect 4724 46264 4725 46304
rect 4683 46255 4725 46264
rect 4867 46304 4925 46305
rect 4867 46264 4876 46304
rect 4916 46264 4925 46304
rect 4867 46263 4925 46264
rect 6883 46304 6941 46305
rect 6883 46264 6892 46304
rect 6932 46264 6941 46304
rect 6883 46263 6941 46264
rect 7363 46304 7421 46305
rect 7363 46264 7372 46304
rect 7412 46264 7421 46304
rect 7363 46263 7421 46264
rect 7555 46304 7613 46305
rect 7555 46264 7564 46304
rect 7604 46264 7613 46304
rect 7555 46263 7613 46264
rect 8139 46304 8181 46313
rect 8139 46264 8140 46304
rect 8180 46264 8181 46304
rect 8139 46255 8181 46264
rect 11883 46304 11925 46313
rect 11883 46264 11884 46304
rect 11924 46264 11925 46304
rect 11883 46255 11925 46264
rect 16779 46304 16821 46313
rect 16779 46264 16780 46304
rect 16820 46264 16821 46304
rect 16779 46255 16821 46264
rect 17251 46304 17309 46305
rect 17251 46264 17260 46304
rect 17300 46264 17309 46304
rect 17251 46263 17309 46264
rect 6595 46238 6653 46239
rect 6595 46198 6604 46238
rect 6644 46198 6653 46238
rect 6595 46197 6653 46198
rect 1152 46136 20452 46160
rect 1152 46096 4928 46136
rect 4968 46096 5010 46136
rect 5050 46096 5092 46136
rect 5132 46096 5174 46136
rect 5214 46096 5256 46136
rect 5296 46096 20048 46136
rect 20088 46096 20130 46136
rect 20170 46096 20212 46136
rect 20252 46096 20294 46136
rect 20334 46096 20376 46136
rect 20416 46096 20452 46136
rect 1152 46072 20452 46096
rect 2859 45968 2901 45977
rect 2859 45928 2860 45968
rect 2900 45928 2901 45968
rect 2859 45919 2901 45928
rect 12651 45968 12693 45977
rect 12651 45928 12652 45968
rect 12692 45928 12693 45968
rect 12651 45919 12693 45928
rect 14283 45968 14325 45977
rect 14283 45928 14284 45968
rect 14324 45928 14325 45968
rect 14283 45919 14325 45928
rect 14467 45968 14525 45969
rect 14467 45928 14476 45968
rect 14516 45928 14525 45968
rect 14467 45927 14525 45928
rect 3339 45884 3381 45893
rect 3339 45844 3340 45884
rect 3380 45844 3381 45884
rect 3339 45835 3381 45844
rect 7563 45884 7605 45893
rect 7563 45844 7564 45884
rect 7604 45844 7605 45884
rect 7563 45835 7605 45844
rect 17259 45884 17301 45893
rect 17259 45844 17260 45884
rect 17300 45844 17301 45884
rect 17259 45835 17301 45844
rect 1411 45800 1469 45801
rect 1411 45760 1420 45800
rect 1460 45760 1469 45800
rect 1411 45759 1469 45760
rect 2659 45800 2717 45801
rect 2659 45760 2668 45800
rect 2708 45760 2717 45800
rect 4003 45800 4061 45801
rect 2659 45759 2717 45760
rect 3531 45786 3573 45795
rect 3531 45746 3532 45786
rect 3572 45746 3573 45786
rect 4003 45760 4012 45800
rect 4052 45760 4061 45800
rect 4003 45759 4061 45760
rect 4971 45800 5013 45809
rect 4971 45760 4972 45800
rect 5012 45760 5013 45800
rect 4971 45751 5013 45760
rect 5067 45800 5109 45809
rect 5067 45760 5068 45800
rect 5108 45760 5109 45800
rect 5067 45751 5109 45760
rect 5835 45800 5877 45809
rect 5835 45760 5836 45800
rect 5876 45760 5877 45800
rect 5835 45751 5877 45760
rect 5931 45800 5973 45809
rect 5931 45760 5932 45800
rect 5972 45760 5973 45800
rect 5931 45751 5973 45760
rect 6315 45800 6357 45809
rect 6315 45760 6316 45800
rect 6356 45760 6357 45800
rect 6315 45751 6357 45760
rect 6411 45800 6453 45809
rect 6411 45760 6412 45800
rect 6452 45760 6453 45800
rect 6411 45751 6453 45760
rect 6883 45800 6941 45801
rect 6883 45760 6892 45800
rect 6932 45760 6941 45800
rect 7939 45800 7997 45801
rect 6883 45759 6941 45760
rect 7371 45786 7413 45795
rect 3531 45737 3573 45746
rect 7371 45746 7372 45786
rect 7412 45746 7413 45786
rect 7939 45760 7948 45800
rect 7988 45760 7997 45800
rect 7939 45759 7997 45760
rect 9187 45800 9245 45801
rect 9187 45760 9196 45800
rect 9236 45760 9245 45800
rect 9187 45759 9245 45760
rect 9571 45800 9629 45801
rect 9571 45760 9580 45800
rect 9620 45760 9629 45800
rect 9571 45759 9629 45760
rect 10819 45800 10877 45801
rect 10819 45760 10828 45800
rect 10868 45760 10877 45800
rect 10819 45759 10877 45760
rect 11203 45800 11261 45801
rect 11203 45760 11212 45800
rect 11252 45760 11261 45800
rect 11203 45759 11261 45760
rect 12451 45800 12509 45801
rect 12451 45760 12460 45800
rect 12500 45760 12509 45800
rect 12451 45759 12509 45760
rect 12835 45800 12893 45801
rect 12835 45760 12844 45800
rect 12884 45760 12893 45800
rect 12835 45759 12893 45760
rect 14083 45800 14141 45801
rect 14083 45760 14092 45800
rect 14132 45760 14141 45800
rect 14083 45759 14141 45760
rect 14667 45800 14709 45809
rect 14667 45760 14668 45800
rect 14708 45760 14709 45800
rect 14667 45751 14709 45760
rect 14763 45800 14805 45809
rect 14763 45760 14764 45800
rect 14804 45760 14805 45800
rect 14763 45751 14805 45760
rect 15531 45800 15573 45809
rect 15531 45760 15532 45800
rect 15572 45760 15573 45800
rect 15531 45751 15573 45760
rect 15627 45800 15669 45809
rect 15627 45760 15628 45800
rect 15668 45760 15669 45800
rect 15627 45751 15669 45760
rect 16011 45800 16053 45809
rect 16011 45760 16012 45800
rect 16052 45760 16053 45800
rect 16011 45751 16053 45760
rect 16107 45800 16149 45809
rect 16107 45760 16108 45800
rect 16148 45760 16149 45800
rect 16107 45751 16149 45760
rect 16579 45800 16637 45801
rect 16579 45760 16588 45800
rect 16628 45760 16637 45800
rect 16579 45759 16637 45760
rect 17067 45795 17109 45804
rect 17067 45755 17068 45795
rect 17108 45755 17109 45795
rect 17067 45746 17109 45755
rect 17451 45800 17493 45809
rect 17451 45760 17452 45800
rect 17492 45760 17493 45800
rect 17451 45751 17493 45760
rect 17739 45800 17781 45809
rect 17739 45760 17740 45800
rect 17780 45760 17781 45800
rect 17739 45751 17781 45760
rect 17931 45800 17973 45809
rect 17931 45760 17932 45800
rect 17972 45760 17973 45800
rect 17931 45751 17973 45760
rect 18027 45800 18069 45809
rect 18027 45760 18028 45800
rect 18068 45760 18069 45800
rect 18027 45751 18069 45760
rect 18219 45800 18261 45809
rect 18219 45760 18220 45800
rect 18260 45760 18261 45800
rect 18219 45751 18261 45760
rect 18403 45800 18461 45801
rect 18403 45760 18412 45800
rect 18452 45760 18461 45800
rect 18403 45759 18461 45760
rect 19651 45800 19709 45801
rect 19651 45760 19660 45800
rect 19700 45760 19709 45800
rect 19651 45759 19709 45760
rect 7371 45737 7413 45746
rect 4491 45716 4533 45725
rect 4491 45676 4492 45716
rect 4532 45676 4533 45716
rect 4491 45667 4533 45676
rect 4587 45716 4629 45725
rect 4587 45676 4588 45716
rect 4628 45676 4629 45716
rect 4587 45667 4629 45676
rect 11019 45632 11061 45641
rect 11019 45592 11020 45632
rect 11060 45592 11061 45632
rect 11019 45583 11061 45592
rect 17923 45632 17981 45633
rect 17923 45592 17932 45632
rect 17972 45592 17981 45632
rect 17923 45591 17981 45592
rect 9387 45548 9429 45557
rect 9387 45508 9388 45548
rect 9428 45508 9429 45548
rect 9387 45499 9429 45508
rect 17739 45548 17781 45557
rect 17739 45508 17740 45548
rect 17780 45508 17781 45548
rect 17739 45499 17781 45508
rect 19851 45548 19893 45557
rect 19851 45508 19852 45548
rect 19892 45508 19893 45548
rect 19851 45499 19893 45508
rect 1152 45380 20352 45404
rect 1152 45340 3688 45380
rect 3728 45340 3770 45380
rect 3810 45340 3852 45380
rect 3892 45340 3934 45380
rect 3974 45340 4016 45380
rect 4056 45340 18808 45380
rect 18848 45340 18890 45380
rect 18930 45340 18972 45380
rect 19012 45340 19054 45380
rect 19094 45340 19136 45380
rect 19176 45340 20352 45380
rect 1152 45316 20352 45340
rect 3435 45212 3477 45221
rect 3435 45172 3436 45212
rect 3476 45172 3477 45212
rect 3435 45163 3477 45172
rect 6987 45212 7029 45221
rect 6987 45172 6988 45212
rect 7028 45172 7029 45212
rect 6987 45163 7029 45172
rect 4003 45128 4061 45129
rect 4003 45088 4012 45128
rect 4052 45088 4061 45128
rect 4003 45087 4061 45088
rect 4395 45128 4437 45137
rect 4395 45088 4396 45128
rect 4436 45088 4437 45128
rect 4395 45079 4437 45088
rect 9771 45044 9813 45053
rect 8763 45002 8805 45011
rect 1987 44960 2045 44961
rect 1987 44920 1996 44960
rect 2036 44920 2045 44960
rect 1987 44919 2045 44920
rect 3235 44960 3293 44961
rect 3235 44920 3244 44960
rect 3284 44920 3293 44960
rect 3235 44919 3293 44920
rect 3723 44960 3765 44969
rect 3723 44920 3724 44960
rect 3764 44920 3765 44960
rect 3723 44911 3765 44920
rect 3915 44960 3957 44969
rect 3915 44920 3916 44960
rect 3956 44920 3957 44960
rect 3915 44911 3957 44920
rect 4011 44960 4053 44969
rect 4011 44920 4012 44960
rect 4052 44920 4053 44960
rect 4011 44911 4053 44920
rect 4395 44952 4437 44961
rect 4395 44912 4396 44952
rect 4436 44912 4437 44952
rect 4395 44903 4437 44912
rect 4683 44960 4725 44969
rect 4683 44920 4684 44960
rect 4724 44920 4725 44960
rect 4683 44911 4725 44920
rect 4971 44960 5013 44969
rect 4971 44920 4972 44960
rect 5012 44920 5013 44960
rect 4971 44911 5013 44920
rect 5539 44960 5597 44961
rect 5539 44920 5548 44960
rect 5588 44920 5597 44960
rect 5539 44919 5597 44920
rect 6787 44960 6845 44961
rect 6787 44920 6796 44960
rect 6836 44920 6845 44960
rect 6787 44919 6845 44920
rect 7179 44960 7221 44969
rect 7179 44920 7180 44960
rect 7220 44920 7221 44960
rect 7179 44911 7221 44920
rect 7275 44960 7317 44969
rect 7275 44920 7276 44960
rect 7316 44920 7317 44960
rect 7275 44911 7317 44920
rect 7371 44960 7413 44969
rect 7371 44920 7372 44960
rect 7412 44920 7413 44960
rect 7371 44911 7413 44920
rect 7467 44960 7509 44969
rect 7467 44920 7468 44960
rect 7508 44920 7509 44960
rect 7467 44911 7509 44920
rect 7651 44960 7709 44961
rect 7651 44920 7660 44960
rect 7700 44920 7709 44960
rect 7651 44919 7709 44920
rect 7755 44960 7797 44969
rect 7755 44920 7756 44960
rect 7796 44920 7797 44960
rect 7755 44911 7797 44920
rect 7947 44960 7989 44969
rect 7947 44920 7948 44960
rect 7988 44920 7989 44960
rect 7947 44911 7989 44920
rect 8131 44960 8189 44961
rect 8131 44920 8140 44960
rect 8180 44920 8189 44960
rect 8131 44919 8189 44920
rect 8235 44960 8277 44969
rect 8235 44920 8236 44960
rect 8276 44920 8277 44960
rect 8763 44962 8764 45002
rect 8804 44962 8805 45002
rect 9771 45004 9772 45044
rect 9812 45004 9813 45044
rect 9771 44995 9813 45004
rect 9867 45044 9909 45053
rect 9867 45004 9868 45044
rect 9908 45004 9909 45044
rect 9867 44995 9909 45004
rect 13803 45044 13845 45053
rect 13803 45004 13804 45044
rect 13844 45004 13845 45044
rect 13803 44995 13845 45004
rect 13899 45044 13941 45053
rect 13899 45004 13900 45044
rect 13940 45004 13941 45044
rect 13899 44995 13941 45004
rect 18891 45044 18933 45053
rect 18891 45004 18892 45044
rect 18932 45004 18933 45044
rect 18891 44995 18933 45004
rect 18987 45044 19029 45053
rect 18987 45004 18988 45044
rect 19028 45004 19029 45044
rect 18987 44995 19029 45004
rect 19947 44974 19989 44983
rect 8763 44953 8805 44962
rect 9283 44960 9341 44961
rect 8235 44911 8277 44920
rect 9283 44920 9292 44960
rect 9332 44920 9341 44960
rect 9283 44919 9341 44920
rect 10251 44960 10293 44969
rect 10251 44920 10252 44960
rect 10292 44920 10293 44960
rect 10251 44911 10293 44920
rect 10347 44960 10389 44969
rect 10347 44920 10348 44960
rect 10388 44920 10389 44960
rect 10347 44911 10389 44920
rect 11395 44960 11453 44961
rect 11395 44920 11404 44960
rect 11444 44920 11453 44960
rect 11395 44919 11453 44920
rect 12643 44960 12701 44961
rect 12643 44920 12652 44960
rect 12692 44920 12701 44960
rect 12643 44919 12701 44920
rect 13323 44960 13365 44969
rect 13323 44920 13324 44960
rect 13364 44920 13365 44960
rect 13323 44911 13365 44920
rect 13419 44960 13461 44969
rect 14859 44965 14901 44974
rect 13419 44920 13420 44960
rect 13460 44920 13461 44960
rect 13419 44911 13461 44920
rect 14371 44960 14429 44961
rect 14371 44920 14380 44960
rect 14420 44920 14429 44960
rect 14371 44919 14429 44920
rect 14859 44925 14860 44965
rect 14900 44925 14901 44965
rect 14859 44916 14901 44925
rect 15243 44960 15285 44969
rect 15243 44920 15244 44960
rect 15284 44920 15285 44960
rect 15243 44911 15285 44920
rect 15435 44960 15477 44969
rect 15435 44920 15436 44960
rect 15476 44920 15477 44960
rect 15435 44911 15477 44920
rect 16675 44960 16733 44961
rect 16675 44920 16684 44960
rect 16724 44920 16733 44960
rect 16675 44919 16733 44920
rect 17923 44960 17981 44961
rect 17923 44920 17932 44960
rect 17972 44920 17981 44960
rect 17923 44919 17981 44920
rect 18411 44960 18453 44969
rect 18411 44920 18412 44960
rect 18452 44920 18453 44960
rect 18411 44911 18453 44920
rect 18507 44960 18549 44969
rect 18507 44920 18508 44960
rect 18548 44920 18549 44960
rect 18507 44911 18549 44920
rect 19459 44960 19517 44961
rect 19459 44920 19468 44960
rect 19508 44920 19517 44960
rect 19947 44934 19948 44974
rect 19988 44934 19989 44974
rect 19947 44925 19989 44934
rect 19459 44919 19517 44920
rect 8619 44876 8661 44885
rect 8619 44836 8620 44876
rect 8660 44836 8661 44876
rect 8619 44827 8661 44836
rect 4203 44792 4245 44801
rect 4203 44752 4204 44792
rect 4244 44752 4245 44792
rect 4203 44743 4245 44752
rect 4875 44792 4917 44801
rect 4875 44752 4876 44792
rect 4916 44752 4917 44792
rect 4875 44743 4917 44752
rect 7843 44792 7901 44793
rect 7843 44752 7852 44792
rect 7892 44752 7901 44792
rect 7843 44751 7901 44752
rect 12843 44792 12885 44801
rect 12843 44752 12844 44792
rect 12884 44752 12885 44792
rect 15339 44792 15381 44801
rect 12843 44743 12885 44752
rect 15051 44750 15093 44759
rect 15051 44710 15052 44750
rect 15092 44710 15093 44750
rect 15339 44752 15340 44792
rect 15380 44752 15381 44792
rect 15339 44743 15381 44752
rect 16291 44792 16349 44793
rect 16291 44752 16300 44792
rect 16340 44752 16349 44792
rect 16291 44751 16349 44752
rect 18123 44792 18165 44801
rect 18123 44752 18124 44792
rect 18164 44752 18165 44792
rect 18123 44743 18165 44752
rect 20139 44792 20181 44801
rect 20139 44752 20140 44792
rect 20180 44752 20181 44792
rect 20139 44743 20181 44752
rect 15051 44701 15093 44710
rect 1152 44624 20452 44648
rect 1152 44584 4928 44624
rect 4968 44584 5010 44624
rect 5050 44584 5092 44624
rect 5132 44584 5174 44624
rect 5214 44584 5256 44624
rect 5296 44584 20048 44624
rect 20088 44584 20130 44624
rect 20170 44584 20212 44624
rect 20252 44584 20294 44624
rect 20334 44584 20376 44624
rect 20416 44584 20452 44624
rect 1152 44560 20452 44584
rect 4587 44456 4629 44465
rect 4587 44416 4588 44456
rect 4628 44416 4629 44456
rect 4587 44407 4629 44416
rect 6315 44456 6357 44465
rect 6315 44416 6316 44456
rect 6356 44416 6357 44456
rect 6315 44407 6357 44416
rect 8331 44456 8373 44465
rect 8331 44416 8332 44456
rect 8372 44416 8373 44456
rect 8331 44407 8373 44416
rect 13603 44456 13661 44457
rect 13603 44416 13612 44456
rect 13652 44416 13661 44456
rect 13603 44415 13661 44416
rect 16107 44456 16149 44465
rect 16107 44416 16108 44456
rect 16148 44416 16149 44456
rect 16107 44407 16149 44416
rect 10347 44372 10389 44381
rect 10347 44332 10348 44372
rect 10388 44332 10389 44372
rect 10347 44323 10389 44332
rect 19947 44372 19989 44381
rect 19947 44332 19948 44372
rect 19988 44332 19989 44372
rect 19947 44323 19989 44332
rect 3139 44288 3197 44289
rect 3139 44248 3148 44288
rect 3188 44248 3197 44288
rect 3139 44247 3197 44248
rect 4387 44288 4445 44289
rect 4387 44248 4396 44288
rect 4436 44248 4445 44288
rect 4387 44247 4445 44248
rect 4867 44288 4925 44289
rect 4867 44248 4876 44288
rect 4916 44248 4925 44288
rect 4867 44247 4925 44248
rect 6115 44288 6173 44289
rect 6115 44248 6124 44288
rect 6164 44248 6173 44288
rect 6115 44247 6173 44248
rect 6883 44288 6941 44289
rect 6883 44248 6892 44288
rect 6932 44248 6941 44288
rect 6883 44247 6941 44248
rect 8131 44288 8189 44289
rect 8131 44248 8140 44288
rect 8180 44248 8189 44288
rect 8131 44247 8189 44248
rect 8619 44288 8661 44297
rect 8619 44248 8620 44288
rect 8660 44248 8661 44288
rect 8619 44239 8661 44248
rect 8715 44288 8757 44297
rect 8715 44248 8716 44288
rect 8756 44248 8757 44288
rect 8715 44239 8757 44248
rect 9099 44288 9141 44297
rect 9099 44248 9100 44288
rect 9140 44248 9141 44288
rect 9099 44239 9141 44248
rect 9195 44288 9237 44297
rect 9195 44248 9196 44288
rect 9236 44248 9237 44288
rect 9195 44239 9237 44248
rect 9667 44288 9725 44289
rect 9667 44248 9676 44288
rect 9716 44248 9725 44288
rect 11779 44288 11837 44289
rect 9667 44247 9725 44248
rect 10155 44274 10197 44283
rect 10155 44234 10156 44274
rect 10196 44234 10197 44274
rect 11779 44248 11788 44288
rect 11828 44248 11837 44288
rect 11779 44247 11837 44248
rect 11971 44288 12029 44289
rect 11971 44248 11980 44288
rect 12020 44248 12029 44288
rect 11971 44247 12029 44248
rect 13219 44288 13277 44289
rect 13219 44248 13228 44288
rect 13268 44248 13277 44288
rect 13219 44247 13277 44248
rect 13803 44288 13845 44297
rect 13803 44248 13804 44288
rect 13844 44248 13845 44288
rect 13803 44239 13845 44248
rect 13899 44288 13941 44297
rect 13899 44248 13900 44288
rect 13940 44248 13941 44288
rect 13899 44239 13941 44248
rect 14091 44288 14133 44297
rect 14091 44248 14092 44288
rect 14132 44248 14133 44288
rect 14091 44239 14133 44248
rect 14187 44288 14229 44297
rect 14187 44248 14188 44288
rect 14228 44248 14229 44288
rect 14187 44239 14229 44248
rect 14283 44288 14325 44297
rect 14283 44248 14284 44288
rect 14324 44248 14325 44288
rect 14283 44239 14325 44248
rect 14379 44288 14421 44297
rect 14379 44248 14380 44288
rect 14420 44248 14421 44288
rect 14379 44239 14421 44248
rect 14659 44288 14717 44289
rect 14659 44248 14668 44288
rect 14708 44248 14717 44288
rect 14659 44247 14717 44248
rect 15907 44288 15965 44289
rect 15907 44248 15916 44288
rect 15956 44248 15965 44288
rect 15907 44247 15965 44248
rect 16779 44288 16821 44297
rect 16779 44248 16780 44288
rect 16820 44248 16821 44288
rect 16779 44239 16821 44248
rect 17163 44288 17205 44297
rect 17163 44248 17164 44288
rect 17204 44248 17205 44288
rect 17163 44239 17205 44248
rect 17259 44288 17301 44297
rect 17259 44248 17260 44288
rect 17300 44248 17301 44288
rect 17259 44239 17301 44248
rect 17451 44288 17493 44297
rect 17451 44248 17452 44288
rect 17492 44248 17493 44288
rect 17451 44239 17493 44248
rect 18219 44288 18261 44297
rect 18219 44248 18220 44288
rect 18260 44248 18261 44288
rect 18219 44239 18261 44248
rect 18315 44288 18357 44297
rect 18315 44248 18316 44288
rect 18356 44248 18357 44288
rect 18315 44239 18357 44248
rect 18699 44288 18741 44297
rect 18699 44248 18700 44288
rect 18740 44248 18741 44288
rect 18699 44239 18741 44248
rect 18795 44288 18837 44297
rect 18795 44248 18796 44288
rect 18836 44248 18837 44288
rect 18795 44239 18837 44248
rect 19267 44288 19325 44289
rect 19267 44248 19276 44288
rect 19316 44248 19325 44288
rect 19267 44247 19325 44248
rect 19803 44278 19845 44287
rect 10155 44225 10197 44234
rect 19803 44238 19804 44278
rect 19844 44238 19845 44278
rect 19803 44229 19845 44238
rect 13419 44120 13461 44129
rect 13419 44080 13420 44120
rect 13460 44080 13461 44120
rect 13419 44071 13461 44080
rect 16299 44120 16341 44129
rect 16299 44080 16300 44120
rect 16340 44080 16341 44120
rect 16299 44071 16341 44080
rect 16779 44120 16821 44129
rect 16779 44080 16780 44120
rect 16820 44080 16821 44120
rect 16779 44071 16821 44080
rect 11691 44036 11733 44045
rect 11691 43996 11692 44036
rect 11732 43996 11733 44036
rect 11691 43987 11733 43996
rect 16587 44036 16629 44045
rect 16587 43996 16588 44036
rect 16628 43996 16629 44036
rect 16587 43987 16629 43996
rect 1152 43868 20352 43892
rect 1152 43828 3688 43868
rect 3728 43828 3770 43868
rect 3810 43828 3852 43868
rect 3892 43828 3934 43868
rect 3974 43828 4016 43868
rect 4056 43828 18808 43868
rect 18848 43828 18890 43868
rect 18930 43828 18972 43868
rect 19012 43828 19054 43868
rect 19094 43828 19136 43868
rect 19176 43828 20352 43868
rect 1152 43804 20352 43828
rect 6699 43700 6741 43709
rect 6699 43660 6700 43700
rect 6740 43660 6741 43700
rect 6699 43651 6741 43660
rect 8331 43700 8373 43709
rect 8331 43660 8332 43700
rect 8372 43660 8373 43700
rect 8331 43651 8373 43660
rect 10155 43700 10197 43709
rect 10155 43660 10156 43700
rect 10196 43660 10197 43700
rect 10155 43651 10197 43660
rect 16107 43700 16149 43709
rect 16107 43660 16108 43700
rect 16148 43660 16149 43700
rect 16107 43651 16149 43660
rect 18603 43700 18645 43709
rect 18603 43660 18604 43700
rect 18644 43660 18645 43700
rect 18603 43651 18645 43660
rect 5067 43616 5109 43625
rect 5067 43576 5068 43616
rect 5108 43576 5109 43616
rect 5067 43567 5109 43576
rect 3619 43448 3677 43449
rect 3619 43408 3628 43448
rect 3668 43408 3677 43448
rect 3619 43407 3677 43408
rect 4867 43448 4925 43449
rect 4867 43408 4876 43448
rect 4916 43408 4925 43448
rect 4867 43407 4925 43408
rect 5251 43448 5309 43449
rect 5251 43408 5260 43448
rect 5300 43408 5309 43448
rect 5251 43407 5309 43408
rect 6499 43448 6557 43449
rect 6499 43408 6508 43448
rect 6548 43408 6557 43448
rect 6499 43407 6557 43408
rect 6883 43448 6941 43449
rect 6883 43408 6892 43448
rect 6932 43408 6941 43448
rect 6883 43407 6941 43408
rect 8131 43448 8189 43449
rect 8131 43408 8140 43448
rect 8180 43408 8189 43448
rect 8131 43407 8189 43408
rect 8707 43448 8765 43449
rect 8707 43408 8716 43448
rect 8756 43408 8765 43448
rect 8707 43407 8765 43408
rect 9955 43448 10013 43449
rect 9955 43408 9964 43448
rect 10004 43408 10013 43448
rect 9955 43407 10013 43408
rect 11299 43448 11357 43449
rect 11299 43408 11308 43448
rect 11348 43408 11357 43448
rect 11299 43407 11357 43408
rect 12547 43448 12605 43449
rect 12547 43408 12556 43448
rect 12596 43408 12605 43448
rect 12547 43407 12605 43408
rect 13131 43448 13173 43457
rect 13131 43408 13132 43448
rect 13172 43408 13173 43448
rect 13323 43448 13365 43457
rect 13131 43399 13173 43408
rect 13227 43427 13269 43436
rect 13227 43387 13228 43427
rect 13268 43387 13269 43427
rect 13323 43408 13324 43448
rect 13364 43408 13365 43448
rect 13323 43399 13365 43408
rect 13419 43448 13461 43457
rect 13419 43408 13420 43448
rect 13460 43408 13461 43448
rect 13419 43399 13461 43408
rect 13699 43448 13757 43449
rect 13699 43408 13708 43448
rect 13748 43408 13757 43448
rect 13699 43407 13757 43408
rect 14091 43448 14133 43457
rect 14091 43408 14092 43448
rect 14132 43408 14133 43448
rect 14091 43399 14133 43408
rect 14187 43448 14229 43457
rect 14187 43408 14188 43448
rect 14228 43408 14229 43448
rect 14187 43399 14229 43408
rect 14283 43448 14325 43457
rect 14283 43408 14284 43448
rect 14324 43408 14325 43448
rect 14283 43399 14325 43408
rect 14659 43448 14717 43449
rect 14659 43408 14668 43448
rect 14708 43408 14717 43448
rect 14659 43407 14717 43408
rect 15907 43448 15965 43449
rect 15907 43408 15916 43448
rect 15956 43408 15965 43448
rect 15907 43407 15965 43408
rect 16587 43448 16629 43457
rect 16587 43408 16588 43448
rect 16628 43408 16629 43448
rect 16587 43399 16629 43408
rect 16779 43448 16821 43457
rect 16779 43408 16780 43448
rect 16820 43408 16821 43448
rect 16779 43399 16821 43408
rect 16867 43448 16925 43449
rect 16867 43408 16876 43448
rect 16916 43408 16925 43448
rect 16867 43407 16925 43408
rect 17155 43448 17213 43449
rect 17155 43408 17164 43448
rect 17204 43408 17213 43448
rect 17155 43407 17213 43408
rect 18403 43448 18461 43449
rect 18403 43408 18412 43448
rect 18452 43408 18461 43448
rect 18403 43407 18461 43408
rect 13227 43378 13269 43387
rect 12747 43280 12789 43289
rect 12747 43240 12748 43280
rect 12788 43240 12789 43280
rect 12747 43231 12789 43240
rect 13603 43280 13661 43281
rect 13603 43240 13612 43280
rect 13652 43240 13661 43280
rect 13603 43239 13661 43240
rect 13891 43280 13949 43281
rect 13891 43240 13900 43280
rect 13940 43240 13949 43280
rect 13891 43239 13949 43240
rect 14371 43280 14429 43281
rect 14371 43240 14380 43280
rect 14420 43240 14429 43280
rect 14371 43239 14429 43240
rect 16291 43280 16349 43281
rect 16291 43240 16300 43280
rect 16340 43240 16349 43280
rect 16291 43239 16349 43240
rect 16675 43280 16733 43281
rect 16675 43240 16684 43280
rect 16724 43240 16733 43280
rect 16675 43239 16733 43240
rect 18979 43280 19037 43281
rect 18979 43240 18988 43280
rect 19028 43240 19037 43280
rect 18979 43239 19037 43240
rect 1152 43112 20452 43136
rect 1152 43072 4928 43112
rect 4968 43072 5010 43112
rect 5050 43072 5092 43112
rect 5132 43072 5174 43112
rect 5214 43072 5256 43112
rect 5296 43072 20048 43112
rect 20088 43072 20130 43112
rect 20170 43072 20212 43112
rect 20252 43072 20294 43112
rect 20334 43072 20376 43112
rect 20416 43072 20452 43112
rect 1152 43048 20452 43072
rect 16291 42944 16349 42945
rect 16291 42904 16300 42944
rect 16340 42904 16349 42944
rect 16291 42903 16349 42904
rect 4875 42860 4917 42869
rect 4875 42820 4876 42860
rect 4916 42820 4917 42860
rect 4875 42811 4917 42820
rect 9579 42860 9621 42869
rect 9579 42820 9580 42860
rect 9620 42820 9621 42860
rect 9579 42811 9621 42820
rect 1411 42776 1469 42777
rect 1411 42736 1420 42776
rect 1460 42736 1469 42776
rect 1411 42735 1469 42736
rect 2659 42776 2717 42777
rect 2659 42736 2668 42776
rect 2708 42736 2717 42776
rect 2659 42735 2717 42736
rect 3147 42776 3189 42785
rect 3147 42736 3148 42776
rect 3188 42736 3189 42776
rect 3147 42727 3189 42736
rect 3243 42776 3285 42785
rect 3243 42736 3244 42776
rect 3284 42736 3285 42776
rect 3243 42727 3285 42736
rect 4195 42776 4253 42777
rect 4195 42736 4204 42776
rect 4244 42736 4253 42776
rect 5347 42776 5405 42777
rect 4195 42735 4253 42736
rect 4683 42762 4725 42771
rect 4683 42722 4684 42762
rect 4724 42722 4725 42762
rect 5347 42736 5356 42776
rect 5396 42736 5405 42776
rect 5347 42735 5405 42736
rect 6595 42776 6653 42777
rect 6595 42736 6604 42776
rect 6644 42736 6653 42776
rect 6595 42735 6653 42736
rect 6787 42776 6845 42777
rect 6787 42736 6796 42776
rect 6836 42736 6845 42776
rect 6787 42735 6845 42736
rect 8035 42776 8093 42777
rect 8035 42736 8044 42776
rect 8084 42736 8093 42776
rect 8035 42735 8093 42736
rect 10723 42776 10781 42777
rect 10723 42736 10732 42776
rect 10772 42736 10781 42776
rect 10723 42735 10781 42736
rect 11971 42776 12029 42777
rect 11971 42736 11980 42776
rect 12020 42736 12029 42776
rect 11971 42735 12029 42736
rect 12739 42776 12797 42777
rect 12739 42736 12748 42776
rect 12788 42736 12797 42776
rect 12739 42735 12797 42736
rect 13987 42776 14045 42777
rect 13987 42736 13996 42776
rect 14036 42736 14045 42776
rect 13987 42735 14045 42736
rect 14659 42776 14717 42777
rect 14659 42736 14668 42776
rect 14708 42736 14717 42776
rect 14659 42735 14717 42736
rect 15907 42776 15965 42777
rect 15907 42736 15916 42776
rect 15956 42736 15965 42776
rect 15907 42735 15965 42736
rect 4683 42713 4725 42722
rect 3627 42692 3669 42701
rect 3627 42652 3628 42692
rect 3668 42652 3669 42692
rect 3627 42643 3669 42652
rect 3723 42692 3765 42701
rect 3723 42652 3724 42692
rect 3764 42652 3765 42692
rect 3723 42643 3765 42652
rect 9099 42692 9141 42701
rect 9099 42652 9100 42692
rect 9140 42652 9141 42692
rect 9099 42643 9141 42652
rect 20035 42692 20093 42693
rect 20035 42652 20044 42692
rect 20084 42652 20093 42692
rect 20035 42651 20093 42652
rect 16395 42608 16437 42617
rect 16395 42568 16396 42608
rect 16436 42568 16437 42608
rect 16395 42559 16437 42568
rect 17259 42608 17301 42617
rect 17259 42568 17260 42608
rect 17300 42568 17301 42608
rect 17259 42559 17301 42568
rect 18987 42608 19029 42617
rect 18987 42568 18988 42608
rect 19028 42568 19029 42608
rect 18987 42559 19029 42568
rect 19755 42608 19797 42617
rect 19755 42568 19756 42608
rect 19796 42568 19797 42608
rect 19755 42559 19797 42568
rect 20235 42608 20277 42617
rect 20235 42568 20236 42608
rect 20276 42568 20277 42608
rect 20235 42559 20277 42568
rect 2859 42524 2901 42533
rect 2859 42484 2860 42524
rect 2900 42484 2901 42524
rect 2859 42475 2901 42484
rect 5163 42524 5205 42533
rect 5163 42484 5164 42524
rect 5204 42484 5205 42524
rect 5163 42475 5205 42484
rect 8235 42524 8277 42533
rect 8235 42484 8236 42524
rect 8276 42484 8277 42524
rect 8235 42475 8277 42484
rect 12171 42524 12213 42533
rect 12171 42484 12172 42524
rect 12212 42484 12213 42524
rect 12171 42475 12213 42484
rect 14187 42524 14229 42533
rect 14187 42484 14188 42524
rect 14228 42484 14229 42524
rect 14187 42475 14229 42484
rect 16107 42524 16149 42533
rect 16107 42484 16108 42524
rect 16148 42484 16149 42524
rect 16107 42475 16149 42484
rect 1152 42356 20352 42380
rect 1152 42316 3688 42356
rect 3728 42316 3770 42356
rect 3810 42316 3852 42356
rect 3892 42316 3934 42356
rect 3974 42316 4016 42356
rect 4056 42316 18808 42356
rect 18848 42316 18890 42356
rect 18930 42316 18972 42356
rect 19012 42316 19054 42356
rect 19094 42316 19136 42356
rect 19176 42316 20352 42356
rect 1152 42292 20352 42316
rect 3915 42188 3957 42197
rect 3915 42148 3916 42188
rect 3956 42148 3957 42188
rect 3915 42139 3957 42148
rect 18123 42188 18165 42197
rect 18123 42148 18124 42188
rect 18164 42148 18165 42188
rect 18123 42139 18165 42148
rect 9099 42104 9141 42113
rect 9099 42064 9100 42104
rect 9140 42064 9141 42104
rect 9099 42055 9141 42064
rect 19851 42104 19893 42113
rect 19851 42064 19852 42104
rect 19892 42064 19893 42104
rect 19851 42055 19893 42064
rect 4779 42020 4821 42029
rect 4779 41980 4780 42020
rect 4820 41980 4821 42020
rect 4779 41971 4821 41980
rect 10251 42020 10293 42029
rect 10251 41980 10252 42020
rect 10292 41980 10293 42020
rect 10251 41971 10293 41980
rect 12843 42020 12885 42029
rect 12843 41980 12844 42020
rect 12884 41980 12885 42020
rect 12843 41971 12885 41980
rect 14955 42020 14997 42029
rect 14955 41980 14956 42020
rect 14996 41980 14997 42020
rect 17923 42020 17981 42021
rect 14955 41971 14997 41980
rect 15963 41978 16005 41987
rect 17923 41980 17932 42020
rect 17972 41980 17981 42020
rect 17923 41979 17981 41980
rect 19267 42020 19325 42021
rect 19267 41980 19276 42020
rect 19316 41980 19325 42020
rect 19267 41979 19325 41980
rect 19651 42020 19709 42021
rect 19651 41980 19660 42020
rect 19700 41980 19709 42020
rect 19651 41979 19709 41980
rect 5739 41950 5781 41959
rect 2467 41936 2525 41937
rect 2467 41896 2476 41936
rect 2516 41896 2525 41936
rect 2467 41895 2525 41896
rect 3715 41936 3773 41937
rect 3715 41896 3724 41936
rect 3764 41896 3773 41936
rect 3715 41895 3773 41896
rect 4203 41936 4245 41945
rect 4203 41896 4204 41936
rect 4244 41896 4245 41936
rect 4203 41887 4245 41896
rect 4299 41936 4341 41945
rect 4299 41896 4300 41936
rect 4340 41896 4341 41936
rect 4299 41887 4341 41896
rect 4683 41936 4725 41945
rect 4683 41896 4684 41936
rect 4724 41896 4725 41936
rect 4683 41887 4725 41896
rect 5251 41936 5309 41937
rect 5251 41896 5260 41936
rect 5300 41896 5309 41936
rect 5739 41910 5740 41950
rect 5780 41910 5781 41950
rect 5739 41901 5781 41910
rect 7363 41936 7421 41937
rect 5251 41895 5309 41896
rect 7363 41896 7372 41936
rect 7412 41896 7421 41936
rect 7363 41895 7421 41896
rect 8611 41936 8669 41937
rect 8611 41896 8620 41936
rect 8660 41896 8669 41936
rect 8611 41895 8669 41896
rect 9675 41936 9717 41945
rect 9675 41896 9676 41936
rect 9716 41896 9717 41936
rect 9675 41887 9717 41896
rect 9771 41936 9813 41945
rect 9771 41896 9772 41936
rect 9812 41896 9813 41936
rect 9771 41887 9813 41896
rect 10155 41936 10197 41945
rect 11211 41941 11253 41950
rect 10155 41896 10156 41936
rect 10196 41896 10197 41936
rect 10155 41887 10197 41896
rect 10723 41936 10781 41937
rect 10723 41896 10732 41936
rect 10772 41896 10781 41936
rect 10723 41895 10781 41896
rect 11211 41901 11212 41941
rect 11252 41901 11253 41941
rect 11211 41892 11253 41901
rect 12267 41936 12309 41945
rect 12267 41896 12268 41936
rect 12308 41896 12309 41936
rect 12267 41887 12309 41896
rect 12363 41936 12405 41945
rect 12363 41896 12364 41936
rect 12404 41896 12405 41936
rect 12363 41887 12405 41896
rect 12747 41936 12789 41945
rect 13803 41941 13845 41950
rect 12747 41896 12748 41936
rect 12788 41896 12789 41936
rect 12747 41887 12789 41896
rect 13315 41936 13373 41937
rect 13315 41896 13324 41936
rect 13364 41896 13373 41936
rect 13315 41895 13373 41896
rect 13803 41901 13804 41941
rect 13844 41901 13845 41941
rect 13803 41892 13845 41901
rect 14379 41936 14421 41945
rect 14379 41896 14380 41936
rect 14420 41896 14421 41936
rect 14379 41887 14421 41896
rect 14475 41936 14517 41945
rect 14475 41896 14476 41936
rect 14516 41896 14517 41936
rect 14475 41887 14517 41896
rect 14859 41936 14901 41945
rect 15963 41938 15964 41978
rect 16004 41938 16005 41978
rect 14859 41896 14860 41936
rect 14900 41896 14901 41936
rect 14859 41887 14901 41896
rect 15427 41936 15485 41937
rect 15427 41896 15436 41936
rect 15476 41896 15485 41936
rect 15963 41929 16005 41938
rect 16483 41936 16541 41937
rect 15427 41895 15485 41896
rect 16483 41896 16492 41936
rect 16532 41896 16541 41936
rect 16483 41895 16541 41896
rect 17731 41936 17789 41937
rect 17731 41896 17740 41936
rect 17780 41896 17789 41936
rect 17731 41895 17789 41896
rect 18987 41936 19029 41945
rect 18987 41896 18988 41936
rect 19028 41896 19029 41936
rect 18987 41887 19029 41896
rect 8811 41852 8853 41861
rect 8811 41812 8812 41852
rect 8852 41812 8853 41852
rect 8811 41803 8853 41812
rect 5931 41768 5973 41777
rect 5931 41728 5932 41768
rect 5972 41728 5973 41768
rect 5931 41719 5973 41728
rect 11403 41768 11445 41777
rect 11403 41728 11404 41768
rect 11444 41728 11445 41768
rect 11403 41719 11445 41728
rect 13995 41768 14037 41777
rect 13995 41728 13996 41768
rect 14036 41728 14037 41768
rect 13995 41719 14037 41728
rect 16107 41768 16149 41777
rect 16107 41728 16108 41768
rect 16148 41728 16149 41768
rect 16107 41719 16149 41728
rect 16299 41768 16341 41777
rect 16299 41728 16300 41768
rect 16340 41728 16341 41768
rect 16299 41719 16341 41728
rect 19467 41768 19509 41777
rect 19467 41728 19468 41768
rect 19508 41728 19509 41768
rect 19467 41719 19509 41728
rect 1152 41600 20452 41624
rect 1152 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20452 41600
rect 1152 41536 20452 41560
rect 3243 41432 3285 41441
rect 3243 41392 3244 41432
rect 3284 41392 3285 41432
rect 3243 41383 3285 41392
rect 11787 41432 11829 41441
rect 11787 41392 11788 41432
rect 11828 41392 11829 41432
rect 11787 41383 11829 41392
rect 13419 41432 13461 41441
rect 13419 41392 13420 41432
rect 13460 41392 13461 41432
rect 13419 41383 13461 41392
rect 16395 41432 16437 41441
rect 16395 41392 16396 41432
rect 16436 41392 16437 41432
rect 16395 41383 16437 41392
rect 18979 41432 19037 41433
rect 18979 41392 18988 41432
rect 19028 41392 19037 41432
rect 18979 41391 19037 41392
rect 19851 41432 19893 41441
rect 19851 41392 19852 41432
rect 19892 41392 19893 41432
rect 19851 41383 19893 41392
rect 5451 41348 5493 41357
rect 5451 41308 5452 41348
rect 5492 41308 5493 41348
rect 5451 41299 5493 41308
rect 8235 41348 8277 41357
rect 8235 41308 8236 41348
rect 8276 41308 8277 41348
rect 8235 41299 8277 41308
rect 10251 41348 10293 41357
rect 10251 41308 10252 41348
rect 10292 41308 10293 41348
rect 10251 41299 10293 41308
rect 16107 41348 16149 41357
rect 16107 41308 16108 41348
rect 16148 41308 16149 41348
rect 16107 41299 16149 41308
rect 1795 41264 1853 41265
rect 1795 41224 1804 41264
rect 1844 41224 1853 41264
rect 1795 41223 1853 41224
rect 3043 41264 3101 41265
rect 3043 41224 3052 41264
rect 3092 41224 3101 41264
rect 3043 41223 3101 41224
rect 3723 41264 3765 41273
rect 3723 41224 3724 41264
rect 3764 41224 3765 41264
rect 3723 41215 3765 41224
rect 3819 41264 3861 41273
rect 3819 41224 3820 41264
rect 3860 41224 3861 41264
rect 3819 41215 3861 41224
rect 4299 41264 4341 41273
rect 4299 41224 4300 41264
rect 4340 41224 4341 41264
rect 4299 41215 4341 41224
rect 4771 41264 4829 41265
rect 4771 41224 4780 41264
rect 4820 41224 4829 41264
rect 6787 41264 6845 41265
rect 4771 41223 4829 41224
rect 5307 41254 5349 41263
rect 5307 41214 5308 41254
rect 5348 41214 5349 41254
rect 6787 41224 6796 41264
rect 6836 41224 6845 41264
rect 6787 41223 6845 41224
rect 8035 41264 8093 41265
rect 8035 41224 8044 41264
rect 8084 41224 8093 41264
rect 8035 41223 8093 41224
rect 8523 41264 8565 41273
rect 8523 41224 8524 41264
rect 8564 41224 8565 41264
rect 8523 41215 8565 41224
rect 8619 41264 8661 41273
rect 8619 41224 8620 41264
rect 8660 41224 8661 41264
rect 8619 41215 8661 41224
rect 9571 41264 9629 41265
rect 9571 41224 9580 41264
rect 9620 41224 9629 41264
rect 9571 41223 9629 41224
rect 10059 41259 10101 41268
rect 10059 41219 10060 41259
rect 10100 41219 10101 41259
rect 11971 41264 12029 41265
rect 11971 41224 11980 41264
rect 12020 41224 12029 41264
rect 11971 41223 12029 41224
rect 13219 41264 13277 41265
rect 13219 41224 13228 41264
rect 13268 41224 13277 41264
rect 13219 41223 13277 41224
rect 14379 41264 14421 41273
rect 14379 41224 14380 41264
rect 14420 41224 14421 41264
rect 5307 41205 5349 41214
rect 10059 41210 10101 41219
rect 14379 41215 14421 41224
rect 14475 41264 14517 41273
rect 14475 41224 14476 41264
rect 14516 41224 14517 41264
rect 14475 41215 14517 41224
rect 14955 41264 14997 41273
rect 14955 41224 14956 41264
rect 14996 41224 14997 41264
rect 14955 41215 14997 41224
rect 15427 41264 15485 41265
rect 15427 41224 15436 41264
rect 15476 41224 15485 41264
rect 15427 41223 15485 41224
rect 15963 41254 16005 41263
rect 15963 41214 15964 41254
rect 16004 41214 16005 41254
rect 15963 41205 16005 41214
rect 4203 41180 4245 41189
rect 4203 41140 4204 41180
rect 4244 41140 4245 41180
rect 4203 41131 4245 41140
rect 9003 41180 9045 41189
rect 9003 41140 9004 41180
rect 9044 41140 9045 41180
rect 9003 41131 9045 41140
rect 9099 41180 9141 41189
rect 9099 41140 9100 41180
rect 9140 41140 9141 41180
rect 9099 41131 9141 41140
rect 14859 41180 14901 41189
rect 14859 41140 14860 41180
rect 14900 41140 14901 41180
rect 14859 41131 14901 41140
rect 19267 41180 19325 41181
rect 19267 41140 19276 41180
rect 19316 41140 19325 41180
rect 19267 41139 19325 41140
rect 19651 41180 19709 41181
rect 19651 41140 19660 41180
rect 19700 41140 19709 41180
rect 19651 41139 19709 41140
rect 17259 41096 17301 41105
rect 17259 41056 17260 41096
rect 17300 41056 17301 41096
rect 17259 41047 17301 41056
rect 19467 41096 19509 41105
rect 19467 41056 19468 41096
rect 19508 41056 19509 41096
rect 19467 41047 19509 41056
rect 1152 40844 20352 40868
rect 1152 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 20352 40844
rect 1152 40780 20352 40804
rect 8235 40676 8277 40685
rect 8235 40636 8236 40676
rect 8276 40636 8277 40676
rect 8235 40627 8277 40636
rect 14091 40676 14133 40685
rect 14091 40636 14092 40676
rect 14132 40636 14133 40676
rect 14091 40627 14133 40636
rect 19563 40676 19605 40685
rect 19563 40636 19564 40676
rect 19604 40636 19605 40676
rect 19563 40627 19605 40636
rect 3339 40592 3381 40601
rect 3339 40552 3340 40592
rect 3380 40552 3381 40592
rect 3339 40543 3381 40552
rect 16395 40592 16437 40601
rect 16395 40552 16396 40592
rect 16436 40552 16437 40592
rect 16395 40543 16437 40552
rect 18027 40592 18069 40601
rect 18027 40552 18028 40592
rect 18068 40552 18069 40592
rect 18027 40543 18069 40552
rect 14955 40508 14997 40517
rect 14955 40468 14956 40508
rect 14996 40468 14997 40508
rect 14955 40459 14997 40468
rect 17827 40508 17885 40509
rect 17827 40468 17836 40508
rect 17876 40468 17885 40508
rect 17827 40467 17885 40468
rect 18979 40508 19037 40509
rect 18979 40468 18988 40508
rect 19028 40468 19037 40508
rect 18979 40467 19037 40468
rect 19363 40508 19421 40509
rect 19363 40468 19372 40508
rect 19412 40468 19421 40508
rect 19363 40467 19421 40468
rect 1891 40424 1949 40425
rect 1891 40384 1900 40424
rect 1940 40384 1949 40424
rect 1891 40383 1949 40384
rect 3139 40424 3197 40425
rect 3139 40384 3148 40424
rect 3188 40384 3197 40424
rect 3139 40383 3197 40384
rect 3523 40424 3581 40425
rect 3523 40384 3532 40424
rect 3572 40384 3581 40424
rect 3523 40383 3581 40384
rect 4771 40424 4829 40425
rect 4771 40384 4780 40424
rect 4820 40384 4829 40424
rect 4771 40383 4829 40384
rect 5155 40424 5213 40425
rect 5155 40384 5164 40424
rect 5204 40384 5213 40424
rect 5155 40383 5213 40384
rect 6403 40424 6461 40425
rect 6403 40384 6412 40424
rect 6452 40384 6461 40424
rect 6403 40383 6461 40384
rect 6787 40424 6845 40425
rect 6787 40384 6796 40424
rect 6836 40384 6845 40424
rect 6787 40383 6845 40384
rect 8035 40424 8093 40425
rect 8035 40384 8044 40424
rect 8084 40384 8093 40424
rect 8035 40383 8093 40384
rect 10723 40424 10781 40425
rect 10723 40384 10732 40424
rect 10772 40384 10781 40424
rect 10723 40383 10781 40384
rect 11971 40424 12029 40425
rect 11971 40384 11980 40424
rect 12020 40384 12029 40424
rect 11971 40383 12029 40384
rect 12643 40424 12701 40425
rect 12643 40384 12652 40424
rect 12692 40384 12701 40424
rect 12643 40383 12701 40384
rect 13891 40424 13949 40425
rect 13891 40384 13900 40424
rect 13940 40384 13949 40424
rect 13891 40383 13949 40384
rect 14379 40424 14421 40433
rect 14379 40384 14380 40424
rect 14420 40384 14421 40424
rect 14379 40375 14421 40384
rect 14475 40424 14517 40433
rect 14475 40384 14476 40424
rect 14516 40384 14517 40424
rect 14475 40375 14517 40384
rect 14859 40424 14901 40433
rect 15915 40429 15957 40438
rect 14859 40384 14860 40424
rect 14900 40384 14901 40424
rect 14859 40375 14901 40384
rect 15427 40424 15485 40425
rect 15427 40384 15436 40424
rect 15476 40384 15485 40424
rect 15427 40383 15485 40384
rect 15915 40389 15916 40429
rect 15956 40389 15957 40429
rect 15915 40380 15957 40389
rect 4971 40340 5013 40349
rect 4971 40300 4972 40340
rect 5012 40300 5013 40340
rect 4971 40291 5013 40300
rect 6603 40340 6645 40349
rect 6603 40300 6604 40340
rect 6644 40300 6645 40340
rect 6603 40291 6645 40300
rect 8419 40256 8477 40257
rect 8419 40216 8428 40256
rect 8468 40216 8477 40256
rect 8419 40215 8477 40216
rect 9099 40256 9141 40265
rect 9099 40216 9100 40256
rect 9140 40216 9141 40256
rect 9099 40207 9141 40216
rect 12171 40256 12213 40265
rect 12171 40216 12172 40256
rect 12212 40216 12213 40256
rect 12171 40207 12213 40216
rect 16107 40256 16149 40265
rect 16107 40216 16108 40256
rect 16148 40216 16149 40256
rect 16107 40207 16149 40216
rect 17251 40256 17309 40257
rect 17251 40216 17260 40256
rect 17300 40216 17309 40256
rect 17251 40215 17309 40216
rect 19179 40256 19221 40265
rect 19179 40216 19180 40256
rect 19220 40216 19221 40256
rect 19179 40207 19221 40216
rect 1152 40088 20452 40112
rect 1152 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20452 40088
rect 1152 40024 20452 40048
rect 2667 39920 2709 39929
rect 2667 39880 2668 39920
rect 2708 39880 2709 39920
rect 2667 39871 2709 39880
rect 9099 39920 9141 39929
rect 9099 39880 9100 39920
rect 9140 39880 9141 39920
rect 9099 39871 9141 39880
rect 14667 39920 14709 39929
rect 14667 39880 14668 39920
rect 14708 39880 14709 39920
rect 14667 39871 14709 39880
rect 16395 39920 16437 39929
rect 16395 39880 16396 39920
rect 16436 39880 16437 39920
rect 16395 39871 16437 39880
rect 17251 39920 17309 39921
rect 17251 39880 17260 39920
rect 17300 39880 17309 39920
rect 17251 39879 17309 39880
rect 18979 39920 19037 39921
rect 18979 39880 18988 39920
rect 19028 39880 19037 39920
rect 18979 39879 19037 39880
rect 5547 39836 5589 39845
rect 5547 39796 5548 39836
rect 5588 39796 5589 39836
rect 5547 39787 5589 39796
rect 8139 39836 8181 39845
rect 8139 39796 8140 39836
rect 8180 39796 8181 39836
rect 8139 39787 8181 39796
rect 11115 39836 11157 39845
rect 11115 39796 11116 39836
rect 11156 39796 11157 39836
rect 11115 39787 11157 39796
rect 14187 39836 14229 39845
rect 14187 39796 14188 39836
rect 14228 39796 14229 39836
rect 14187 39787 14229 39796
rect 1219 39752 1277 39753
rect 1219 39712 1228 39752
rect 1268 39712 1277 39752
rect 1219 39711 1277 39712
rect 2467 39752 2525 39753
rect 2467 39712 2476 39752
rect 2516 39712 2525 39752
rect 2467 39711 2525 39712
rect 3819 39752 3861 39761
rect 3819 39712 3820 39752
rect 3860 39712 3861 39752
rect 3819 39703 3861 39712
rect 3915 39752 3957 39761
rect 3915 39712 3916 39752
rect 3956 39712 3957 39752
rect 3915 39703 3957 39712
rect 4395 39752 4437 39761
rect 4395 39712 4396 39752
rect 4436 39712 4437 39752
rect 4395 39703 4437 39712
rect 4867 39752 4925 39753
rect 4867 39712 4876 39752
rect 4916 39712 4925 39752
rect 4867 39711 4925 39712
rect 5355 39747 5397 39756
rect 5355 39707 5356 39747
rect 5396 39707 5397 39747
rect 5355 39698 5397 39707
rect 6411 39752 6453 39761
rect 6411 39712 6412 39752
rect 6452 39712 6453 39752
rect 6411 39703 6453 39712
rect 6507 39752 6549 39761
rect 6507 39712 6508 39752
rect 6548 39712 6549 39752
rect 6507 39703 6549 39712
rect 6891 39752 6933 39761
rect 6891 39712 6892 39752
rect 6932 39712 6933 39752
rect 6891 39703 6933 39712
rect 7459 39752 7517 39753
rect 7459 39712 7468 39752
rect 7508 39712 7517 39752
rect 9387 39752 9429 39761
rect 7459 39711 7517 39712
rect 7947 39738 7989 39747
rect 7947 39698 7948 39738
rect 7988 39698 7989 39738
rect 9387 39712 9388 39752
rect 9428 39712 9429 39752
rect 9387 39703 9429 39712
rect 9483 39752 9525 39761
rect 9483 39712 9484 39752
rect 9524 39712 9525 39752
rect 9483 39703 9525 39712
rect 9963 39752 10005 39761
rect 9963 39712 9964 39752
rect 10004 39712 10005 39752
rect 9963 39703 10005 39712
rect 10435 39752 10493 39753
rect 10435 39712 10444 39752
rect 10484 39712 10493 39752
rect 12459 39752 12501 39761
rect 10435 39711 10493 39712
rect 10923 39738 10965 39747
rect 7947 39689 7989 39698
rect 10923 39698 10924 39738
rect 10964 39698 10965 39738
rect 12459 39712 12460 39752
rect 12500 39712 12501 39752
rect 12459 39703 12501 39712
rect 12555 39752 12597 39761
rect 12555 39712 12556 39752
rect 12596 39712 12597 39752
rect 12555 39703 12597 39712
rect 13035 39752 13077 39761
rect 13035 39712 13036 39752
rect 13076 39712 13077 39752
rect 13035 39703 13077 39712
rect 13507 39752 13565 39753
rect 13507 39712 13516 39752
rect 13556 39712 13565 39752
rect 14851 39752 14909 39753
rect 13507 39711 13565 39712
rect 13995 39738 14037 39747
rect 10923 39689 10965 39698
rect 13995 39698 13996 39738
rect 14036 39698 14037 39738
rect 14851 39712 14860 39752
rect 14900 39712 14909 39752
rect 14851 39711 14909 39712
rect 16099 39752 16157 39753
rect 16099 39712 16108 39752
rect 16148 39712 16157 39752
rect 16099 39711 16157 39712
rect 13995 39689 14037 39698
rect 4299 39668 4341 39677
rect 4299 39628 4300 39668
rect 4340 39628 4341 39668
rect 4299 39619 4341 39628
rect 6987 39668 7029 39677
rect 6987 39628 6988 39668
rect 7028 39628 7029 39668
rect 6987 39619 7029 39628
rect 9867 39668 9909 39677
rect 9867 39628 9868 39668
rect 9908 39628 9909 39668
rect 9867 39619 9909 39628
rect 12939 39668 12981 39677
rect 12939 39628 12940 39668
rect 12980 39628 12981 39668
rect 12939 39619 12981 39628
rect 19267 39668 19325 39669
rect 19267 39628 19276 39668
rect 19316 39628 19325 39668
rect 19267 39627 19325 39628
rect 19651 39668 19709 39669
rect 19651 39628 19660 39668
rect 19700 39628 19709 39668
rect 19651 39627 19709 39628
rect 9003 39584 9045 39593
rect 9003 39544 9004 39584
rect 9044 39544 9045 39584
rect 9003 39535 9045 39544
rect 16299 39584 16341 39593
rect 16299 39544 16300 39584
rect 16340 39544 16341 39584
rect 16299 39535 16341 39544
rect 17355 39584 17397 39593
rect 17355 39544 17356 39584
rect 17396 39544 17397 39584
rect 17355 39535 17397 39544
rect 19851 39584 19893 39593
rect 19851 39544 19852 39584
rect 19892 39544 19893 39584
rect 19851 39535 19893 39544
rect 19467 39500 19509 39509
rect 19467 39460 19468 39500
rect 19508 39460 19509 39500
rect 19467 39451 19509 39460
rect 1152 39332 20352 39356
rect 1152 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 20352 39332
rect 1152 39268 20352 39292
rect 7179 39080 7221 39089
rect 7179 39040 7180 39080
rect 7220 39040 7221 39080
rect 7179 39031 7221 39040
rect 8811 39080 8853 39089
rect 8811 39040 8812 39080
rect 8852 39040 8853 39080
rect 8811 39031 8853 39040
rect 12459 39080 12501 39089
rect 12459 39040 12460 39080
rect 12500 39040 12501 39080
rect 12459 39031 12501 39040
rect 16299 39080 16341 39089
rect 16299 39040 16300 39080
rect 16340 39040 16341 39080
rect 16299 39031 16341 39040
rect 17259 39080 17301 39089
rect 17259 39040 17260 39080
rect 17300 39040 17301 39080
rect 17259 39031 17301 39040
rect 19851 39080 19893 39089
rect 19851 39040 19852 39080
rect 19892 39040 19893 39080
rect 19851 39031 19893 39040
rect 3051 38996 3093 39005
rect 3051 38956 3052 38996
rect 3092 38956 3093 38996
rect 3051 38947 3093 38956
rect 14955 38996 14997 39005
rect 14955 38956 14956 38996
rect 14996 38956 14997 38996
rect 14955 38947 14997 38956
rect 19267 38996 19325 38997
rect 19267 38956 19276 38996
rect 19316 38956 19325 38996
rect 19267 38955 19325 38956
rect 19651 38996 19709 38997
rect 19651 38956 19660 38996
rect 19700 38956 19709 38996
rect 19651 38955 19709 38956
rect 20035 38996 20093 38997
rect 20035 38956 20044 38996
rect 20084 38956 20093 38996
rect 20035 38955 20093 38956
rect 2475 38912 2517 38921
rect 2475 38872 2476 38912
rect 2516 38872 2517 38912
rect 2475 38863 2517 38872
rect 2571 38912 2613 38921
rect 2571 38872 2572 38912
rect 2612 38872 2613 38912
rect 2571 38863 2613 38872
rect 2955 38912 2997 38921
rect 4011 38917 4053 38926
rect 15963 38921 16005 38930
rect 2955 38872 2956 38912
rect 2996 38872 2997 38912
rect 2955 38863 2997 38872
rect 3523 38912 3581 38913
rect 3523 38872 3532 38912
rect 3572 38872 3581 38912
rect 3523 38871 3581 38872
rect 4011 38877 4012 38917
rect 4052 38877 4053 38917
rect 4011 38868 4053 38877
rect 5731 38912 5789 38913
rect 5731 38872 5740 38912
rect 5780 38872 5789 38912
rect 5731 38871 5789 38872
rect 6979 38912 7037 38913
rect 6979 38872 6988 38912
rect 7028 38872 7037 38912
rect 6979 38871 7037 38872
rect 7363 38912 7421 38913
rect 7363 38872 7372 38912
rect 7412 38872 7421 38912
rect 7363 38871 7421 38872
rect 8611 38912 8669 38913
rect 8611 38872 8620 38912
rect 8660 38872 8669 38912
rect 8611 38871 8669 38872
rect 8995 38912 9053 38913
rect 8995 38872 9004 38912
rect 9044 38872 9053 38912
rect 8995 38871 9053 38872
rect 10243 38912 10301 38913
rect 10243 38872 10252 38912
rect 10292 38872 10301 38912
rect 10243 38871 10301 38872
rect 11011 38912 11069 38913
rect 11011 38872 11020 38912
rect 11060 38872 11069 38912
rect 11011 38871 11069 38872
rect 12259 38912 12317 38913
rect 12259 38872 12268 38912
rect 12308 38872 12317 38912
rect 12259 38871 12317 38872
rect 12643 38912 12701 38913
rect 12643 38872 12652 38912
rect 12692 38872 12701 38912
rect 12643 38871 12701 38872
rect 13891 38912 13949 38913
rect 13891 38872 13900 38912
rect 13940 38872 13949 38912
rect 13891 38871 13949 38872
rect 14379 38912 14421 38921
rect 14379 38872 14380 38912
rect 14420 38872 14421 38912
rect 14379 38863 14421 38872
rect 14475 38912 14517 38921
rect 14475 38872 14476 38912
rect 14516 38872 14517 38912
rect 14475 38863 14517 38872
rect 14859 38912 14901 38921
rect 14859 38872 14860 38912
rect 14900 38872 14901 38912
rect 14859 38863 14901 38872
rect 15427 38912 15485 38913
rect 15427 38872 15436 38912
rect 15476 38872 15485 38912
rect 15963 38881 15964 38921
rect 16004 38881 16005 38921
rect 15963 38872 16005 38881
rect 17443 38912 17501 38913
rect 17443 38872 17452 38912
rect 17492 38872 17501 38912
rect 15427 38871 15485 38872
rect 17443 38871 17501 38872
rect 18691 38912 18749 38913
rect 18691 38872 18700 38912
rect 18740 38872 18749 38912
rect 18691 38871 18749 38872
rect 4203 38828 4245 38837
rect 4203 38788 4204 38828
rect 4244 38788 4245 38828
rect 4203 38779 4245 38788
rect 14091 38828 14133 38837
rect 14091 38788 14092 38828
rect 14132 38788 14133 38828
rect 14091 38779 14133 38788
rect 16107 38828 16149 38837
rect 16107 38788 16108 38828
rect 16148 38788 16149 38828
rect 16107 38779 16149 38788
rect 10443 38744 10485 38753
rect 10443 38704 10444 38744
rect 10484 38704 10485 38744
rect 10443 38695 10485 38704
rect 18979 38744 19037 38745
rect 18979 38704 18988 38744
rect 19028 38704 19037 38744
rect 18979 38703 19037 38704
rect 19467 38744 19509 38753
rect 19467 38704 19468 38744
rect 19508 38704 19509 38744
rect 19467 38695 19509 38704
rect 20235 38744 20277 38753
rect 20235 38704 20236 38744
rect 20276 38704 20277 38744
rect 20235 38695 20277 38704
rect 1152 38576 20452 38600
rect 1152 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20452 38576
rect 1152 38512 20452 38536
rect 2667 38408 2709 38417
rect 2667 38368 2668 38408
rect 2708 38368 2709 38408
rect 2667 38359 2709 38368
rect 4683 38408 4725 38417
rect 4683 38368 4684 38408
rect 4724 38368 4725 38408
rect 4683 38359 4725 38368
rect 8995 38408 9053 38409
rect 8995 38368 9004 38408
rect 9044 38368 9053 38408
rect 8995 38367 9053 38368
rect 16107 38408 16149 38417
rect 16107 38368 16108 38408
rect 16148 38368 16149 38408
rect 16107 38359 16149 38368
rect 16395 38408 16437 38417
rect 16395 38368 16396 38408
rect 16436 38368 16437 38408
rect 16395 38359 16437 38368
rect 17251 38408 17309 38409
rect 17251 38368 17260 38408
rect 17300 38368 17309 38408
rect 17251 38367 17309 38368
rect 18979 38408 19037 38409
rect 18979 38368 18988 38408
rect 19028 38368 19037 38408
rect 18979 38367 19037 38368
rect 19467 38408 19509 38417
rect 19467 38368 19468 38408
rect 19508 38368 19509 38408
rect 19467 38359 19509 38368
rect 7947 38324 7989 38333
rect 7947 38284 7948 38324
rect 7988 38284 7989 38324
rect 7947 38275 7989 38284
rect 11883 38324 11925 38333
rect 11883 38284 11884 38324
rect 11924 38284 11925 38324
rect 11883 38275 11925 38284
rect 13995 38324 14037 38333
rect 13995 38284 13996 38324
rect 14036 38284 14037 38324
rect 13995 38275 14037 38284
rect 1219 38240 1277 38241
rect 1219 38200 1228 38240
rect 1268 38200 1277 38240
rect 1219 38199 1277 38200
rect 2467 38240 2525 38241
rect 2467 38200 2476 38240
rect 2516 38200 2525 38240
rect 2467 38199 2525 38200
rect 2955 38240 2997 38249
rect 2955 38200 2956 38240
rect 2996 38200 2997 38240
rect 2955 38191 2997 38200
rect 3051 38240 3093 38249
rect 3051 38200 3052 38240
rect 3092 38200 3093 38240
rect 3051 38191 3093 38200
rect 3435 38240 3477 38249
rect 3435 38200 3436 38240
rect 3476 38200 3477 38240
rect 3435 38191 3477 38200
rect 3531 38240 3573 38249
rect 3531 38200 3532 38240
rect 3572 38200 3573 38240
rect 3531 38191 3573 38200
rect 4003 38240 4061 38241
rect 4003 38200 4012 38240
rect 4052 38200 4061 38240
rect 6219 38240 6261 38249
rect 4003 38199 4061 38200
rect 4491 38226 4533 38235
rect 4491 38186 4492 38226
rect 4532 38186 4533 38226
rect 6219 38200 6220 38240
rect 6260 38200 6261 38240
rect 6219 38191 6261 38200
rect 6315 38240 6357 38249
rect 6315 38200 6316 38240
rect 6356 38200 6357 38240
rect 6315 38191 6357 38200
rect 6699 38240 6741 38249
rect 6699 38200 6700 38240
rect 6740 38200 6741 38240
rect 6699 38191 6741 38200
rect 6795 38240 6837 38249
rect 6795 38200 6796 38240
rect 6836 38200 6837 38240
rect 6795 38191 6837 38200
rect 7267 38240 7325 38241
rect 7267 38200 7276 38240
rect 7316 38200 7325 38240
rect 8139 38240 8181 38249
rect 7267 38199 7325 38200
rect 7755 38226 7797 38235
rect 4491 38177 4533 38186
rect 7755 38186 7756 38226
rect 7796 38186 7797 38226
rect 8139 38200 8140 38240
rect 8180 38200 8181 38240
rect 8139 38191 8181 38200
rect 8331 38240 8373 38249
rect 8331 38200 8332 38240
rect 8372 38200 8373 38240
rect 8331 38191 8373 38200
rect 9675 38240 9717 38249
rect 9675 38200 9676 38240
rect 9716 38200 9717 38240
rect 9675 38191 9717 38200
rect 9859 38240 9917 38241
rect 9859 38200 9868 38240
rect 9908 38200 9917 38240
rect 9859 38199 9917 38200
rect 10155 38240 10197 38249
rect 10155 38200 10156 38240
rect 10196 38200 10197 38240
rect 10155 38191 10197 38200
rect 10251 38240 10293 38249
rect 10251 38200 10252 38240
rect 10292 38200 10293 38240
rect 10251 38191 10293 38200
rect 11203 38240 11261 38241
rect 11203 38200 11212 38240
rect 11252 38200 11261 38240
rect 11203 38199 11261 38200
rect 11691 38235 11733 38244
rect 11691 38195 11692 38235
rect 11732 38195 11733 38235
rect 11691 38186 11733 38195
rect 12267 38240 12309 38249
rect 12267 38200 12268 38240
rect 12308 38200 12309 38240
rect 12267 38191 12309 38200
rect 12363 38240 12405 38249
rect 12363 38200 12364 38240
rect 12404 38200 12405 38240
rect 12363 38191 12405 38200
rect 13315 38240 13373 38241
rect 13315 38200 13324 38240
rect 13364 38200 13373 38240
rect 14659 38240 14717 38241
rect 13315 38199 13373 38200
rect 13803 38226 13845 38235
rect 13803 38186 13804 38226
rect 13844 38186 13845 38226
rect 14659 38200 14668 38240
rect 14708 38200 14717 38240
rect 14659 38199 14717 38200
rect 15907 38240 15965 38241
rect 15907 38200 15916 38240
rect 15956 38200 15965 38240
rect 15907 38199 15965 38200
rect 7755 38177 7797 38186
rect 13803 38177 13845 38186
rect 10635 38156 10677 38165
rect 10635 38116 10636 38156
rect 10676 38116 10677 38156
rect 10635 38107 10677 38116
rect 10731 38156 10773 38165
rect 10731 38116 10732 38156
rect 10772 38116 10773 38156
rect 10731 38107 10773 38116
rect 12747 38156 12789 38165
rect 12747 38116 12748 38156
rect 12788 38116 12789 38156
rect 12747 38107 12789 38116
rect 12843 38156 12885 38165
rect 12843 38116 12844 38156
rect 12884 38116 12885 38156
rect 12843 38107 12885 38116
rect 18595 38156 18653 38157
rect 18595 38116 18604 38156
rect 18644 38116 18653 38156
rect 18595 38115 18653 38116
rect 19267 38156 19325 38157
rect 19267 38116 19276 38156
rect 19316 38116 19325 38156
rect 19267 38115 19325 38116
rect 19651 38156 19709 38157
rect 19651 38116 19660 38156
rect 19700 38116 19709 38156
rect 19651 38115 19709 38116
rect 20035 38156 20093 38157
rect 20035 38116 20044 38156
rect 20084 38116 20093 38156
rect 20035 38115 20093 38116
rect 19083 38072 19125 38081
rect 19083 38032 19084 38072
rect 19124 38032 19125 38072
rect 19083 38023 19125 38032
rect 20235 38072 20277 38081
rect 20235 38032 20236 38072
rect 20276 38032 20277 38072
rect 20235 38023 20277 38032
rect 8139 37988 8181 37997
rect 8139 37948 8140 37988
rect 8180 37948 8181 37988
rect 8139 37939 8181 37948
rect 9771 37988 9813 37997
rect 9771 37948 9772 37988
rect 9812 37948 9813 37988
rect 9771 37939 9813 37948
rect 18795 37988 18837 37997
rect 18795 37948 18796 37988
rect 18836 37948 18837 37988
rect 18795 37939 18837 37948
rect 19851 37988 19893 37997
rect 19851 37948 19852 37988
rect 19892 37948 19893 37988
rect 19851 37939 19893 37948
rect 1152 37820 20352 37844
rect 1152 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 20352 37820
rect 1152 37756 20352 37780
rect 3915 37652 3957 37661
rect 3915 37612 3916 37652
rect 3956 37612 3957 37652
rect 3915 37603 3957 37612
rect 5547 37652 5589 37661
rect 5547 37612 5548 37652
rect 5588 37612 5589 37652
rect 5547 37603 5589 37612
rect 7179 37652 7221 37661
rect 7179 37612 7180 37652
rect 7220 37612 7221 37652
rect 7179 37603 7221 37612
rect 8811 37652 8853 37661
rect 8811 37612 8812 37652
rect 8852 37612 8853 37652
rect 8811 37603 8853 37612
rect 12075 37652 12117 37661
rect 12075 37612 12076 37652
rect 12116 37612 12117 37652
rect 12075 37603 12117 37612
rect 13707 37652 13749 37661
rect 13707 37612 13708 37652
rect 13748 37612 13749 37652
rect 13707 37603 13749 37612
rect 10155 37568 10197 37577
rect 10155 37528 10156 37568
rect 10196 37528 10197 37568
rect 10155 37519 10197 37528
rect 19083 37568 19125 37577
rect 19083 37528 19084 37568
rect 19124 37528 19125 37568
rect 19083 37519 19125 37528
rect 15819 37484 15861 37493
rect 15819 37444 15820 37484
rect 15860 37444 15861 37484
rect 15819 37435 15861 37444
rect 15915 37484 15957 37493
rect 15915 37444 15916 37484
rect 15956 37444 15957 37484
rect 15915 37435 15957 37444
rect 19267 37484 19325 37485
rect 19267 37444 19276 37484
rect 19316 37444 19325 37484
rect 19267 37443 19325 37444
rect 19651 37484 19709 37485
rect 19651 37444 19660 37484
rect 19700 37444 19709 37484
rect 19651 37443 19709 37444
rect 20035 37484 20093 37485
rect 20035 37444 20044 37484
rect 20084 37444 20093 37484
rect 20035 37443 20093 37444
rect 16923 37409 16965 37418
rect 2467 37400 2525 37401
rect 2467 37360 2476 37400
rect 2516 37360 2525 37400
rect 2467 37359 2525 37360
rect 3715 37400 3773 37401
rect 3715 37360 3724 37400
rect 3764 37360 3773 37400
rect 3715 37359 3773 37360
rect 4099 37400 4157 37401
rect 4099 37360 4108 37400
rect 4148 37360 4157 37400
rect 4099 37359 4157 37360
rect 5347 37400 5405 37401
rect 5347 37360 5356 37400
rect 5396 37360 5405 37400
rect 5347 37359 5405 37360
rect 5731 37400 5789 37401
rect 5731 37360 5740 37400
rect 5780 37360 5789 37400
rect 5731 37359 5789 37360
rect 6979 37400 7037 37401
rect 6979 37360 6988 37400
rect 7028 37360 7037 37400
rect 6979 37359 7037 37360
rect 7363 37400 7421 37401
rect 7363 37360 7372 37400
rect 7412 37360 7421 37400
rect 7363 37359 7421 37360
rect 8611 37400 8669 37401
rect 8611 37360 8620 37400
rect 8660 37360 8669 37400
rect 8611 37359 8669 37360
rect 9379 37400 9437 37401
rect 9379 37360 9388 37400
rect 9428 37360 9437 37400
rect 9379 37359 9437 37360
rect 9579 37400 9621 37409
rect 9579 37360 9580 37400
rect 9620 37360 9621 37400
rect 9579 37351 9621 37360
rect 9667 37400 9725 37401
rect 9667 37360 9676 37400
rect 9716 37360 9725 37400
rect 9667 37359 9725 37360
rect 10627 37400 10685 37401
rect 10627 37360 10636 37400
rect 10676 37360 10685 37400
rect 10627 37359 10685 37360
rect 11875 37400 11933 37401
rect 11875 37360 11884 37400
rect 11924 37360 11933 37400
rect 11875 37359 11933 37360
rect 12259 37400 12317 37401
rect 12259 37360 12268 37400
rect 12308 37360 12317 37400
rect 12259 37359 12317 37360
rect 13507 37400 13565 37401
rect 13507 37360 13516 37400
rect 13556 37360 13565 37400
rect 13507 37359 13565 37360
rect 15339 37400 15381 37409
rect 15339 37360 15340 37400
rect 15380 37360 15381 37400
rect 15339 37351 15381 37360
rect 15435 37400 15477 37409
rect 15435 37360 15436 37400
rect 15476 37360 15477 37400
rect 15435 37351 15477 37360
rect 16387 37400 16445 37401
rect 16387 37360 16396 37400
rect 16436 37360 16445 37400
rect 16923 37369 16924 37409
rect 16964 37369 16965 37409
rect 16923 37360 16965 37369
rect 16387 37359 16445 37360
rect 17067 37316 17109 37325
rect 17067 37276 17068 37316
rect 17108 37276 17109 37316
rect 17067 37267 17109 37276
rect 8995 37232 9053 37233
rect 8995 37192 9004 37232
rect 9044 37192 9053 37232
rect 8995 37191 9053 37192
rect 9387 37232 9429 37241
rect 9387 37192 9388 37232
rect 9428 37192 9429 37232
rect 9387 37183 9429 37192
rect 10051 37232 10109 37233
rect 10051 37192 10060 37232
rect 10100 37192 10109 37232
rect 10051 37191 10109 37192
rect 17251 37232 17309 37233
rect 17251 37192 17260 37232
rect 17300 37192 17309 37232
rect 17251 37191 17309 37192
rect 19467 37232 19509 37241
rect 19467 37192 19468 37232
rect 19508 37192 19509 37232
rect 19467 37183 19509 37192
rect 19851 37232 19893 37241
rect 19851 37192 19852 37232
rect 19892 37192 19893 37232
rect 19851 37183 19893 37192
rect 20235 37232 20277 37241
rect 20235 37192 20236 37232
rect 20276 37192 20277 37232
rect 20235 37183 20277 37192
rect 1152 37064 20452 37088
rect 1152 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20452 37064
rect 1152 37000 20452 37024
rect 2667 36896 2709 36905
rect 2667 36856 2668 36896
rect 2708 36856 2709 36896
rect 2667 36847 2709 36856
rect 9571 36896 9629 36897
rect 9571 36856 9580 36896
rect 9620 36856 9629 36896
rect 9571 36855 9629 36856
rect 19083 36896 19125 36905
rect 19083 36856 19084 36896
rect 19124 36856 19125 36896
rect 19083 36847 19125 36856
rect 12939 36812 12981 36821
rect 12939 36772 12940 36812
rect 12980 36772 12981 36812
rect 12939 36763 12981 36772
rect 14955 36812 14997 36821
rect 14955 36772 14956 36812
rect 14996 36772 14997 36812
rect 14955 36763 14997 36772
rect 16971 36812 17013 36821
rect 16971 36772 16972 36812
rect 17012 36772 17013 36812
rect 16971 36763 17013 36772
rect 1219 36728 1277 36729
rect 1219 36688 1228 36728
rect 1268 36688 1277 36728
rect 1219 36687 1277 36688
rect 2467 36728 2525 36729
rect 2467 36688 2476 36728
rect 2516 36688 2525 36728
rect 2467 36687 2525 36688
rect 3331 36728 3389 36729
rect 3331 36688 3340 36728
rect 3380 36688 3389 36728
rect 3331 36687 3389 36688
rect 4579 36728 4637 36729
rect 4579 36688 4588 36728
rect 4628 36688 4637 36728
rect 4579 36687 4637 36688
rect 5539 36728 5597 36729
rect 5539 36688 5548 36728
rect 5588 36688 5597 36728
rect 5539 36687 5597 36688
rect 6787 36728 6845 36729
rect 6787 36688 6796 36728
rect 6836 36688 6845 36728
rect 6787 36687 6845 36688
rect 7363 36728 7421 36729
rect 7363 36688 7372 36728
rect 7412 36688 7421 36728
rect 7363 36687 7421 36688
rect 8611 36728 8669 36729
rect 8611 36688 8620 36728
rect 8660 36688 8669 36728
rect 8611 36687 8669 36688
rect 9771 36728 9813 36737
rect 9771 36688 9772 36728
rect 9812 36688 9813 36728
rect 9771 36679 9813 36688
rect 9867 36728 9909 36737
rect 9867 36688 9868 36728
rect 9908 36688 9909 36728
rect 9867 36679 9909 36688
rect 10627 36728 10685 36729
rect 10627 36688 10636 36728
rect 10676 36688 10685 36728
rect 10627 36687 10685 36688
rect 10923 36728 10965 36737
rect 10923 36688 10924 36728
rect 10964 36688 10965 36728
rect 10923 36679 10965 36688
rect 11019 36728 11061 36737
rect 11019 36688 11020 36728
rect 11060 36688 11061 36728
rect 11019 36679 11061 36688
rect 11491 36728 11549 36729
rect 11491 36688 11500 36728
rect 11540 36688 11549 36728
rect 11491 36687 11549 36688
rect 12739 36728 12797 36729
rect 12739 36688 12748 36728
rect 12788 36688 12797 36728
rect 12739 36687 12797 36688
rect 13227 36728 13269 36737
rect 13227 36688 13228 36728
rect 13268 36688 13269 36728
rect 13227 36679 13269 36688
rect 13323 36728 13365 36737
rect 13323 36688 13324 36728
rect 13364 36688 13365 36728
rect 13323 36679 13365 36688
rect 14275 36728 14333 36729
rect 14275 36688 14284 36728
rect 14324 36688 14333 36728
rect 15243 36728 15285 36737
rect 14275 36687 14333 36688
rect 14763 36714 14805 36723
rect 14763 36674 14764 36714
rect 14804 36674 14805 36714
rect 15243 36688 15244 36728
rect 15284 36688 15285 36728
rect 15243 36679 15285 36688
rect 15339 36728 15381 36737
rect 15339 36688 15340 36728
rect 15380 36688 15381 36728
rect 15339 36679 15381 36688
rect 15723 36728 15765 36737
rect 15723 36688 15724 36728
rect 15764 36688 15765 36728
rect 15723 36679 15765 36688
rect 15819 36728 15861 36737
rect 15819 36688 15820 36728
rect 15860 36688 15861 36728
rect 15819 36679 15861 36688
rect 16291 36728 16349 36729
rect 16291 36688 16300 36728
rect 16340 36688 16349 36728
rect 16291 36687 16349 36688
rect 16779 36714 16821 36723
rect 14763 36665 14805 36674
rect 16779 36674 16780 36714
rect 16820 36674 16821 36714
rect 16779 36665 16821 36674
rect 13707 36644 13749 36653
rect 13707 36604 13708 36644
rect 13748 36604 13749 36644
rect 13707 36595 13749 36604
rect 13803 36644 13845 36653
rect 13803 36604 13804 36644
rect 13844 36604 13845 36644
rect 13803 36595 13845 36604
rect 6987 36560 7029 36569
rect 6987 36520 6988 36560
rect 7028 36520 7029 36560
rect 6987 36511 7029 36520
rect 8811 36560 8853 36569
rect 8811 36520 8812 36560
rect 8852 36520 8853 36560
rect 8811 36511 8853 36520
rect 9003 36560 9045 36569
rect 9003 36520 9004 36560
rect 9044 36520 9045 36560
rect 9003 36511 9045 36520
rect 10059 36560 10101 36569
rect 10059 36520 10060 36560
rect 10100 36520 10101 36560
rect 10059 36511 10101 36520
rect 17259 36560 17301 36569
rect 17259 36520 17260 36560
rect 17300 36520 17301 36560
rect 17259 36511 17301 36520
rect 4779 36476 4821 36485
rect 4779 36436 4780 36476
rect 4820 36436 4821 36476
rect 4779 36427 4821 36436
rect 11299 36476 11357 36477
rect 11299 36436 11308 36476
rect 11348 36436 11357 36476
rect 11299 36435 11357 36436
rect 1152 36308 20352 36332
rect 1152 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 20352 36308
rect 1152 36244 20352 36268
rect 2667 36140 2709 36149
rect 2667 36100 2668 36140
rect 2708 36100 2709 36140
rect 2667 36091 2709 36100
rect 7179 36140 7221 36149
rect 7179 36100 7180 36140
rect 7220 36100 7221 36140
rect 7179 36091 7221 36100
rect 14283 36140 14325 36149
rect 14283 36100 14284 36140
rect 14324 36100 14325 36140
rect 14283 36091 14325 36100
rect 15147 36140 15189 36149
rect 15147 36100 15148 36140
rect 15188 36100 15189 36140
rect 15147 36091 15189 36100
rect 19755 36140 19797 36149
rect 19755 36100 19756 36140
rect 19796 36100 19797 36140
rect 19755 36091 19797 36100
rect 20139 36140 20181 36149
rect 20139 36100 20140 36140
rect 20180 36100 20181 36140
rect 20139 36091 20181 36100
rect 8811 36056 8853 36065
rect 8811 36016 8812 36056
rect 8852 36016 8853 36056
rect 8811 36007 8853 36016
rect 10051 36056 10109 36057
rect 10051 36016 10060 36056
rect 10100 36016 10109 36056
rect 10051 36015 10109 36016
rect 18123 35972 18165 35981
rect 4539 35930 4581 35939
rect 1219 35888 1277 35889
rect 1219 35848 1228 35888
rect 1268 35848 1277 35888
rect 1219 35847 1277 35848
rect 2467 35888 2525 35889
rect 2467 35848 2476 35888
rect 2516 35848 2525 35888
rect 2467 35847 2525 35848
rect 2955 35888 2997 35897
rect 2955 35848 2956 35888
rect 2996 35848 2997 35888
rect 2955 35839 2997 35848
rect 3051 35888 3093 35897
rect 3051 35848 3052 35888
rect 3092 35848 3093 35888
rect 3051 35839 3093 35848
rect 3435 35888 3477 35897
rect 3435 35848 3436 35888
rect 3476 35848 3477 35888
rect 3435 35839 3477 35848
rect 3531 35888 3573 35897
rect 4539 35890 4540 35930
rect 4580 35890 4581 35930
rect 18123 35932 18124 35972
rect 18164 35932 18165 35972
rect 18123 35923 18165 35932
rect 19555 35972 19613 35973
rect 19555 35932 19564 35972
rect 19604 35932 19613 35972
rect 19555 35931 19613 35932
rect 19939 35972 19997 35973
rect 19939 35932 19948 35972
rect 19988 35932 19997 35972
rect 19939 35931 19997 35932
rect 3531 35848 3532 35888
rect 3572 35848 3573 35888
rect 3531 35839 3573 35848
rect 4003 35888 4061 35889
rect 4003 35848 4012 35888
rect 4052 35848 4061 35888
rect 4539 35881 4581 35890
rect 5251 35888 5309 35889
rect 4003 35847 4061 35848
rect 5251 35848 5260 35888
rect 5300 35848 5309 35888
rect 5251 35847 5309 35848
rect 6499 35888 6557 35889
rect 6499 35848 6508 35888
rect 6548 35848 6557 35888
rect 6499 35847 6557 35848
rect 6883 35888 6941 35889
rect 6883 35848 6892 35888
rect 6932 35848 6941 35888
rect 6883 35847 6941 35848
rect 6987 35888 7029 35897
rect 6987 35848 6988 35888
rect 7028 35848 7029 35888
rect 6987 35839 7029 35848
rect 7179 35888 7221 35897
rect 7179 35848 7180 35888
rect 7220 35848 7221 35888
rect 7179 35839 7221 35848
rect 7363 35888 7421 35889
rect 7363 35848 7372 35888
rect 7412 35848 7421 35888
rect 7363 35847 7421 35848
rect 8611 35888 8669 35889
rect 8611 35848 8620 35888
rect 8660 35848 8669 35888
rect 8611 35847 8669 35848
rect 9379 35888 9437 35889
rect 9379 35848 9388 35888
rect 9428 35848 9437 35888
rect 9379 35847 9437 35848
rect 9675 35888 9717 35897
rect 9675 35848 9676 35888
rect 9716 35848 9717 35888
rect 9675 35839 9717 35848
rect 10531 35888 10589 35889
rect 10531 35848 10540 35888
rect 10580 35848 10589 35888
rect 10531 35847 10589 35848
rect 11779 35888 11837 35889
rect 11779 35848 11788 35888
rect 11828 35848 11837 35888
rect 11779 35847 11837 35848
rect 11979 35888 12021 35897
rect 11979 35848 11980 35888
rect 12020 35848 12021 35888
rect 11979 35839 12021 35848
rect 12171 35888 12213 35897
rect 12171 35848 12172 35888
rect 12212 35848 12213 35888
rect 12171 35839 12213 35848
rect 12459 35888 12501 35897
rect 12459 35848 12460 35888
rect 12500 35848 12501 35888
rect 12835 35888 12893 35889
rect 12459 35839 12501 35848
rect 12651 35877 12693 35886
rect 12651 35837 12652 35877
rect 12692 35837 12693 35877
rect 12835 35848 12844 35888
rect 12884 35848 12893 35888
rect 12835 35847 12893 35848
rect 14083 35888 14141 35889
rect 14083 35848 14092 35888
rect 14132 35848 14141 35888
rect 14083 35847 14141 35848
rect 15331 35888 15389 35889
rect 15331 35848 15340 35888
rect 15380 35848 15389 35888
rect 15331 35847 15389 35848
rect 16579 35888 16637 35889
rect 16579 35848 16588 35888
rect 16628 35848 16637 35888
rect 16579 35847 16637 35848
rect 17643 35888 17685 35897
rect 17643 35848 17644 35888
rect 17684 35848 17685 35888
rect 17643 35839 17685 35848
rect 17739 35888 17781 35897
rect 17739 35848 17740 35888
rect 17780 35848 17781 35888
rect 17739 35839 17781 35848
rect 18219 35888 18261 35897
rect 19179 35893 19221 35902
rect 18219 35848 18220 35888
rect 18260 35848 18261 35888
rect 18219 35839 18261 35848
rect 18691 35888 18749 35889
rect 18691 35848 18700 35888
rect 18740 35848 18749 35888
rect 18691 35847 18749 35848
rect 19179 35853 19180 35893
rect 19220 35853 19221 35893
rect 19179 35844 19221 35853
rect 12651 35828 12693 35837
rect 9771 35804 9813 35813
rect 9771 35764 9772 35804
rect 9812 35764 9813 35804
rect 9771 35755 9813 35764
rect 4683 35720 4725 35729
rect 4683 35680 4684 35720
rect 4724 35680 4725 35720
rect 4683 35671 4725 35680
rect 6699 35720 6741 35729
rect 6699 35680 6700 35720
rect 6740 35680 6741 35720
rect 6699 35671 6741 35680
rect 8995 35720 9053 35721
rect 8995 35680 9004 35720
rect 9044 35680 9053 35720
rect 8995 35679 9053 35680
rect 10347 35720 10389 35729
rect 10347 35680 10348 35720
rect 10388 35680 10389 35720
rect 10347 35671 10389 35680
rect 12075 35720 12117 35729
rect 12075 35680 12076 35720
rect 12116 35680 12117 35720
rect 12075 35671 12117 35680
rect 12555 35720 12597 35729
rect 12555 35680 12556 35720
rect 12596 35680 12597 35720
rect 12555 35671 12597 35680
rect 17251 35720 17309 35721
rect 17251 35680 17260 35720
rect 17300 35680 17309 35720
rect 17251 35679 17309 35680
rect 19371 35720 19413 35729
rect 19371 35680 19372 35720
rect 19412 35680 19413 35720
rect 19371 35671 19413 35680
rect 1152 35552 20452 35576
rect 1152 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20452 35552
rect 1152 35488 20452 35512
rect 4299 35300 4341 35309
rect 4299 35260 4300 35300
rect 4340 35260 4341 35300
rect 4299 35251 4341 35260
rect 7563 35300 7605 35309
rect 7563 35260 7564 35300
rect 7604 35260 7605 35300
rect 7563 35251 7605 35260
rect 8235 35300 8277 35309
rect 8235 35260 8236 35300
rect 8276 35260 8277 35300
rect 8235 35251 8277 35260
rect 9771 35300 9813 35309
rect 9771 35260 9772 35300
rect 9812 35260 9813 35300
rect 9771 35251 9813 35260
rect 14571 35300 14613 35309
rect 14571 35260 14572 35300
rect 14612 35260 14613 35300
rect 14571 35251 14613 35260
rect 16395 35300 16437 35309
rect 16395 35260 16396 35300
rect 16436 35260 16437 35300
rect 16395 35251 16437 35260
rect 17547 35300 17589 35309
rect 17547 35260 17548 35300
rect 17588 35260 17589 35300
rect 17547 35251 17589 35260
rect 2571 35216 2613 35225
rect 2571 35176 2572 35216
rect 2612 35176 2613 35216
rect 2571 35167 2613 35176
rect 2667 35216 2709 35225
rect 2667 35176 2668 35216
rect 2708 35176 2709 35216
rect 2667 35167 2709 35176
rect 3619 35216 3677 35217
rect 3619 35176 3628 35216
rect 3668 35176 3677 35216
rect 4779 35216 4821 35225
rect 3619 35175 3677 35176
rect 4107 35202 4149 35211
rect 4107 35162 4108 35202
rect 4148 35162 4149 35202
rect 4779 35176 4780 35216
rect 4820 35176 4821 35216
rect 4779 35167 4821 35176
rect 5067 35216 5109 35225
rect 5067 35176 5068 35216
rect 5108 35176 5109 35216
rect 5067 35167 5109 35176
rect 5259 35216 5301 35225
rect 5259 35176 5260 35216
rect 5300 35176 5301 35216
rect 5259 35167 5301 35176
rect 5451 35216 5493 35225
rect 5451 35176 5452 35216
rect 5492 35176 5493 35216
rect 5451 35167 5493 35176
rect 5539 35216 5597 35217
rect 5539 35176 5548 35216
rect 5588 35176 5597 35216
rect 5539 35175 5597 35176
rect 5835 35216 5877 35225
rect 5835 35176 5836 35216
rect 5876 35176 5877 35216
rect 5835 35167 5877 35176
rect 5931 35216 5973 35225
rect 5931 35176 5932 35216
rect 5972 35176 5973 35216
rect 6883 35216 6941 35217
rect 5931 35167 5973 35176
rect 6315 35174 6357 35183
rect 6883 35176 6892 35216
rect 6932 35176 6941 35216
rect 6883 35175 6941 35176
rect 7371 35211 7413 35220
rect 4107 35153 4149 35162
rect 2083 35132 2141 35133
rect 2083 35092 2092 35132
rect 2132 35092 2141 35132
rect 2083 35091 2141 35092
rect 3051 35132 3093 35141
rect 3051 35092 3052 35132
rect 3092 35092 3093 35132
rect 3051 35083 3093 35092
rect 3147 35132 3189 35141
rect 3147 35092 3148 35132
rect 3188 35092 3189 35132
rect 6315 35134 6316 35174
rect 6356 35134 6357 35174
rect 7371 35171 7372 35211
rect 7412 35171 7413 35211
rect 7843 35216 7901 35217
rect 7843 35176 7852 35216
rect 7892 35176 7901 35216
rect 7843 35175 7901 35176
rect 8139 35216 8181 35225
rect 8139 35176 8140 35216
rect 8180 35176 8181 35216
rect 7371 35162 7413 35171
rect 8139 35167 8181 35176
rect 9379 35216 9437 35217
rect 9379 35176 9388 35216
rect 9428 35176 9437 35216
rect 9379 35175 9437 35176
rect 9675 35216 9717 35225
rect 9675 35176 9676 35216
rect 9716 35176 9717 35216
rect 9675 35167 9717 35176
rect 10251 35216 10293 35225
rect 10251 35176 10252 35216
rect 10292 35176 10293 35216
rect 10251 35167 10293 35176
rect 10339 35216 10397 35217
rect 10339 35176 10348 35216
rect 10388 35176 10397 35216
rect 10339 35175 10397 35176
rect 10531 35216 10589 35217
rect 10531 35176 10540 35216
rect 10580 35176 10589 35216
rect 10531 35175 10589 35176
rect 11779 35216 11837 35217
rect 11779 35176 11788 35216
rect 11828 35176 11837 35216
rect 11779 35175 11837 35176
rect 12171 35216 12213 35225
rect 12171 35176 12172 35216
rect 12212 35176 12213 35216
rect 12171 35167 12213 35176
rect 12363 35216 12405 35225
rect 12363 35176 12364 35216
rect 12404 35176 12405 35216
rect 12363 35167 12405 35176
rect 12451 35216 12509 35217
rect 12451 35176 12460 35216
rect 12500 35176 12509 35216
rect 12451 35175 12509 35176
rect 13123 35216 13181 35217
rect 13123 35176 13132 35216
rect 13172 35176 13181 35216
rect 13123 35175 13181 35176
rect 14371 35216 14429 35217
rect 14371 35176 14380 35216
rect 14420 35176 14429 35216
rect 14371 35175 14429 35176
rect 14947 35216 15005 35217
rect 14947 35176 14956 35216
rect 14996 35176 15005 35216
rect 14947 35175 15005 35176
rect 16195 35216 16253 35217
rect 16195 35176 16204 35216
rect 16244 35176 16253 35216
rect 16195 35175 16253 35176
rect 17731 35216 17789 35217
rect 17731 35176 17740 35216
rect 17780 35176 17789 35216
rect 17731 35175 17789 35176
rect 18979 35216 19037 35217
rect 18979 35176 18988 35216
rect 19028 35176 19037 35216
rect 18979 35175 19037 35176
rect 6315 35125 6357 35134
rect 6411 35132 6453 35141
rect 3147 35083 3189 35092
rect 6411 35092 6412 35132
rect 6452 35092 6453 35132
rect 6411 35083 6453 35092
rect 19459 35132 19517 35133
rect 19459 35092 19468 35132
rect 19508 35092 19517 35132
rect 19459 35091 19517 35092
rect 19843 35132 19901 35133
rect 19843 35092 19852 35132
rect 19892 35092 19901 35132
rect 19843 35091 19901 35092
rect 5259 35048 5301 35057
rect 5259 35008 5260 35048
rect 5300 35008 5301 35048
rect 5259 34999 5301 35008
rect 9003 35048 9045 35057
rect 9003 35008 9004 35048
rect 9044 35008 9045 35048
rect 9003 34999 9045 35008
rect 12843 35048 12885 35057
rect 12843 35008 12844 35048
rect 12884 35008 12885 35048
rect 12843 34999 12885 35008
rect 17259 35048 17301 35057
rect 17259 35008 17260 35048
rect 17300 35008 17301 35048
rect 17259 34999 17301 35008
rect 19659 35048 19701 35057
rect 19659 35008 19660 35048
rect 19700 35008 19701 35048
rect 19659 34999 19701 35008
rect 20043 35048 20085 35057
rect 20043 35008 20044 35048
rect 20084 35008 20085 35048
rect 20043 34999 20085 35008
rect 1899 34964 1941 34973
rect 1899 34924 1900 34964
rect 1940 34924 1941 34964
rect 1899 34915 1941 34924
rect 5067 34964 5109 34973
rect 5067 34924 5068 34964
rect 5108 34924 5109 34964
rect 5067 34915 5109 34924
rect 8515 34964 8573 34965
rect 8515 34924 8524 34964
rect 8564 34924 8573 34964
rect 8515 34923 8573 34924
rect 10051 34964 10109 34965
rect 10051 34924 10060 34964
rect 10100 34924 10109 34964
rect 10051 34923 10109 34924
rect 11979 34964 12021 34973
rect 11979 34924 11980 34964
rect 12020 34924 12021 34964
rect 11979 34915 12021 34924
rect 12171 34964 12213 34973
rect 12171 34924 12172 34964
rect 12212 34924 12213 34964
rect 12171 34915 12213 34924
rect 1152 34796 20352 34820
rect 1152 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 20352 34796
rect 1152 34732 20352 34756
rect 2667 34628 2709 34637
rect 2667 34588 2668 34628
rect 2708 34588 2709 34628
rect 2667 34579 2709 34588
rect 5931 34628 5973 34637
rect 5931 34588 5932 34628
rect 5972 34588 5973 34628
rect 5931 34579 5973 34588
rect 16875 34628 16917 34637
rect 16875 34588 16876 34628
rect 16916 34588 16917 34628
rect 16875 34579 16917 34588
rect 19659 34628 19701 34637
rect 19659 34588 19660 34628
rect 19700 34588 19701 34628
rect 19659 34579 19701 34588
rect 9963 34544 10005 34553
rect 9963 34504 9964 34544
rect 10004 34504 10005 34544
rect 9963 34495 10005 34504
rect 8331 34460 8373 34469
rect 8331 34420 8332 34460
rect 8372 34420 8373 34460
rect 8331 34411 8373 34420
rect 15051 34460 15093 34469
rect 15051 34420 15052 34460
rect 15092 34420 15093 34460
rect 15051 34411 15093 34420
rect 16675 34460 16733 34461
rect 16675 34420 16684 34460
rect 16724 34420 16733 34460
rect 16675 34419 16733 34420
rect 19459 34460 19517 34461
rect 19459 34420 19468 34460
rect 19508 34420 19517 34460
rect 19459 34419 19517 34420
rect 19843 34460 19901 34461
rect 19843 34420 19852 34460
rect 19892 34420 19901 34460
rect 19843 34419 19901 34420
rect 1219 34376 1277 34377
rect 1219 34336 1228 34376
rect 1268 34336 1277 34376
rect 1219 34335 1277 34336
rect 2467 34376 2525 34377
rect 2467 34336 2476 34376
rect 2516 34336 2525 34376
rect 2467 34335 2525 34336
rect 3043 34376 3101 34377
rect 3043 34336 3052 34376
rect 3092 34336 3101 34376
rect 3043 34335 3101 34336
rect 4291 34376 4349 34377
rect 4291 34336 4300 34376
rect 4340 34336 4349 34376
rect 4291 34335 4349 34336
rect 4483 34376 4541 34377
rect 4483 34336 4492 34376
rect 4532 34336 4541 34376
rect 4483 34335 4541 34336
rect 5731 34376 5789 34377
rect 5731 34336 5740 34376
rect 5780 34336 5789 34376
rect 5731 34335 5789 34336
rect 6115 34376 6173 34377
rect 6115 34336 6124 34376
rect 6164 34336 6173 34376
rect 6115 34335 6173 34336
rect 7363 34376 7421 34377
rect 7363 34336 7372 34376
rect 7412 34336 7421 34376
rect 7363 34335 7421 34336
rect 7755 34376 7797 34385
rect 7755 34336 7756 34376
rect 7796 34336 7797 34376
rect 7755 34327 7797 34336
rect 8043 34376 8085 34385
rect 8043 34336 8044 34376
rect 8084 34336 8085 34376
rect 8043 34327 8085 34336
rect 8515 34376 8573 34377
rect 8515 34336 8524 34376
rect 8564 34336 8573 34376
rect 8515 34335 8573 34336
rect 9763 34376 9821 34377
rect 9763 34336 9772 34376
rect 9812 34336 9821 34376
rect 9763 34335 9821 34336
rect 10251 34376 10293 34385
rect 10251 34336 10252 34376
rect 10292 34336 10293 34376
rect 10251 34327 10293 34336
rect 10347 34376 10389 34385
rect 10347 34336 10348 34376
rect 10388 34336 10389 34376
rect 10347 34327 10389 34336
rect 10731 34376 10773 34385
rect 10731 34336 10732 34376
rect 10772 34336 10773 34376
rect 10731 34327 10773 34336
rect 10827 34376 10869 34385
rect 11787 34381 11829 34390
rect 10827 34336 10828 34376
rect 10868 34336 10869 34376
rect 10827 34327 10869 34336
rect 11299 34376 11357 34377
rect 11299 34336 11308 34376
rect 11348 34336 11357 34376
rect 11299 34335 11357 34336
rect 11787 34341 11788 34381
rect 11828 34341 11829 34381
rect 11787 34332 11829 34341
rect 12163 34376 12221 34377
rect 12163 34336 12172 34376
rect 12212 34336 12221 34376
rect 12163 34335 12221 34336
rect 12267 34376 12309 34385
rect 12267 34336 12268 34376
rect 12308 34336 12309 34376
rect 12267 34327 12309 34336
rect 12459 34376 12501 34385
rect 12459 34336 12460 34376
rect 12500 34336 12501 34376
rect 12459 34327 12501 34336
rect 12739 34376 12797 34377
rect 12739 34336 12748 34376
rect 12788 34336 12797 34376
rect 12739 34335 12797 34336
rect 13987 34376 14045 34377
rect 13987 34336 13996 34376
rect 14036 34336 14045 34376
rect 13987 34335 14045 34336
rect 14475 34376 14517 34385
rect 14475 34336 14476 34376
rect 14516 34336 14517 34376
rect 14475 34327 14517 34336
rect 14571 34376 14613 34385
rect 14571 34336 14572 34376
rect 14612 34336 14613 34376
rect 14571 34327 14613 34336
rect 14955 34376 14997 34385
rect 16011 34381 16053 34390
rect 19131 34385 19173 34394
rect 14955 34336 14956 34376
rect 14996 34336 14997 34376
rect 14955 34327 14997 34336
rect 15523 34376 15581 34377
rect 15523 34336 15532 34376
rect 15572 34336 15581 34376
rect 15523 34335 15581 34336
rect 16011 34341 16012 34381
rect 16052 34341 16053 34381
rect 16011 34332 16053 34341
rect 17547 34376 17589 34385
rect 17547 34336 17548 34376
rect 17588 34336 17589 34376
rect 17547 34327 17589 34336
rect 17643 34376 17685 34385
rect 17643 34336 17644 34376
rect 17684 34336 17685 34376
rect 17643 34327 17685 34336
rect 18027 34376 18069 34385
rect 18027 34336 18028 34376
rect 18068 34336 18069 34376
rect 18027 34327 18069 34336
rect 18123 34376 18165 34385
rect 18123 34336 18124 34376
rect 18164 34336 18165 34376
rect 18123 34327 18165 34336
rect 18595 34376 18653 34377
rect 18595 34336 18604 34376
rect 18644 34336 18653 34376
rect 19131 34345 19132 34385
rect 19172 34345 19173 34385
rect 19131 34336 19173 34345
rect 18595 34335 18653 34336
rect 11979 34292 12021 34301
rect 11979 34252 11980 34292
rect 12020 34252 12021 34292
rect 11979 34243 12021 34252
rect 14187 34292 14229 34301
rect 14187 34252 14188 34292
rect 14228 34252 14229 34292
rect 14187 34243 14229 34252
rect 2859 34208 2901 34217
rect 2859 34168 2860 34208
rect 2900 34168 2901 34208
rect 2859 34159 2901 34168
rect 5931 34208 5973 34217
rect 5931 34168 5932 34208
rect 5972 34168 5973 34208
rect 5931 34159 5973 34168
rect 7563 34208 7605 34217
rect 7563 34168 7564 34208
rect 7604 34168 7605 34208
rect 7563 34159 7605 34168
rect 7947 34208 7989 34217
rect 7947 34168 7948 34208
rect 7988 34168 7989 34208
rect 7947 34159 7989 34168
rect 12355 34208 12413 34209
rect 12355 34168 12364 34208
rect 12404 34168 12413 34208
rect 12355 34167 12413 34168
rect 16203 34208 16245 34217
rect 16203 34168 16204 34208
rect 16244 34168 16245 34208
rect 16203 34159 16245 34168
rect 19275 34208 19317 34217
rect 19275 34168 19276 34208
rect 19316 34168 19317 34208
rect 19275 34159 19317 34168
rect 20043 34208 20085 34217
rect 20043 34168 20044 34208
rect 20084 34168 20085 34208
rect 20043 34159 20085 34168
rect 1152 34040 20452 34064
rect 1152 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20452 34040
rect 1152 33976 20452 34000
rect 2859 33872 2901 33881
rect 2859 33832 2860 33872
rect 2900 33832 2901 33872
rect 2859 33823 2901 33832
rect 3243 33872 3285 33881
rect 3243 33832 3244 33872
rect 3284 33832 3285 33872
rect 3243 33823 3285 33832
rect 5251 33872 5309 33873
rect 5251 33832 5260 33872
rect 5300 33832 5309 33872
rect 5251 33831 5309 33832
rect 9763 33872 9821 33873
rect 9763 33832 9772 33872
rect 9812 33832 9821 33872
rect 9763 33831 9821 33832
rect 15915 33872 15957 33881
rect 15915 33832 15916 33872
rect 15956 33832 15957 33872
rect 15915 33823 15957 33832
rect 18603 33872 18645 33881
rect 18603 33832 18604 33872
rect 18644 33832 18645 33872
rect 18603 33823 18645 33832
rect 19563 33872 19605 33881
rect 19563 33832 19564 33872
rect 19604 33832 19605 33872
rect 19563 33823 19605 33832
rect 19947 33872 19989 33881
rect 19947 33832 19948 33872
rect 19988 33832 19989 33872
rect 19947 33823 19989 33832
rect 7563 33788 7605 33797
rect 7563 33748 7564 33788
rect 7604 33748 7605 33788
rect 7563 33739 7605 33748
rect 1219 33704 1277 33705
rect 1219 33664 1228 33704
rect 1268 33664 1277 33704
rect 1219 33663 1277 33664
rect 2467 33704 2525 33705
rect 2467 33664 2476 33704
rect 2516 33664 2525 33704
rect 2467 33663 2525 33664
rect 2947 33704 3005 33705
rect 2947 33664 2956 33704
rect 2996 33664 3005 33704
rect 2947 33663 3005 33664
rect 3435 33699 3477 33708
rect 3435 33659 3436 33699
rect 3476 33659 3477 33699
rect 3907 33704 3965 33705
rect 3907 33664 3916 33704
rect 3956 33664 3965 33704
rect 3907 33663 3965 33664
rect 4875 33704 4917 33713
rect 4875 33664 4876 33704
rect 4916 33664 4917 33704
rect 3435 33650 3477 33659
rect 4875 33655 4917 33664
rect 4971 33704 5013 33713
rect 4971 33664 4972 33704
rect 5012 33664 5013 33704
rect 4971 33655 5013 33664
rect 5355 33704 5397 33713
rect 5355 33664 5356 33704
rect 5396 33664 5397 33704
rect 5355 33655 5397 33664
rect 5451 33704 5493 33713
rect 5451 33664 5452 33704
rect 5492 33664 5493 33704
rect 5451 33655 5493 33664
rect 5547 33704 5589 33713
rect 5547 33664 5548 33704
rect 5588 33664 5589 33704
rect 5547 33655 5589 33664
rect 5835 33704 5877 33713
rect 5835 33664 5836 33704
rect 5876 33664 5877 33704
rect 5835 33655 5877 33664
rect 5931 33704 5973 33713
rect 5931 33664 5932 33704
rect 5972 33664 5973 33704
rect 5931 33655 5973 33664
rect 6883 33704 6941 33705
rect 6883 33664 6892 33704
rect 6932 33664 6941 33704
rect 7747 33704 7805 33705
rect 6883 33663 6941 33664
rect 7419 33694 7461 33703
rect 7419 33654 7420 33694
rect 7460 33654 7461 33694
rect 7747 33664 7756 33704
rect 7796 33664 7805 33704
rect 7747 33663 7805 33664
rect 8995 33704 9053 33705
rect 8995 33664 9004 33704
rect 9044 33664 9053 33704
rect 8995 33663 9053 33664
rect 9483 33704 9525 33713
rect 9483 33664 9484 33704
rect 9524 33664 9525 33704
rect 9483 33655 9525 33664
rect 9579 33704 9621 33713
rect 9579 33664 9580 33704
rect 9620 33664 9621 33704
rect 9579 33655 9621 33664
rect 10819 33704 10877 33705
rect 10819 33664 10828 33704
rect 10868 33664 10877 33704
rect 10819 33663 10877 33664
rect 12067 33704 12125 33705
rect 12067 33664 12076 33704
rect 12116 33664 12125 33704
rect 12067 33663 12125 33664
rect 14083 33704 14141 33705
rect 14083 33664 14092 33704
rect 14132 33664 14141 33704
rect 14083 33663 14141 33664
rect 14467 33704 14525 33705
rect 14467 33664 14476 33704
rect 14516 33664 14525 33704
rect 14467 33663 14525 33664
rect 15715 33704 15773 33705
rect 15715 33664 15724 33704
rect 15764 33664 15773 33704
rect 15715 33663 15773 33664
rect 17155 33704 17213 33705
rect 17155 33664 17164 33704
rect 17204 33664 17213 33704
rect 17155 33663 17213 33664
rect 18403 33704 18461 33705
rect 18403 33664 18412 33704
rect 18452 33664 18461 33704
rect 18403 33663 18461 33664
rect 12835 33662 12893 33663
rect 7419 33645 7461 33654
rect 4395 33620 4437 33629
rect 4395 33580 4396 33620
rect 4436 33580 4437 33620
rect 4395 33571 4437 33580
rect 4491 33620 4533 33629
rect 4491 33580 4492 33620
rect 4532 33580 4533 33620
rect 4491 33571 4533 33580
rect 6315 33620 6357 33629
rect 6315 33580 6316 33620
rect 6356 33580 6357 33620
rect 6315 33571 6357 33580
rect 6411 33620 6453 33629
rect 12835 33622 12844 33662
rect 12884 33622 12893 33662
rect 12835 33621 12893 33622
rect 19374 33633 19432 33634
rect 6411 33580 6412 33620
rect 6452 33580 6453 33620
rect 6411 33571 6453 33580
rect 12451 33620 12509 33621
rect 12451 33580 12460 33620
rect 12500 33580 12509 33620
rect 19374 33593 19383 33633
rect 19423 33593 19432 33633
rect 19374 33592 19432 33593
rect 19747 33620 19805 33621
rect 12451 33579 12509 33580
rect 19747 33580 19756 33620
rect 19796 33580 19805 33620
rect 19747 33579 19805 33580
rect 2667 33452 2709 33461
rect 2667 33412 2668 33452
rect 2708 33412 2709 33452
rect 2667 33403 2709 33412
rect 9195 33452 9237 33461
rect 9195 33412 9196 33452
rect 9236 33412 9237 33452
rect 9195 33403 9237 33412
rect 12267 33452 12309 33461
rect 12267 33412 12268 33452
rect 12308 33412 12309 33452
rect 12267 33403 12309 33412
rect 12651 33452 12693 33461
rect 12651 33412 12652 33452
rect 12692 33412 12693 33452
rect 12651 33403 12693 33412
rect 14283 33452 14325 33461
rect 14283 33412 14284 33452
rect 14324 33412 14325 33452
rect 14283 33403 14325 33412
rect 1152 33284 20352 33308
rect 1152 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 20352 33284
rect 1152 33220 20352 33244
rect 2667 33116 2709 33125
rect 2667 33076 2668 33116
rect 2708 33076 2709 33116
rect 2667 33067 2709 33076
rect 3915 33116 3957 33125
rect 3915 33076 3916 33116
rect 3956 33076 3957 33116
rect 3915 33067 3957 33076
rect 5547 33116 5589 33125
rect 5547 33076 5548 33116
rect 5588 33076 5589 33116
rect 5547 33067 5589 33076
rect 18795 33116 18837 33125
rect 18795 33076 18796 33116
rect 18836 33076 18837 33116
rect 18795 33067 18837 33076
rect 19179 33116 19221 33125
rect 19179 33076 19180 33116
rect 19220 33076 19221 33116
rect 19179 33067 19221 33076
rect 19563 33116 19605 33125
rect 19563 33076 19564 33116
rect 19604 33076 19605 33116
rect 19563 33067 19605 33076
rect 19755 33032 19797 33041
rect 19755 32992 19756 33032
rect 19796 32992 19797 33032
rect 19755 32983 19797 32992
rect 8043 32948 8085 32957
rect 8043 32908 8044 32948
rect 8084 32908 8085 32948
rect 10539 32948 10581 32957
rect 8043 32899 8085 32908
rect 9051 32906 9093 32915
rect 2467 32864 2525 32865
rect 2467 32824 2476 32864
rect 2516 32824 2525 32864
rect 2467 32823 2525 32824
rect 3051 32864 3093 32873
rect 3051 32824 3052 32864
rect 3092 32824 3093 32864
rect 1219 32822 1277 32823
rect 1219 32782 1228 32822
rect 1268 32782 1277 32822
rect 3051 32815 3093 32824
rect 3147 32864 3189 32873
rect 3147 32824 3148 32864
rect 3188 32824 3189 32864
rect 3147 32815 3189 32824
rect 3373 32871 3415 32880
rect 3373 32831 3374 32871
rect 3414 32831 3415 32871
rect 3373 32822 3415 32831
rect 3531 32864 3573 32873
rect 3531 32824 3532 32864
rect 3572 32824 3573 32864
rect 3531 32815 3573 32824
rect 3627 32864 3669 32873
rect 3627 32824 3628 32864
rect 3668 32824 3669 32864
rect 3627 32815 3669 32824
rect 3811 32864 3869 32865
rect 3811 32824 3820 32864
rect 3860 32824 3869 32864
rect 3811 32823 3869 32824
rect 3907 32864 3965 32865
rect 3907 32824 3916 32864
rect 3956 32824 3965 32864
rect 3907 32823 3965 32824
rect 4099 32864 4157 32865
rect 4099 32824 4108 32864
rect 4148 32824 4157 32864
rect 4099 32823 4157 32824
rect 5347 32864 5405 32865
rect 5347 32824 5356 32864
rect 5396 32824 5405 32864
rect 5347 32823 5405 32824
rect 5731 32864 5789 32865
rect 5731 32824 5740 32864
rect 5780 32824 5789 32864
rect 5731 32823 5789 32824
rect 6979 32864 7037 32865
rect 6979 32824 6988 32864
rect 7028 32824 7037 32864
rect 6979 32823 7037 32824
rect 7467 32864 7509 32873
rect 7467 32824 7468 32864
rect 7508 32824 7509 32864
rect 7467 32815 7509 32824
rect 7563 32864 7605 32873
rect 7563 32824 7564 32864
rect 7604 32824 7605 32864
rect 7563 32815 7605 32824
rect 7947 32864 7989 32873
rect 9051 32866 9052 32906
rect 9092 32866 9093 32906
rect 10539 32908 10540 32948
rect 10580 32908 10581 32948
rect 10539 32899 10581 32908
rect 10635 32948 10677 32957
rect 10635 32908 10636 32948
rect 10676 32908 10677 32948
rect 10635 32899 10677 32908
rect 17163 32948 17205 32957
rect 17163 32908 17164 32948
rect 17204 32908 17205 32948
rect 13603 32906 13661 32907
rect 7947 32824 7948 32864
rect 7988 32824 7989 32864
rect 7947 32815 7989 32824
rect 8515 32864 8573 32865
rect 8515 32824 8524 32864
rect 8564 32824 8573 32864
rect 9051 32857 9093 32866
rect 10059 32864 10101 32873
rect 8515 32823 8573 32824
rect 10059 32824 10060 32864
rect 10100 32824 10101 32864
rect 10059 32815 10101 32824
rect 10155 32864 10197 32873
rect 11595 32869 11637 32878
rect 10155 32824 10156 32864
rect 10196 32824 10197 32864
rect 10155 32815 10197 32824
rect 11107 32864 11165 32865
rect 11107 32824 11116 32864
rect 11156 32824 11165 32864
rect 11107 32823 11165 32824
rect 11595 32829 11596 32869
rect 11636 32829 11637 32869
rect 13603 32866 13612 32906
rect 13652 32866 13661 32906
rect 17163 32899 17205 32908
rect 17259 32948 17301 32957
rect 17259 32908 17260 32948
rect 17300 32908 17301 32948
rect 17259 32899 17301 32908
rect 18595 32948 18653 32949
rect 18595 32908 18604 32948
rect 18644 32908 18653 32948
rect 18595 32907 18653 32908
rect 18979 32948 19037 32949
rect 18979 32908 18988 32948
rect 19028 32908 19037 32948
rect 18979 32907 19037 32908
rect 19363 32948 19421 32949
rect 19363 32908 19372 32948
rect 19412 32908 19421 32948
rect 19363 32907 19421 32908
rect 20035 32948 20093 32949
rect 20035 32908 20044 32948
rect 20084 32908 20093 32948
rect 20035 32907 20093 32908
rect 13603 32865 13661 32866
rect 14851 32885 14909 32886
rect 11595 32820 11637 32829
rect 11971 32864 12029 32865
rect 11971 32824 11980 32864
rect 12020 32824 12029 32864
rect 11971 32823 12029 32824
rect 13219 32864 13277 32865
rect 13219 32824 13228 32864
rect 13268 32824 13277 32864
rect 14851 32845 14860 32885
rect 14900 32845 14909 32885
rect 18219 32878 18261 32887
rect 14851 32844 14909 32845
rect 16683 32864 16725 32873
rect 13219 32823 13277 32824
rect 16683 32824 16684 32864
rect 16724 32824 16725 32864
rect 16683 32815 16725 32824
rect 16779 32864 16821 32873
rect 16779 32824 16780 32864
rect 16820 32824 16821 32864
rect 16779 32815 16821 32824
rect 17731 32864 17789 32865
rect 17731 32824 17740 32864
rect 17780 32824 17789 32864
rect 18219 32838 18220 32878
rect 18260 32838 18261 32878
rect 18219 32829 18261 32838
rect 17731 32823 17789 32824
rect 1219 32781 1277 32782
rect 7179 32780 7221 32789
rect 7179 32740 7180 32780
rect 7220 32740 7221 32780
rect 7179 32731 7221 32740
rect 11787 32780 11829 32789
rect 11787 32740 11788 32780
rect 11828 32740 11829 32780
rect 11787 32731 11829 32740
rect 18411 32780 18453 32789
rect 18411 32740 18412 32780
rect 18452 32740 18453 32780
rect 18411 32731 18453 32740
rect 2851 32696 2909 32697
rect 2851 32656 2860 32696
rect 2900 32656 2909 32696
rect 2851 32655 2909 32656
rect 9195 32696 9237 32705
rect 9195 32656 9196 32696
rect 9236 32656 9237 32696
rect 9195 32647 9237 32656
rect 13419 32696 13461 32705
rect 13419 32656 13420 32696
rect 13460 32656 13461 32696
rect 13419 32647 13461 32656
rect 15051 32696 15093 32705
rect 15051 32656 15052 32696
rect 15092 32656 15093 32696
rect 15051 32647 15093 32656
rect 20235 32696 20277 32705
rect 20235 32656 20236 32696
rect 20276 32656 20277 32696
rect 20235 32647 20277 32656
rect 1152 32528 20452 32552
rect 1152 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20452 32528
rect 1152 32464 20452 32488
rect 2667 32360 2709 32369
rect 2667 32320 2668 32360
rect 2708 32320 2709 32360
rect 2667 32311 2709 32320
rect 4299 32360 4341 32369
rect 4299 32320 4300 32360
rect 4340 32320 4341 32360
rect 4299 32311 4341 32320
rect 4971 32360 5013 32369
rect 4971 32320 4972 32360
rect 5012 32320 5013 32360
rect 4971 32311 5013 32320
rect 8035 32360 8093 32361
rect 8035 32320 8044 32360
rect 8084 32320 8093 32360
rect 8035 32319 8093 32320
rect 9867 32360 9909 32369
rect 9867 32320 9868 32360
rect 9908 32320 9909 32360
rect 9867 32311 9909 32320
rect 11595 32360 11637 32369
rect 11595 32320 11596 32360
rect 11636 32320 11637 32360
rect 11595 32311 11637 32320
rect 11971 32360 12029 32361
rect 11971 32320 11980 32360
rect 12020 32320 12029 32360
rect 11971 32319 12029 32320
rect 12739 32360 12797 32361
rect 12739 32320 12748 32360
rect 12788 32320 12797 32360
rect 12739 32319 12797 32320
rect 17163 32360 17205 32369
rect 17163 32320 17164 32360
rect 17204 32320 17205 32360
rect 17163 32311 17205 32320
rect 20235 32360 20277 32369
rect 20235 32320 20236 32360
rect 20276 32320 20277 32360
rect 20235 32311 20277 32320
rect 14955 32276 14997 32285
rect 14955 32236 14956 32276
rect 14996 32236 14997 32276
rect 14955 32227 14997 32236
rect 16971 32276 17013 32285
rect 16971 32236 16972 32276
rect 17012 32236 17013 32276
rect 16971 32227 17013 32236
rect 1219 32192 1277 32193
rect 1219 32152 1228 32192
rect 1268 32152 1277 32192
rect 1219 32151 1277 32152
rect 2467 32192 2525 32193
rect 2467 32152 2476 32192
rect 2516 32152 2525 32192
rect 2467 32151 2525 32152
rect 2851 32192 2909 32193
rect 2851 32152 2860 32192
rect 2900 32152 2909 32192
rect 2851 32151 2909 32152
rect 4099 32192 4157 32193
rect 4099 32152 4108 32192
rect 4148 32152 4157 32192
rect 4099 32151 4157 32152
rect 4491 32192 4533 32201
rect 4491 32152 4492 32192
rect 4532 32152 4533 32192
rect 4491 32143 4533 32152
rect 4587 32192 4629 32201
rect 4587 32152 4588 32192
rect 4628 32152 4629 32192
rect 4587 32143 4629 32152
rect 4779 32192 4821 32201
rect 4779 32152 4780 32192
rect 4820 32152 4821 32192
rect 4779 32143 4821 32152
rect 5059 32192 5117 32193
rect 5059 32152 5068 32192
rect 5108 32152 5117 32192
rect 5059 32151 5117 32152
rect 7755 32192 7797 32201
rect 7755 32152 7756 32192
rect 7796 32152 7797 32192
rect 7755 32143 7797 32152
rect 7851 32192 7893 32201
rect 7851 32152 7852 32192
rect 7892 32152 7893 32192
rect 7851 32143 7893 32152
rect 8419 32192 8477 32193
rect 8419 32152 8428 32192
rect 8468 32152 8477 32192
rect 8419 32151 8477 32152
rect 9667 32192 9725 32193
rect 9667 32152 9676 32192
rect 9716 32152 9725 32192
rect 9667 32151 9725 32152
rect 10147 32192 10205 32193
rect 10147 32152 10156 32192
rect 10196 32152 10205 32192
rect 10147 32151 10205 32152
rect 11395 32192 11453 32193
rect 11395 32152 11404 32192
rect 11444 32152 11453 32192
rect 11395 32151 11453 32152
rect 12459 32192 12501 32201
rect 12459 32152 12460 32192
rect 12500 32152 12501 32192
rect 12459 32143 12501 32152
rect 12555 32192 12597 32201
rect 12555 32152 12556 32192
rect 12596 32152 12597 32192
rect 12555 32143 12597 32152
rect 13227 32192 13269 32201
rect 13227 32152 13228 32192
rect 13268 32152 13269 32192
rect 13227 32143 13269 32152
rect 13323 32192 13365 32201
rect 13323 32152 13324 32192
rect 13364 32152 13365 32192
rect 13323 32143 13365 32152
rect 13707 32192 13749 32201
rect 13707 32152 13708 32192
rect 13748 32152 13749 32192
rect 13707 32143 13749 32152
rect 13803 32192 13845 32201
rect 13803 32152 13804 32192
rect 13844 32152 13845 32192
rect 13803 32143 13845 32152
rect 14275 32192 14333 32193
rect 14275 32152 14284 32192
rect 14324 32152 14333 32192
rect 15243 32192 15285 32201
rect 14275 32151 14333 32152
rect 14811 32182 14853 32191
rect 14811 32142 14812 32182
rect 14852 32142 14853 32182
rect 15243 32152 15244 32192
rect 15284 32152 15285 32192
rect 15243 32143 15285 32152
rect 15339 32192 15381 32201
rect 15339 32152 15340 32192
rect 15380 32152 15381 32192
rect 15339 32143 15381 32152
rect 15723 32192 15765 32201
rect 15723 32152 15724 32192
rect 15764 32152 15765 32192
rect 15723 32143 15765 32152
rect 15819 32192 15861 32201
rect 15819 32152 15820 32192
rect 15860 32152 15861 32192
rect 15819 32143 15861 32152
rect 16291 32192 16349 32193
rect 16291 32152 16300 32192
rect 16340 32152 16349 32192
rect 17347 32192 17405 32193
rect 16291 32151 16349 32152
rect 16779 32178 16821 32187
rect 14811 32133 14853 32142
rect 16779 32138 16780 32178
rect 16820 32138 16821 32178
rect 17347 32152 17356 32192
rect 17396 32152 17405 32192
rect 17347 32151 17405 32152
rect 18595 32192 18653 32193
rect 18595 32152 18604 32192
rect 18644 32152 18653 32192
rect 18595 32151 18653 32152
rect 18787 32192 18845 32193
rect 18787 32152 18796 32192
rect 18836 32152 18845 32192
rect 18787 32151 18845 32152
rect 20035 32192 20093 32193
rect 20035 32152 20044 32192
rect 20084 32152 20093 32192
rect 20035 32151 20093 32152
rect 16779 32129 16821 32138
rect 4483 32024 4541 32025
rect 4483 31984 4492 32024
rect 4532 31984 4541 32024
rect 4483 31983 4541 31984
rect 1152 31772 20352 31796
rect 1152 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 20352 31772
rect 1152 31708 20352 31732
rect 5443 31520 5501 31521
rect 5443 31480 5452 31520
rect 5492 31480 5501 31520
rect 5443 31479 5501 31480
rect 13131 31520 13173 31529
rect 13131 31480 13132 31520
rect 13172 31480 13173 31520
rect 13131 31471 13173 31480
rect 14763 31520 14805 31529
rect 14763 31480 14764 31520
rect 14804 31480 14805 31520
rect 14763 31471 14805 31480
rect 16971 31520 17013 31529
rect 16971 31480 16972 31520
rect 17012 31480 17013 31520
rect 16971 31471 17013 31480
rect 19947 31520 19989 31529
rect 19947 31480 19948 31520
rect 19988 31480 19989 31520
rect 19947 31471 19989 31480
rect 2955 31436 2997 31445
rect 2955 31396 2956 31436
rect 2996 31396 2997 31436
rect 2955 31387 2997 31396
rect 4291 31436 4349 31437
rect 4291 31396 4300 31436
rect 4340 31396 4349 31436
rect 4291 31395 4349 31396
rect 11211 31436 11253 31445
rect 11211 31396 11212 31436
rect 11252 31396 11253 31436
rect 17739 31436 17781 31445
rect 11211 31387 11253 31396
rect 12219 31394 12261 31403
rect 3963 31361 4005 31370
rect 2379 31352 2421 31361
rect 2379 31312 2380 31352
rect 2420 31312 2421 31352
rect 2379 31303 2421 31312
rect 2475 31352 2517 31361
rect 2475 31312 2476 31352
rect 2516 31312 2517 31352
rect 2475 31303 2517 31312
rect 2859 31352 2901 31361
rect 2859 31312 2860 31352
rect 2900 31312 2901 31352
rect 2859 31303 2901 31312
rect 3427 31352 3485 31353
rect 3427 31312 3436 31352
rect 3476 31312 3485 31352
rect 3963 31321 3964 31361
rect 4004 31321 4005 31361
rect 3963 31312 4005 31321
rect 4771 31352 4829 31353
rect 4771 31312 4780 31352
rect 4820 31312 4829 31352
rect 3427 31311 3485 31312
rect 4771 31311 4829 31312
rect 5067 31352 5109 31361
rect 5067 31312 5068 31352
rect 5108 31312 5109 31352
rect 5067 31303 5109 31312
rect 5635 31352 5693 31353
rect 5635 31312 5644 31352
rect 5684 31312 5693 31352
rect 5635 31311 5693 31312
rect 6883 31352 6941 31353
rect 6883 31312 6892 31352
rect 6932 31312 6941 31352
rect 6883 31311 6941 31312
rect 7267 31352 7325 31353
rect 7267 31312 7276 31352
rect 7316 31312 7325 31352
rect 7267 31311 7325 31312
rect 8515 31352 8573 31353
rect 8515 31312 8524 31352
rect 8564 31312 8573 31352
rect 8515 31311 8573 31312
rect 8899 31352 8957 31353
rect 8899 31312 8908 31352
rect 8948 31312 8957 31352
rect 8899 31311 8957 31312
rect 10147 31352 10205 31353
rect 10147 31312 10156 31352
rect 10196 31312 10205 31352
rect 10147 31311 10205 31312
rect 10635 31352 10677 31361
rect 10635 31312 10636 31352
rect 10676 31312 10677 31352
rect 10635 31303 10677 31312
rect 10731 31352 10773 31361
rect 10731 31312 10732 31352
rect 10772 31312 10773 31352
rect 10731 31303 10773 31312
rect 11115 31352 11157 31361
rect 12219 31354 12220 31394
rect 12260 31354 12261 31394
rect 17739 31396 17740 31436
rect 17780 31396 17781 31436
rect 17739 31387 17781 31396
rect 19363 31436 19421 31437
rect 19363 31396 19372 31436
rect 19412 31396 19421 31436
rect 19363 31395 19421 31396
rect 19747 31436 19805 31437
rect 19747 31396 19756 31436
rect 19796 31396 19805 31436
rect 19747 31395 19805 31396
rect 11115 31312 11116 31352
rect 11156 31312 11157 31352
rect 11115 31303 11157 31312
rect 11683 31352 11741 31353
rect 11683 31312 11692 31352
rect 11732 31312 11741 31352
rect 12219 31345 12261 31354
rect 13315 31352 13373 31353
rect 11683 31311 11741 31312
rect 13315 31312 13324 31352
rect 13364 31312 13373 31352
rect 13315 31311 13373 31312
rect 14563 31352 14621 31353
rect 14563 31312 14572 31352
rect 14612 31312 14621 31352
rect 14563 31311 14621 31312
rect 15523 31352 15581 31353
rect 15523 31312 15532 31352
rect 15572 31312 15581 31352
rect 15523 31311 15581 31312
rect 16771 31352 16829 31353
rect 16771 31312 16780 31352
rect 16820 31312 16829 31352
rect 16771 31311 16829 31312
rect 17259 31352 17301 31361
rect 17259 31312 17260 31352
rect 17300 31312 17301 31352
rect 17259 31303 17301 31312
rect 17355 31352 17397 31361
rect 17355 31312 17356 31352
rect 17396 31312 17397 31352
rect 17355 31303 17397 31312
rect 17835 31352 17877 31361
rect 18795 31357 18837 31366
rect 17835 31312 17836 31352
rect 17876 31312 17877 31352
rect 17835 31303 17877 31312
rect 18307 31352 18365 31353
rect 18307 31312 18316 31352
rect 18356 31312 18365 31352
rect 18307 31311 18365 31312
rect 18795 31317 18796 31357
rect 18836 31317 18837 31357
rect 18795 31308 18837 31317
rect 4107 31268 4149 31277
rect 4107 31228 4108 31268
rect 4148 31228 4149 31268
rect 4107 31219 4149 31228
rect 5163 31268 5205 31277
rect 5163 31228 5164 31268
rect 5204 31228 5205 31268
rect 5163 31219 5205 31228
rect 10347 31268 10389 31277
rect 10347 31228 10348 31268
rect 10388 31228 10389 31268
rect 10347 31219 10389 31228
rect 4491 31184 4533 31193
rect 4491 31144 4492 31184
rect 4532 31144 4533 31184
rect 4491 31135 4533 31144
rect 7083 31184 7125 31193
rect 7083 31144 7084 31184
rect 7124 31144 7125 31184
rect 7083 31135 7125 31144
rect 8715 31184 8757 31193
rect 8715 31144 8716 31184
rect 8756 31144 8757 31184
rect 8715 31135 8757 31144
rect 12363 31184 12405 31193
rect 12363 31144 12364 31184
rect 12404 31144 12405 31184
rect 12363 31135 12405 31144
rect 13027 31184 13085 31185
rect 13027 31144 13036 31184
rect 13076 31144 13085 31184
rect 13027 31143 13085 31144
rect 18987 31184 19029 31193
rect 18987 31144 18988 31184
rect 19028 31144 19029 31184
rect 18987 31135 19029 31144
rect 19563 31184 19605 31193
rect 19563 31144 19564 31184
rect 19604 31144 19605 31184
rect 19563 31135 19605 31144
rect 1152 31016 20452 31040
rect 1152 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20452 31016
rect 1152 30952 20452 30976
rect 1803 30848 1845 30857
rect 1803 30808 1804 30848
rect 1844 30808 1845 30848
rect 1803 30799 1845 30808
rect 14763 30848 14805 30857
rect 14763 30808 14764 30848
rect 14804 30808 14805 30848
rect 14763 30799 14805 30808
rect 16395 30848 16437 30857
rect 16395 30808 16396 30848
rect 16436 30808 16437 30848
rect 16395 30799 16437 30808
rect 17355 30848 17397 30857
rect 17355 30808 17356 30848
rect 17396 30808 17397 30848
rect 17355 30799 17397 30808
rect 19275 30848 19317 30857
rect 19275 30808 19276 30848
rect 19316 30808 19317 30848
rect 19275 30799 19317 30808
rect 19659 30848 19701 30857
rect 19659 30808 19660 30848
rect 19700 30808 19701 30848
rect 19659 30799 19701 30808
rect 6795 30764 6837 30773
rect 6795 30724 6796 30764
rect 6836 30724 6837 30764
rect 6795 30715 6837 30724
rect 9387 30764 9429 30773
rect 9387 30724 9388 30764
rect 9428 30724 9429 30764
rect 9387 30715 9429 30724
rect 12363 30764 12405 30773
rect 12363 30724 12364 30764
rect 12404 30724 12405 30764
rect 12363 30715 12405 30724
rect 3331 30680 3389 30681
rect 3331 30640 3340 30680
rect 3380 30640 3389 30680
rect 3331 30639 3389 30640
rect 4579 30680 4637 30681
rect 4579 30640 4588 30680
rect 4628 30640 4637 30680
rect 4579 30639 4637 30640
rect 5067 30680 5109 30689
rect 5067 30640 5068 30680
rect 5108 30640 5109 30680
rect 5067 30631 5109 30640
rect 5163 30680 5205 30689
rect 5163 30640 5164 30680
rect 5204 30640 5205 30680
rect 5163 30631 5205 30640
rect 6115 30680 6173 30681
rect 6115 30640 6124 30680
rect 6164 30640 6173 30680
rect 6987 30680 7029 30689
rect 6115 30639 6173 30640
rect 6603 30666 6645 30675
rect 6603 30626 6604 30666
rect 6644 30626 6645 30666
rect 6987 30640 6988 30680
rect 7028 30640 7029 30680
rect 6987 30631 7029 30640
rect 7083 30680 7125 30689
rect 7083 30640 7084 30680
rect 7124 30640 7125 30680
rect 7083 30631 7125 30640
rect 7179 30680 7221 30689
rect 7179 30640 7180 30680
rect 7220 30640 7221 30680
rect 7179 30631 7221 30640
rect 7275 30680 7317 30689
rect 7275 30640 7276 30680
rect 7316 30640 7317 30680
rect 7275 30631 7317 30640
rect 7659 30680 7701 30689
rect 7659 30640 7660 30680
rect 7700 30640 7701 30680
rect 8139 30680 8181 30689
rect 7659 30631 7701 30640
rect 7755 30661 7797 30670
rect 6603 30617 6645 30626
rect 7755 30621 7756 30661
rect 7796 30621 7797 30661
rect 8139 30640 8140 30680
rect 8180 30640 8181 30680
rect 8139 30631 8181 30640
rect 8707 30680 8765 30681
rect 8707 30640 8716 30680
rect 8756 30640 8765 30680
rect 8707 30639 8765 30640
rect 9195 30675 9237 30684
rect 9195 30635 9196 30675
rect 9236 30635 9237 30675
rect 9195 30626 9237 30635
rect 10635 30680 10677 30689
rect 10635 30640 10636 30680
rect 10676 30640 10677 30680
rect 10635 30631 10677 30640
rect 10731 30680 10773 30689
rect 10731 30640 10732 30680
rect 10772 30640 10773 30680
rect 10731 30631 10773 30640
rect 11115 30680 11157 30689
rect 11115 30640 11116 30680
rect 11156 30640 11157 30680
rect 11115 30631 11157 30640
rect 11211 30680 11253 30689
rect 11211 30640 11212 30680
rect 11252 30640 11253 30680
rect 11211 30631 11253 30640
rect 11683 30680 11741 30681
rect 11683 30640 11692 30680
rect 11732 30640 11741 30680
rect 13315 30680 13373 30681
rect 11683 30639 11741 30640
rect 12219 30638 12261 30647
rect 13315 30640 13324 30680
rect 13364 30640 13373 30680
rect 13315 30639 13373 30640
rect 14563 30680 14621 30681
rect 14563 30640 14572 30680
rect 14612 30640 14621 30680
rect 14563 30639 14621 30640
rect 14947 30680 15005 30681
rect 14947 30640 14956 30680
rect 14996 30640 15005 30680
rect 14947 30639 15005 30640
rect 16195 30680 16253 30681
rect 16195 30640 16204 30680
rect 16244 30640 16253 30680
rect 16195 30639 16253 30640
rect 17827 30680 17885 30681
rect 17827 30640 17836 30680
rect 17876 30640 17885 30680
rect 17827 30639 17885 30640
rect 19075 30680 19133 30681
rect 19075 30640 19084 30680
rect 19124 30640 19133 30680
rect 19075 30639 19133 30640
rect 7755 30612 7797 30621
rect 5547 30596 5589 30605
rect 5547 30556 5548 30596
rect 5588 30556 5589 30596
rect 5547 30547 5589 30556
rect 5643 30596 5685 30605
rect 5643 30556 5644 30596
rect 5684 30556 5685 30596
rect 5643 30547 5685 30556
rect 8235 30596 8277 30605
rect 8235 30556 8236 30596
rect 8276 30556 8277 30596
rect 12219 30598 12220 30638
rect 12260 30598 12261 30638
rect 12219 30589 12261 30598
rect 16771 30596 16829 30597
rect 8235 30547 8277 30556
rect 16771 30556 16780 30596
rect 16820 30556 16829 30596
rect 16771 30555 16829 30556
rect 17155 30596 17213 30597
rect 17155 30556 17164 30596
rect 17204 30556 17213 30596
rect 17155 30555 17213 30556
rect 19459 30596 19517 30597
rect 19459 30556 19468 30596
rect 19508 30556 19517 30596
rect 19459 30555 19517 30556
rect 19843 30596 19901 30597
rect 19843 30556 19852 30596
rect 19892 30556 19901 30596
rect 19843 30555 19901 30556
rect 4779 30428 4821 30437
rect 4779 30388 4780 30428
rect 4820 30388 4821 30428
rect 4779 30379 4821 30388
rect 16971 30428 17013 30437
rect 16971 30388 16972 30428
rect 17012 30388 17013 30428
rect 16971 30379 17013 30388
rect 20043 30428 20085 30437
rect 20043 30388 20044 30428
rect 20084 30388 20085 30428
rect 20043 30379 20085 30388
rect 1152 30260 20352 30284
rect 1152 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 20352 30260
rect 1152 30196 20352 30220
rect 3435 30092 3477 30101
rect 3435 30052 3436 30092
rect 3476 30052 3477 30092
rect 3435 30043 3477 30052
rect 6211 30092 6269 30093
rect 6211 30052 6220 30092
rect 6260 30052 6269 30092
rect 6211 30051 6269 30052
rect 6411 30092 6453 30101
rect 6411 30052 6412 30092
rect 6452 30052 6453 30092
rect 6411 30043 6453 30052
rect 10539 30092 10581 30101
rect 10539 30052 10540 30092
rect 10580 30052 10581 30092
rect 10539 30043 10581 30052
rect 12459 30092 12501 30101
rect 12459 30052 12460 30092
rect 12500 30052 12501 30092
rect 12459 30043 12501 30052
rect 19851 30092 19893 30101
rect 19851 30052 19852 30092
rect 19892 30052 19893 30092
rect 19851 30043 19893 30052
rect 20235 30092 20277 30101
rect 20235 30052 20236 30092
rect 20276 30052 20277 30092
rect 20235 30043 20277 30052
rect 1803 30008 1845 30017
rect 1803 29968 1804 30008
rect 1844 29968 1845 30008
rect 1803 29959 1845 29968
rect 14859 29924 14901 29933
rect 14859 29884 14860 29924
rect 14900 29884 14901 29924
rect 14859 29875 14901 29884
rect 16771 29924 16829 29925
rect 16771 29884 16780 29924
rect 16820 29884 16829 29924
rect 16771 29883 16829 29884
rect 17155 29924 17213 29925
rect 17155 29884 17164 29924
rect 17204 29884 17213 29924
rect 17155 29883 17213 29884
rect 18219 29924 18261 29933
rect 18219 29884 18220 29924
rect 18260 29884 18261 29924
rect 18219 29875 18261 29884
rect 19651 29924 19709 29925
rect 19651 29884 19660 29924
rect 19700 29884 19709 29924
rect 19651 29883 19709 29884
rect 20035 29924 20093 29925
rect 20035 29884 20044 29924
rect 20084 29884 20093 29924
rect 20035 29883 20093 29884
rect 1987 29840 2045 29841
rect 1987 29800 1996 29840
rect 2036 29800 2045 29840
rect 1987 29799 2045 29800
rect 3235 29840 3293 29841
rect 3235 29800 3244 29840
rect 3284 29800 3293 29840
rect 3235 29799 3293 29800
rect 3723 29840 3765 29849
rect 3723 29800 3724 29840
rect 3764 29800 3765 29840
rect 3723 29791 3765 29800
rect 3819 29840 3861 29849
rect 3819 29800 3820 29840
rect 3860 29800 3861 29840
rect 3819 29791 3861 29800
rect 3915 29840 3957 29849
rect 3915 29800 3916 29840
rect 3956 29800 3957 29840
rect 3915 29791 3957 29800
rect 4099 29840 4157 29841
rect 4099 29800 4108 29840
rect 4148 29800 4157 29840
rect 4099 29799 4157 29800
rect 5347 29840 5405 29841
rect 5347 29800 5356 29840
rect 5396 29800 5405 29840
rect 5347 29799 5405 29800
rect 5835 29840 5877 29849
rect 5835 29800 5836 29840
rect 5876 29800 5877 29840
rect 5835 29791 5877 29800
rect 5931 29840 5973 29849
rect 5931 29800 5932 29840
rect 5972 29800 5973 29840
rect 5931 29791 5973 29800
rect 6027 29840 6069 29849
rect 6027 29800 6028 29840
rect 6068 29800 6069 29840
rect 6027 29791 6069 29800
rect 6499 29840 6557 29841
rect 6499 29800 6508 29840
rect 6548 29800 6557 29840
rect 6499 29799 6557 29800
rect 7267 29840 7325 29841
rect 7267 29800 7276 29840
rect 7316 29800 7325 29840
rect 7267 29799 7325 29800
rect 8515 29840 8573 29841
rect 8515 29800 8524 29840
rect 8564 29800 8573 29840
rect 8515 29799 8573 29800
rect 9091 29840 9149 29841
rect 9091 29800 9100 29840
rect 9140 29800 9149 29840
rect 9091 29799 9149 29800
rect 10339 29840 10397 29841
rect 10339 29800 10348 29840
rect 10388 29800 10397 29840
rect 10339 29799 10397 29800
rect 11011 29840 11069 29841
rect 11011 29800 11020 29840
rect 11060 29800 11069 29840
rect 11011 29799 11069 29800
rect 12259 29840 12317 29841
rect 12259 29800 12268 29840
rect 12308 29800 12317 29840
rect 12259 29799 12317 29800
rect 13699 29840 13757 29841
rect 13699 29800 13708 29840
rect 13748 29800 13757 29840
rect 13699 29799 13757 29800
rect 13803 29840 13845 29849
rect 13803 29800 13804 29840
rect 13844 29800 13845 29840
rect 13803 29791 13845 29800
rect 13995 29840 14037 29849
rect 13995 29800 13996 29840
rect 14036 29800 14037 29840
rect 13995 29791 14037 29800
rect 14283 29840 14325 29849
rect 14283 29800 14284 29840
rect 14324 29800 14325 29840
rect 14283 29791 14325 29800
rect 14379 29840 14421 29849
rect 14379 29800 14380 29840
rect 14420 29800 14421 29840
rect 14379 29791 14421 29800
rect 14763 29840 14805 29849
rect 15819 29845 15861 29854
rect 19227 29849 19269 29858
rect 14763 29800 14764 29840
rect 14804 29800 14805 29840
rect 14763 29791 14805 29800
rect 15331 29840 15389 29841
rect 15331 29800 15340 29840
rect 15380 29800 15389 29840
rect 15331 29799 15389 29800
rect 15819 29805 15820 29845
rect 15860 29805 15861 29845
rect 15819 29796 15861 29805
rect 17643 29840 17685 29849
rect 17643 29800 17644 29840
rect 17684 29800 17685 29840
rect 17643 29791 17685 29800
rect 17739 29840 17781 29849
rect 17739 29800 17740 29840
rect 17780 29800 17781 29840
rect 17739 29791 17781 29800
rect 18123 29840 18165 29849
rect 18123 29800 18124 29840
rect 18164 29800 18165 29840
rect 18123 29791 18165 29800
rect 18691 29840 18749 29841
rect 18691 29800 18700 29840
rect 18740 29800 18749 29840
rect 19227 29809 19228 29849
rect 19268 29809 19269 29849
rect 19227 29800 19269 29809
rect 18691 29799 18749 29800
rect 5547 29756 5589 29765
rect 5547 29716 5548 29756
rect 5588 29716 5589 29756
rect 5547 29707 5589 29716
rect 13899 29756 13941 29765
rect 13899 29716 13900 29756
rect 13940 29716 13941 29756
rect 13899 29707 13941 29716
rect 3619 29672 3677 29673
rect 3619 29632 3628 29672
rect 3668 29632 3677 29672
rect 3619 29631 3677 29632
rect 8715 29672 8757 29681
rect 8715 29632 8716 29672
rect 8756 29632 8757 29672
rect 8715 29623 8757 29632
rect 16011 29672 16053 29681
rect 16011 29632 16012 29672
rect 16052 29632 16053 29672
rect 16011 29623 16053 29632
rect 16971 29672 17013 29681
rect 16971 29632 16972 29672
rect 17012 29632 17013 29672
rect 16971 29623 17013 29632
rect 17355 29672 17397 29681
rect 17355 29632 17356 29672
rect 17396 29632 17397 29672
rect 17355 29623 17397 29632
rect 19371 29672 19413 29681
rect 19371 29632 19372 29672
rect 19412 29632 19413 29672
rect 19371 29623 19413 29632
rect 1152 29504 20452 29528
rect 1152 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20452 29504
rect 1152 29440 20452 29464
rect 1803 29336 1845 29345
rect 1803 29296 1804 29336
rect 1844 29296 1845 29336
rect 1803 29287 1845 29296
rect 1987 29336 2045 29337
rect 1987 29296 1996 29336
rect 2036 29296 2045 29336
rect 1987 29295 2045 29296
rect 4771 29336 4829 29337
rect 4771 29296 4780 29336
rect 4820 29296 4829 29336
rect 4771 29295 4829 29296
rect 4963 29336 5021 29337
rect 4963 29296 4972 29336
rect 5012 29296 5021 29336
rect 4963 29295 5021 29296
rect 11979 29336 12021 29345
rect 11979 29296 11980 29336
rect 12020 29296 12021 29336
rect 11979 29287 12021 29296
rect 14187 29336 14229 29345
rect 14187 29296 14188 29336
rect 14228 29296 14229 29336
rect 14187 29287 14229 29296
rect 15619 29336 15677 29337
rect 15619 29296 15628 29336
rect 15668 29296 15677 29336
rect 15619 29295 15677 29296
rect 19851 29336 19893 29345
rect 19851 29296 19852 29336
rect 19892 29296 19893 29336
rect 19851 29287 19893 29296
rect 6891 29252 6933 29261
rect 6891 29212 6892 29252
rect 6932 29212 6933 29252
rect 6891 29203 6933 29212
rect 8907 29252 8949 29261
rect 8907 29212 8908 29252
rect 8948 29212 8949 29252
rect 8907 29203 8949 29212
rect 14859 29252 14901 29261
rect 14859 29212 14860 29252
rect 14900 29212 14901 29252
rect 14859 29203 14901 29212
rect 18219 29252 18261 29261
rect 18219 29212 18220 29252
rect 18260 29212 18261 29252
rect 18219 29203 18261 29212
rect 2187 29168 2229 29177
rect 2187 29128 2188 29168
rect 2228 29128 2229 29168
rect 2467 29168 2525 29169
rect 2187 29119 2229 29128
rect 2319 29158 2361 29167
rect 2319 29118 2320 29158
rect 2360 29118 2361 29158
rect 2467 29128 2476 29168
rect 2516 29128 2525 29168
rect 2467 29127 2525 29128
rect 3715 29168 3773 29169
rect 3715 29128 3724 29168
rect 3764 29128 3773 29168
rect 3715 29127 3773 29128
rect 4491 29168 4533 29177
rect 4491 29128 4492 29168
rect 4532 29128 4533 29168
rect 4491 29119 4533 29128
rect 4587 29168 4629 29177
rect 4587 29128 4588 29168
rect 4628 29128 4629 29168
rect 4587 29119 4629 29128
rect 5163 29168 5205 29177
rect 5163 29128 5164 29168
rect 5204 29128 5205 29168
rect 5163 29119 5205 29128
rect 5259 29168 5301 29177
rect 5259 29128 5260 29168
rect 5300 29128 5301 29168
rect 5259 29119 5301 29128
rect 5443 29168 5501 29169
rect 5443 29128 5452 29168
rect 5492 29128 5501 29168
rect 5443 29127 5501 29128
rect 6691 29168 6749 29169
rect 6691 29128 6700 29168
rect 6740 29128 6749 29168
rect 6691 29127 6749 29128
rect 7179 29168 7221 29177
rect 7179 29128 7180 29168
rect 7220 29128 7221 29168
rect 7179 29119 7221 29128
rect 7275 29168 7317 29177
rect 7275 29128 7276 29168
rect 7316 29128 7317 29168
rect 7275 29119 7317 29128
rect 7659 29168 7701 29177
rect 7659 29128 7660 29168
rect 7700 29128 7701 29168
rect 7659 29119 7701 29128
rect 7755 29168 7797 29177
rect 7755 29128 7756 29168
rect 7796 29128 7797 29168
rect 7755 29119 7797 29128
rect 8227 29168 8285 29169
rect 8227 29128 8236 29168
rect 8276 29128 8285 29168
rect 8227 29127 8285 29128
rect 8715 29163 8757 29172
rect 8715 29123 8716 29163
rect 8756 29123 8757 29163
rect 2319 29109 2361 29118
rect 8715 29114 8757 29123
rect 10251 29168 10293 29177
rect 10251 29128 10252 29168
rect 10292 29128 10293 29168
rect 10251 29119 10293 29128
rect 10347 29168 10389 29177
rect 10347 29128 10348 29168
rect 10388 29128 10389 29168
rect 10347 29119 10389 29128
rect 10731 29168 10773 29177
rect 10731 29128 10732 29168
rect 10772 29128 10773 29168
rect 10731 29119 10773 29128
rect 10827 29168 10869 29177
rect 10827 29128 10828 29168
rect 10868 29128 10869 29168
rect 10827 29119 10869 29128
rect 11299 29168 11357 29169
rect 11299 29128 11308 29168
rect 11348 29128 11357 29168
rect 12739 29168 12797 29169
rect 11299 29127 11357 29128
rect 11787 29154 11829 29163
rect 11787 29114 11788 29154
rect 11828 29114 11829 29154
rect 12739 29128 12748 29168
rect 12788 29128 12797 29168
rect 12739 29127 12797 29128
rect 13987 29168 14045 29169
rect 13987 29128 13996 29168
rect 14036 29128 14045 29168
rect 13987 29127 14045 29128
rect 14467 29168 14525 29169
rect 14467 29128 14476 29168
rect 14516 29128 14525 29168
rect 14467 29127 14525 29128
rect 14763 29168 14805 29177
rect 14763 29128 14764 29168
rect 14804 29128 14805 29168
rect 14763 29119 14805 29128
rect 16491 29168 16533 29177
rect 16491 29128 16492 29168
rect 16532 29128 16533 29168
rect 16491 29119 16533 29128
rect 16587 29168 16629 29177
rect 16587 29128 16588 29168
rect 16628 29128 16629 29168
rect 16587 29119 16629 29128
rect 17539 29168 17597 29169
rect 17539 29128 17548 29168
rect 17588 29128 17597 29168
rect 18403 29168 18461 29169
rect 17539 29127 17597 29128
rect 18027 29154 18069 29163
rect 11787 29105 11829 29114
rect 18027 29114 18028 29154
rect 18068 29114 18069 29154
rect 18403 29128 18412 29168
rect 18452 29128 18461 29168
rect 18403 29127 18461 29128
rect 18027 29105 18069 29114
rect 19651 29126 19709 29127
rect 16971 29084 17013 29093
rect 16971 29044 16972 29084
rect 17012 29044 17013 29084
rect 16971 29035 17013 29044
rect 17067 29084 17109 29093
rect 19651 29086 19660 29126
rect 19700 29086 19709 29126
rect 19651 29085 19709 29086
rect 17067 29044 17068 29084
rect 17108 29044 17109 29084
rect 17067 29035 17109 29044
rect 20035 29084 20093 29085
rect 20035 29044 20044 29084
rect 20084 29044 20093 29084
rect 20035 29043 20093 29044
rect 3915 29000 3957 29009
rect 3915 28960 3916 29000
rect 3956 28960 3957 29000
rect 3915 28951 3957 28960
rect 15723 29000 15765 29009
rect 15723 28960 15724 29000
rect 15764 28960 15765 29000
rect 15723 28951 15765 28960
rect 20235 28916 20277 28925
rect 20235 28876 20236 28916
rect 20276 28876 20277 28916
rect 15139 28874 15197 28875
rect 15139 28834 15148 28874
rect 15188 28834 15197 28874
rect 20235 28867 20277 28876
rect 15139 28833 15197 28834
rect 1152 28748 20352 28772
rect 1152 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 20352 28748
rect 1152 28684 20352 28708
rect 11691 28580 11733 28589
rect 11691 28540 11692 28580
rect 11732 28540 11733 28580
rect 11691 28531 11733 28540
rect 12171 28580 12213 28589
rect 12171 28540 12172 28580
rect 12212 28540 12213 28580
rect 12171 28531 12213 28540
rect 15435 28580 15477 28589
rect 15435 28540 15436 28580
rect 15476 28540 15477 28580
rect 15435 28531 15477 28540
rect 15915 28580 15957 28589
rect 15915 28540 15916 28580
rect 15956 28540 15957 28580
rect 15915 28531 15957 28540
rect 18987 28580 19029 28589
rect 18987 28540 18988 28580
rect 19028 28540 19029 28580
rect 18987 28531 19029 28540
rect 19755 28580 19797 28589
rect 19755 28540 19756 28580
rect 19796 28540 19797 28580
rect 19755 28531 19797 28540
rect 20139 28580 20181 28589
rect 20139 28540 20140 28580
rect 20180 28540 20181 28580
rect 20139 28531 20181 28540
rect 1803 28496 1845 28505
rect 1803 28456 1804 28496
rect 1844 28456 1845 28496
rect 1803 28447 1845 28456
rect 15627 28496 15669 28505
rect 15627 28456 15628 28496
rect 15668 28456 15669 28496
rect 15627 28447 15669 28456
rect 3531 28412 3573 28421
rect 3531 28372 3532 28412
rect 3572 28372 3573 28412
rect 3531 28363 3573 28372
rect 19171 28412 19229 28413
rect 19171 28372 19180 28412
rect 19220 28372 19229 28412
rect 19171 28371 19229 28372
rect 19555 28412 19613 28413
rect 19555 28372 19564 28412
rect 19604 28372 19613 28412
rect 19555 28371 19613 28372
rect 19939 28412 19997 28413
rect 19939 28372 19948 28412
rect 19988 28372 19997 28412
rect 19939 28371 19997 28372
rect 3051 28328 3093 28337
rect 3051 28288 3052 28328
rect 3092 28288 3093 28328
rect 3051 28279 3093 28288
rect 3147 28328 3189 28337
rect 3147 28288 3148 28328
rect 3188 28288 3189 28328
rect 3147 28279 3189 28288
rect 3627 28328 3669 28337
rect 4587 28333 4629 28342
rect 3627 28288 3628 28328
rect 3668 28288 3669 28328
rect 3627 28279 3669 28288
rect 4099 28328 4157 28329
rect 4099 28288 4108 28328
rect 4148 28288 4157 28328
rect 4099 28287 4157 28288
rect 4587 28293 4588 28333
rect 4628 28293 4629 28333
rect 4587 28284 4629 28293
rect 5059 28328 5117 28329
rect 5059 28288 5068 28328
rect 5108 28288 5117 28328
rect 5059 28287 5117 28288
rect 6307 28328 6365 28329
rect 6307 28288 6316 28328
rect 6356 28288 6365 28328
rect 6307 28287 6365 28288
rect 6795 28328 6837 28337
rect 6795 28288 6796 28328
rect 6836 28288 6837 28328
rect 6795 28279 6837 28288
rect 6891 28328 6933 28337
rect 6891 28288 6892 28328
rect 6932 28288 6933 28328
rect 6891 28279 6933 28288
rect 7275 28328 7317 28337
rect 7275 28288 7276 28328
rect 7316 28288 7317 28328
rect 7275 28279 7317 28288
rect 7371 28328 7413 28337
rect 8331 28333 8373 28342
rect 7371 28288 7372 28328
rect 7412 28288 7413 28328
rect 7371 28279 7413 28288
rect 7843 28328 7901 28329
rect 7843 28288 7852 28328
rect 7892 28288 7901 28328
rect 7843 28287 7901 28288
rect 8331 28293 8332 28333
rect 8372 28293 8373 28333
rect 8331 28284 8373 28293
rect 10243 28328 10301 28329
rect 10243 28288 10252 28328
rect 10292 28288 10301 28328
rect 10243 28287 10301 28288
rect 11491 28328 11549 28329
rect 11491 28288 11500 28328
rect 11540 28288 11549 28328
rect 11491 28287 11549 28288
rect 11883 28328 11925 28337
rect 11883 28288 11884 28328
rect 11924 28288 11925 28328
rect 11883 28279 11925 28288
rect 12171 28328 12213 28337
rect 12171 28288 12172 28328
rect 12212 28288 12213 28328
rect 12171 28279 12213 28288
rect 12547 28328 12605 28329
rect 12547 28288 12556 28328
rect 12596 28288 12605 28328
rect 12547 28287 12605 28288
rect 13795 28328 13853 28329
rect 13795 28288 13804 28328
rect 13844 28288 13853 28328
rect 13795 28287 13853 28288
rect 13987 28328 14045 28329
rect 13987 28288 13996 28328
rect 14036 28288 14045 28328
rect 13987 28287 14045 28288
rect 15235 28328 15293 28329
rect 15235 28288 15244 28328
rect 15284 28288 15293 28328
rect 15235 28287 15293 28288
rect 16099 28328 16157 28329
rect 16099 28288 16108 28328
rect 16148 28288 16157 28328
rect 16099 28287 16157 28288
rect 17347 28328 17405 28329
rect 17347 28288 17356 28328
rect 17396 28288 17405 28328
rect 17347 28287 17405 28288
rect 17539 28328 17597 28329
rect 17539 28288 17548 28328
rect 17588 28288 17597 28328
rect 17539 28287 17597 28288
rect 18787 28328 18845 28329
rect 18787 28288 18796 28328
rect 18836 28288 18845 28328
rect 18787 28287 18845 28288
rect 4779 28244 4821 28253
rect 4779 28204 4780 28244
rect 4820 28204 4821 28244
rect 4779 28195 4821 28204
rect 6507 28244 6549 28253
rect 6507 28204 6508 28244
rect 6548 28204 6549 28244
rect 6507 28195 6549 28204
rect 1699 28160 1757 28161
rect 1699 28120 1708 28160
rect 1748 28120 1757 28160
rect 1699 28119 1757 28120
rect 8523 28160 8565 28169
rect 8523 28120 8524 28160
rect 8564 28120 8565 28160
rect 8523 28111 8565 28120
rect 12363 28160 12405 28169
rect 12363 28120 12364 28160
rect 12404 28120 12405 28160
rect 12363 28111 12405 28120
rect 19371 28160 19413 28169
rect 19371 28120 19372 28160
rect 19412 28120 19413 28160
rect 19371 28111 19413 28120
rect 1152 27992 20452 28016
rect 1152 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20452 27992
rect 1152 27928 20452 27952
rect 3147 27824 3189 27833
rect 3147 27784 3148 27824
rect 3188 27784 3189 27824
rect 3147 27775 3189 27784
rect 8235 27824 8277 27833
rect 8235 27784 8236 27824
rect 8276 27784 8277 27824
rect 8235 27775 8277 27784
rect 15435 27824 15477 27833
rect 15435 27784 15436 27824
rect 15476 27784 15477 27824
rect 15435 27775 15477 27784
rect 16579 27824 16637 27825
rect 16579 27784 16588 27824
rect 16628 27784 16637 27824
rect 16579 27783 16637 27784
rect 20043 27824 20085 27833
rect 20043 27784 20044 27824
rect 20084 27784 20085 27824
rect 20043 27775 20085 27784
rect 6507 27740 6549 27749
rect 6507 27700 6508 27740
rect 6548 27700 6549 27740
rect 6507 27691 6549 27700
rect 9867 27740 9909 27749
rect 9867 27700 9868 27740
rect 9908 27700 9909 27740
rect 9867 27691 9909 27700
rect 11883 27740 11925 27749
rect 11883 27700 11884 27740
rect 11924 27700 11925 27740
rect 11883 27691 11925 27700
rect 16011 27740 16053 27749
rect 16011 27700 16012 27740
rect 16052 27700 16053 27740
rect 16011 27691 16053 27700
rect 17451 27740 17493 27749
rect 17451 27700 17452 27740
rect 17492 27700 17493 27740
rect 17451 27691 17493 27700
rect 1699 27656 1757 27657
rect 1699 27616 1708 27656
rect 1748 27616 1757 27656
rect 1699 27615 1757 27616
rect 2947 27656 3005 27657
rect 2947 27616 2956 27656
rect 2996 27616 3005 27656
rect 2947 27615 3005 27616
rect 3339 27656 3381 27665
rect 3339 27616 3340 27656
rect 3380 27616 3381 27656
rect 3339 27607 3381 27616
rect 3531 27656 3573 27665
rect 3531 27616 3532 27656
rect 3572 27616 3573 27656
rect 3531 27607 3573 27616
rect 3715 27656 3773 27657
rect 3715 27616 3724 27656
rect 3764 27616 3773 27656
rect 3715 27615 3773 27616
rect 4963 27656 5021 27657
rect 4963 27616 4972 27656
rect 5012 27616 5021 27656
rect 4963 27615 5021 27616
rect 5443 27656 5501 27657
rect 5443 27616 5452 27656
rect 5492 27616 5501 27656
rect 5443 27615 5501 27616
rect 5739 27656 5781 27665
rect 5739 27616 5740 27656
rect 5780 27616 5781 27656
rect 5739 27607 5781 27616
rect 5835 27656 5877 27665
rect 5835 27616 5836 27656
rect 5876 27616 5877 27656
rect 5835 27607 5877 27616
rect 6307 27656 6365 27657
rect 6307 27616 6316 27656
rect 6356 27616 6365 27656
rect 6307 27615 6365 27616
rect 6411 27656 6453 27665
rect 6411 27616 6412 27656
rect 6452 27616 6453 27656
rect 6411 27607 6453 27616
rect 6603 27656 6645 27665
rect 6603 27616 6604 27656
rect 6644 27616 6645 27656
rect 6603 27607 6645 27616
rect 6787 27656 6845 27657
rect 6787 27616 6796 27656
rect 6836 27616 6845 27656
rect 6787 27615 6845 27616
rect 8035 27656 8093 27657
rect 8035 27616 8044 27656
rect 8084 27616 8093 27656
rect 8035 27615 8093 27616
rect 8419 27656 8477 27657
rect 8419 27616 8428 27656
rect 8468 27616 8477 27656
rect 8419 27615 8477 27616
rect 9667 27656 9725 27657
rect 9667 27616 9676 27656
rect 9716 27616 9725 27656
rect 9667 27615 9725 27616
rect 10155 27656 10197 27665
rect 10155 27616 10156 27656
rect 10196 27616 10197 27656
rect 10155 27607 10197 27616
rect 10251 27656 10293 27665
rect 10251 27616 10252 27656
rect 10292 27616 10293 27656
rect 10251 27607 10293 27616
rect 10731 27656 10773 27665
rect 10731 27616 10732 27656
rect 10772 27616 10773 27656
rect 10731 27607 10773 27616
rect 11203 27656 11261 27657
rect 11203 27616 11212 27656
rect 11252 27616 11261 27656
rect 12067 27656 12125 27657
rect 11203 27615 11261 27616
rect 11691 27642 11733 27651
rect 11691 27602 11692 27642
rect 11732 27602 11733 27642
rect 12067 27616 12076 27656
rect 12116 27616 12125 27656
rect 12067 27615 12125 27616
rect 13315 27656 13373 27657
rect 13315 27616 13324 27656
rect 13364 27616 13373 27656
rect 13315 27615 13373 27616
rect 13987 27656 14045 27657
rect 13987 27616 13996 27656
rect 14036 27616 14045 27656
rect 13987 27615 14045 27616
rect 15235 27656 15293 27657
rect 15235 27616 15244 27656
rect 15284 27616 15293 27656
rect 15235 27615 15293 27616
rect 15915 27656 15957 27665
rect 15915 27616 15916 27656
rect 15956 27616 15957 27656
rect 15915 27607 15957 27616
rect 16107 27656 16149 27665
rect 16107 27616 16108 27656
rect 16148 27616 16149 27656
rect 16683 27656 16725 27665
rect 16107 27607 16149 27616
rect 16491 27645 16533 27654
rect 11691 27593 11733 27602
rect 16491 27605 16492 27645
rect 16532 27605 16533 27645
rect 16683 27616 16684 27656
rect 16724 27616 16725 27656
rect 16683 27607 16725 27616
rect 16771 27656 16829 27657
rect 16771 27616 16780 27656
rect 16820 27616 16829 27656
rect 18115 27656 18173 27657
rect 16771 27615 16829 27616
rect 17643 27642 17685 27651
rect 16491 27596 16533 27605
rect 17643 27602 17644 27642
rect 17684 27602 17685 27642
rect 18115 27616 18124 27656
rect 18164 27616 18173 27656
rect 18115 27615 18173 27616
rect 18603 27656 18645 27665
rect 18603 27616 18604 27656
rect 18644 27616 18645 27656
rect 18603 27607 18645 27616
rect 18699 27656 18741 27665
rect 18699 27616 18700 27656
rect 18740 27616 18741 27656
rect 18699 27607 18741 27616
rect 19083 27656 19125 27665
rect 19083 27616 19084 27656
rect 19124 27616 19125 27656
rect 19083 27607 19125 27616
rect 19179 27656 19221 27665
rect 19179 27616 19180 27656
rect 19220 27616 19221 27656
rect 19179 27607 19221 27616
rect 17643 27593 17685 27602
rect 10635 27572 10677 27581
rect 10635 27532 10636 27572
rect 10676 27532 10677 27572
rect 10635 27523 10677 27532
rect 17059 27572 17117 27573
rect 17059 27532 17068 27572
rect 17108 27532 17117 27572
rect 17059 27531 17117 27532
rect 19459 27572 19517 27573
rect 19459 27532 19468 27572
rect 19508 27532 19517 27572
rect 19459 27531 19517 27532
rect 19843 27572 19901 27573
rect 19843 27532 19852 27572
rect 19892 27532 19901 27572
rect 19843 27531 19901 27532
rect 5163 27488 5205 27497
rect 5163 27448 5164 27488
rect 5204 27448 5205 27488
rect 5163 27439 5205 27448
rect 15723 27488 15765 27497
rect 15723 27448 15724 27488
rect 15764 27448 15765 27488
rect 15723 27439 15765 27448
rect 19659 27488 19701 27497
rect 19659 27448 19660 27488
rect 19700 27448 19701 27488
rect 19659 27439 19701 27448
rect 3531 27404 3573 27413
rect 3531 27364 3532 27404
rect 3572 27364 3573 27404
rect 3531 27355 3573 27364
rect 6115 27404 6173 27405
rect 6115 27364 6124 27404
rect 6164 27364 6173 27404
rect 6115 27363 6173 27364
rect 13515 27404 13557 27413
rect 13515 27364 13516 27404
rect 13556 27364 13557 27404
rect 13515 27355 13557 27364
rect 17259 27404 17301 27413
rect 17259 27364 17260 27404
rect 17300 27364 17301 27404
rect 17259 27355 17301 27364
rect 1152 27236 20352 27260
rect 1152 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 20352 27236
rect 1152 27172 20352 27196
rect 3435 27068 3477 27077
rect 3435 27028 3436 27068
rect 3476 27028 3477 27068
rect 3435 27019 3477 27028
rect 5067 27068 5109 27077
rect 5067 27028 5068 27068
rect 5108 27028 5109 27068
rect 5067 27019 5109 27028
rect 5643 27068 5685 27077
rect 5643 27028 5644 27068
rect 5684 27028 5685 27068
rect 5643 27019 5685 27028
rect 11499 27068 11541 27077
rect 11499 27028 11500 27068
rect 11540 27028 11541 27068
rect 11499 27019 11541 27028
rect 15435 27068 15477 27077
rect 15435 27028 15436 27068
rect 15476 27028 15477 27068
rect 15435 27019 15477 27028
rect 1707 26984 1749 26993
rect 1707 26944 1708 26984
rect 1748 26944 1749 26984
rect 1707 26935 1749 26944
rect 16963 26984 17021 26985
rect 16963 26944 16972 26984
rect 17012 26944 17021 26984
rect 16963 26943 17021 26944
rect 8235 26900 8277 26909
rect 8235 26860 8236 26900
rect 8276 26860 8277 26900
rect 8235 26851 8277 26860
rect 15235 26900 15293 26901
rect 15235 26860 15244 26900
rect 15284 26860 15293 26900
rect 15235 26859 15293 26860
rect 19363 26900 19421 26901
rect 19363 26860 19372 26900
rect 19412 26860 19421 26900
rect 19363 26859 19421 26860
rect 19747 26900 19805 26901
rect 19747 26860 19756 26900
rect 19796 26860 19805 26900
rect 19747 26859 19805 26860
rect 14379 26830 14421 26839
rect 1227 26816 1269 26825
rect 1227 26776 1228 26816
rect 1268 26776 1269 26816
rect 1227 26767 1269 26776
rect 1323 26816 1365 26825
rect 1323 26776 1324 26816
rect 1364 26776 1365 26816
rect 1323 26767 1365 26776
rect 1419 26816 1461 26825
rect 1419 26776 1420 26816
rect 1460 26776 1461 26816
rect 1419 26767 1461 26776
rect 1515 26816 1557 26825
rect 1515 26776 1516 26816
rect 1556 26776 1557 26816
rect 1515 26767 1557 26776
rect 1987 26816 2045 26817
rect 1987 26776 1996 26816
rect 2036 26776 2045 26816
rect 1987 26775 2045 26776
rect 3235 26816 3293 26817
rect 3235 26776 3244 26816
rect 3284 26776 3293 26816
rect 3235 26775 3293 26776
rect 3619 26816 3677 26817
rect 3619 26776 3628 26816
rect 3668 26776 3677 26816
rect 3619 26775 3677 26776
rect 4867 26816 4925 26817
rect 4867 26776 4876 26816
rect 4916 26776 4925 26816
rect 4867 26775 4925 26776
rect 5355 26816 5397 26825
rect 5355 26776 5356 26816
rect 5396 26776 5397 26816
rect 5355 26767 5397 26776
rect 5643 26816 5685 26825
rect 5643 26776 5644 26816
rect 5684 26776 5685 26816
rect 5643 26767 5685 26776
rect 6019 26816 6077 26817
rect 6019 26776 6028 26816
rect 6068 26776 6077 26816
rect 6019 26775 6077 26776
rect 7267 26816 7325 26817
rect 7267 26776 7276 26816
rect 7316 26776 7325 26816
rect 7267 26775 7325 26776
rect 7755 26816 7797 26825
rect 7755 26776 7756 26816
rect 7796 26776 7797 26816
rect 7755 26767 7797 26776
rect 7851 26816 7893 26825
rect 7851 26776 7852 26816
rect 7892 26776 7893 26816
rect 7851 26767 7893 26776
rect 8331 26816 8373 26825
rect 9291 26821 9333 26830
rect 8331 26776 8332 26816
rect 8372 26776 8373 26816
rect 8331 26767 8373 26776
rect 8803 26816 8861 26817
rect 8803 26776 8812 26816
rect 8852 26776 8861 26816
rect 8803 26775 8861 26776
rect 9291 26781 9292 26821
rect 9332 26781 9333 26821
rect 9291 26772 9333 26781
rect 10051 26816 10109 26817
rect 10051 26776 10060 26816
rect 10100 26776 10109 26816
rect 10051 26775 10109 26776
rect 11299 26816 11357 26817
rect 11299 26776 11308 26816
rect 11348 26776 11357 26816
rect 11299 26775 11357 26776
rect 12843 26816 12885 26825
rect 12843 26776 12844 26816
rect 12884 26776 12885 26816
rect 12843 26767 12885 26776
rect 12939 26816 12981 26825
rect 12939 26776 12940 26816
rect 12980 26776 12981 26816
rect 12939 26767 12981 26776
rect 13323 26816 13365 26825
rect 13323 26776 13324 26816
rect 13364 26776 13365 26816
rect 13323 26767 13365 26776
rect 13419 26816 13461 26825
rect 13419 26776 13420 26816
rect 13460 26776 13461 26816
rect 13419 26767 13461 26776
rect 13891 26816 13949 26817
rect 13891 26776 13900 26816
rect 13940 26776 13949 26816
rect 14379 26790 14380 26830
rect 14420 26790 14421 26830
rect 14379 26781 14421 26790
rect 14763 26816 14805 26825
rect 13891 26775 13949 26776
rect 14763 26776 14764 26816
rect 14804 26776 14805 26816
rect 14763 26767 14805 26776
rect 14859 26816 14901 26825
rect 14859 26776 14860 26816
rect 14900 26776 14901 26816
rect 14859 26767 14901 26776
rect 16291 26816 16349 26817
rect 16291 26776 16300 26816
rect 16340 26776 16349 26816
rect 16291 26775 16349 26776
rect 16587 26816 16629 26825
rect 16587 26776 16588 26816
rect 16628 26776 16629 26816
rect 16587 26767 16629 26776
rect 16683 26816 16725 26825
rect 16683 26776 16684 26816
rect 16724 26776 16725 26816
rect 16683 26767 16725 26776
rect 17259 26816 17301 26825
rect 17259 26776 17260 26816
rect 17300 26776 17301 26816
rect 17259 26767 17301 26776
rect 17355 26816 17397 26825
rect 17355 26776 17356 26816
rect 17396 26776 17397 26816
rect 17355 26767 17397 26776
rect 17739 26816 17781 26825
rect 17739 26776 17740 26816
rect 17780 26776 17781 26816
rect 17739 26767 17781 26776
rect 17835 26816 17877 26825
rect 18795 26821 18837 26830
rect 17835 26776 17836 26816
rect 17876 26776 17877 26816
rect 17835 26767 17877 26776
rect 18307 26816 18365 26817
rect 18307 26776 18316 26816
rect 18356 26776 18365 26816
rect 18307 26775 18365 26776
rect 18795 26781 18796 26821
rect 18836 26781 18837 26821
rect 18795 26772 18837 26781
rect 7467 26732 7509 26741
rect 7467 26692 7468 26732
rect 7508 26692 7509 26732
rect 7467 26683 7509 26692
rect 14571 26732 14613 26741
rect 14571 26692 14572 26732
rect 14612 26692 14613 26732
rect 14571 26683 14613 26692
rect 1699 26648 1757 26649
rect 1699 26608 1708 26648
rect 1748 26608 1757 26648
rect 1699 26607 1757 26608
rect 5067 26648 5109 26657
rect 5067 26608 5068 26648
rect 5108 26608 5109 26648
rect 5067 26599 5109 26608
rect 9483 26648 9525 26657
rect 9483 26608 9484 26648
rect 9524 26608 9525 26648
rect 9483 26599 9525 26608
rect 15043 26648 15101 26649
rect 15043 26608 15052 26648
rect 15092 26608 15101 26648
rect 15043 26607 15101 26608
rect 15619 26648 15677 26649
rect 15619 26608 15628 26648
rect 15668 26608 15677 26648
rect 15619 26607 15677 26608
rect 15907 26648 15965 26649
rect 15907 26608 15916 26648
rect 15956 26608 15965 26648
rect 15907 26607 15965 26608
rect 18987 26648 19029 26657
rect 18987 26608 18988 26648
rect 19028 26608 19029 26648
rect 18987 26599 19029 26608
rect 19563 26648 19605 26657
rect 19563 26608 19564 26648
rect 19604 26608 19605 26648
rect 19563 26599 19605 26608
rect 19947 26648 19989 26657
rect 19947 26608 19948 26648
rect 19988 26608 19989 26648
rect 19947 26599 19989 26608
rect 1152 26480 20452 26504
rect 1152 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20452 26480
rect 1152 26416 20452 26440
rect 1699 26312 1757 26313
rect 1699 26272 1708 26312
rect 1748 26272 1757 26312
rect 1699 26271 1757 26272
rect 3435 26312 3477 26321
rect 3435 26272 3436 26312
rect 3476 26272 3477 26312
rect 3435 26263 3477 26272
rect 3627 26312 3669 26321
rect 3627 26272 3628 26312
rect 3668 26272 3669 26312
rect 3627 26263 3669 26272
rect 8523 26312 8565 26321
rect 8523 26272 8524 26312
rect 8564 26272 8565 26312
rect 8523 26263 8565 26272
rect 10155 26312 10197 26321
rect 10155 26272 10156 26312
rect 10196 26272 10197 26312
rect 10155 26263 10197 26272
rect 17067 26312 17109 26321
rect 17067 26272 17068 26312
rect 17108 26272 17109 26312
rect 17067 26263 17109 26272
rect 18699 26312 18741 26321
rect 18699 26272 18700 26312
rect 18740 26272 18741 26312
rect 18699 26263 18741 26272
rect 19171 26312 19229 26313
rect 19171 26272 19180 26312
rect 19220 26272 19229 26312
rect 19171 26271 19229 26272
rect 1227 26228 1269 26237
rect 1227 26188 1228 26228
rect 1268 26188 1269 26228
rect 1227 26179 1269 26188
rect 1323 26144 1365 26153
rect 1323 26104 1324 26144
rect 1364 26104 1365 26144
rect 1323 26095 1365 26104
rect 1419 26144 1461 26153
rect 1419 26104 1420 26144
rect 1460 26104 1461 26144
rect 1419 26095 1461 26104
rect 1515 26144 1557 26153
rect 1515 26104 1516 26144
rect 1556 26104 1557 26144
rect 1515 26095 1557 26104
rect 1987 26144 2045 26145
rect 1987 26104 1996 26144
rect 2036 26104 2045 26144
rect 1987 26103 2045 26104
rect 3235 26144 3293 26145
rect 3235 26104 3244 26144
rect 3284 26104 3293 26144
rect 3235 26103 3293 26104
rect 3811 26144 3869 26145
rect 3811 26104 3820 26144
rect 3860 26104 3869 26144
rect 3811 26103 3869 26104
rect 5059 26144 5117 26145
rect 5059 26104 5068 26144
rect 5108 26104 5117 26144
rect 5059 26103 5117 26104
rect 5443 26144 5501 26145
rect 5443 26104 5452 26144
rect 5492 26104 5501 26144
rect 5443 26103 5501 26104
rect 6691 26144 6749 26145
rect 6691 26104 6700 26144
rect 6740 26104 6749 26144
rect 6691 26103 6749 26104
rect 7075 26144 7133 26145
rect 7075 26104 7084 26144
rect 7124 26104 7133 26144
rect 7075 26103 7133 26104
rect 8323 26144 8381 26145
rect 8323 26104 8332 26144
rect 8372 26104 8381 26144
rect 8323 26103 8381 26104
rect 8707 26144 8765 26145
rect 8707 26104 8716 26144
rect 8756 26104 8765 26144
rect 8707 26103 8765 26104
rect 9955 26144 10013 26145
rect 9955 26104 9964 26144
rect 10004 26104 10013 26144
rect 9955 26103 10013 26104
rect 12747 26144 12789 26153
rect 12747 26104 12748 26144
rect 12788 26104 12789 26144
rect 12747 26095 12789 26104
rect 12843 26144 12885 26153
rect 12843 26104 12844 26144
rect 12884 26104 12885 26144
rect 12843 26095 12885 26104
rect 13123 26144 13181 26145
rect 13123 26104 13132 26144
rect 13172 26104 13181 26144
rect 13123 26103 13181 26104
rect 13419 26144 13461 26153
rect 13419 26104 13420 26144
rect 13460 26104 13461 26144
rect 13419 26095 13461 26104
rect 13611 26144 13653 26153
rect 13611 26104 13612 26144
rect 13652 26104 13653 26144
rect 13611 26095 13653 26104
rect 13795 26144 13853 26145
rect 13795 26104 13804 26144
rect 13844 26104 13853 26144
rect 13795 26103 13853 26104
rect 15043 26144 15101 26145
rect 15043 26104 15052 26144
rect 15092 26104 15101 26144
rect 15043 26103 15101 26104
rect 15619 26144 15677 26145
rect 15619 26104 15628 26144
rect 15668 26104 15677 26144
rect 15619 26103 15677 26104
rect 16867 26144 16925 26145
rect 16867 26104 16876 26144
rect 16916 26104 16925 26144
rect 16867 26103 16925 26104
rect 17251 26144 17309 26145
rect 17251 26104 17260 26144
rect 17300 26104 17309 26144
rect 17251 26103 17309 26104
rect 18499 26144 18557 26145
rect 18499 26104 18508 26144
rect 18548 26104 18557 26144
rect 18499 26103 18557 26104
rect 18891 26144 18933 26153
rect 18891 26104 18892 26144
rect 18932 26104 18933 26144
rect 18891 26095 18933 26104
rect 18987 26144 19029 26153
rect 18987 26104 18988 26144
rect 19028 26104 19029 26144
rect 18987 26095 19029 26104
rect 19755 26144 19797 26153
rect 19755 26104 19756 26144
rect 19796 26104 19797 26144
rect 19755 26095 19797 26104
rect 19851 26144 19893 26153
rect 19851 26104 19852 26144
rect 19892 26104 19893 26144
rect 19851 26095 19893 26104
rect 19947 26144 19989 26153
rect 19947 26104 19948 26144
rect 19988 26104 19989 26144
rect 19947 26095 19989 26104
rect 20043 26144 20085 26153
rect 20043 26104 20044 26144
rect 20084 26104 20085 26144
rect 20043 26095 20085 26104
rect 19363 26060 19421 26061
rect 19363 26020 19372 26060
rect 19412 26020 19421 26060
rect 19363 26019 19421 26020
rect 6891 25892 6933 25901
rect 6891 25852 6892 25892
rect 6932 25852 6933 25892
rect 6891 25843 6933 25852
rect 12451 25892 12509 25893
rect 12451 25852 12460 25892
rect 12500 25852 12509 25892
rect 12451 25851 12509 25852
rect 13611 25892 13653 25901
rect 13611 25852 13612 25892
rect 13652 25852 13653 25892
rect 13611 25843 13653 25852
rect 15243 25892 15285 25901
rect 15243 25852 15244 25892
rect 15284 25852 15285 25892
rect 15243 25843 15285 25852
rect 19563 25892 19605 25901
rect 19563 25852 19564 25892
rect 19604 25852 19605 25892
rect 19563 25843 19605 25852
rect 1152 25724 20352 25748
rect 1152 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 20352 25724
rect 1152 25660 20352 25684
rect 1995 25556 2037 25565
rect 1995 25516 1996 25556
rect 2036 25516 2037 25556
rect 1995 25507 2037 25516
rect 11595 25556 11637 25565
rect 11595 25516 11596 25556
rect 11636 25516 11637 25556
rect 11595 25507 11637 25516
rect 17451 25556 17493 25565
rect 17451 25516 17452 25556
rect 17492 25516 17493 25556
rect 17451 25507 17493 25516
rect 19083 25556 19125 25565
rect 19083 25516 19084 25556
rect 19124 25516 19125 25556
rect 19083 25507 19125 25516
rect 1707 25472 1749 25481
rect 1707 25432 1708 25472
rect 1748 25432 1749 25472
rect 1707 25423 1749 25432
rect 13035 25388 13077 25397
rect 13035 25348 13036 25388
rect 13076 25348 13077 25388
rect 13035 25339 13077 25348
rect 4011 25318 4053 25327
rect 1227 25304 1269 25313
rect 1227 25264 1228 25304
rect 1268 25264 1269 25304
rect 1227 25255 1269 25264
rect 1419 25304 1461 25313
rect 1419 25264 1420 25304
rect 1460 25264 1461 25304
rect 1419 25255 1461 25264
rect 1515 25304 1557 25313
rect 1515 25264 1516 25304
rect 1556 25264 1557 25304
rect 1515 25255 1557 25264
rect 2179 25304 2237 25305
rect 2179 25264 2188 25304
rect 2228 25264 2237 25304
rect 2179 25263 2237 25264
rect 3427 25304 3485 25305
rect 3427 25264 3436 25304
rect 3476 25264 3485 25304
rect 4011 25278 4012 25318
rect 4052 25278 4053 25318
rect 4011 25269 4053 25278
rect 4483 25304 4541 25305
rect 3427 25263 3485 25264
rect 4483 25264 4492 25304
rect 4532 25264 4541 25304
rect 4483 25263 4541 25264
rect 4971 25304 5013 25313
rect 4971 25264 4972 25304
rect 5012 25264 5013 25304
rect 4971 25255 5013 25264
rect 5067 25304 5109 25313
rect 5067 25264 5068 25304
rect 5108 25264 5109 25304
rect 5067 25255 5109 25264
rect 5451 25304 5493 25313
rect 5451 25264 5452 25304
rect 5492 25264 5493 25304
rect 5451 25255 5493 25264
rect 5547 25304 5589 25313
rect 5547 25264 5548 25304
rect 5588 25264 5589 25304
rect 5547 25255 5589 25264
rect 5835 25304 5877 25313
rect 5835 25264 5836 25304
rect 5876 25264 5877 25304
rect 5835 25255 5877 25264
rect 5931 25304 5973 25313
rect 5931 25264 5932 25304
rect 5972 25264 5973 25304
rect 5931 25255 5973 25264
rect 6987 25304 7029 25313
rect 6987 25264 6988 25304
rect 7028 25264 7029 25304
rect 6987 25255 7029 25264
rect 7083 25304 7125 25313
rect 7083 25264 7084 25304
rect 7124 25264 7125 25304
rect 7083 25255 7125 25264
rect 7467 25304 7509 25313
rect 7467 25264 7468 25304
rect 7508 25264 7509 25304
rect 7467 25255 7509 25264
rect 7563 25304 7605 25313
rect 8523 25309 8565 25318
rect 7563 25264 7564 25304
rect 7604 25264 7605 25304
rect 7563 25255 7605 25264
rect 8035 25304 8093 25305
rect 8035 25264 8044 25304
rect 8084 25264 8093 25304
rect 8035 25263 8093 25264
rect 8523 25269 8524 25309
rect 8564 25269 8565 25309
rect 11979 25309 12021 25318
rect 8523 25260 8565 25269
rect 10147 25304 10205 25305
rect 10147 25264 10156 25304
rect 10196 25264 10205 25304
rect 10147 25263 10205 25264
rect 11395 25304 11453 25305
rect 11395 25264 11404 25304
rect 11444 25264 11453 25304
rect 11395 25263 11453 25264
rect 11979 25269 11980 25309
rect 12020 25269 12021 25309
rect 11979 25260 12021 25269
rect 12451 25304 12509 25305
rect 12451 25264 12460 25304
rect 12500 25264 12509 25304
rect 12451 25263 12509 25264
rect 12939 25304 12981 25313
rect 12939 25264 12940 25304
rect 12980 25264 12981 25304
rect 12939 25255 12981 25264
rect 13419 25304 13461 25313
rect 13419 25264 13420 25304
rect 13460 25264 13461 25304
rect 13419 25255 13461 25264
rect 13515 25304 13557 25313
rect 13515 25264 13516 25304
rect 13556 25264 13557 25304
rect 13515 25255 13557 25264
rect 13987 25304 14045 25305
rect 13987 25264 13996 25304
rect 14036 25264 14045 25304
rect 13987 25263 14045 25264
rect 15235 25304 15293 25305
rect 15235 25264 15244 25304
rect 15284 25264 15293 25304
rect 15235 25263 15293 25264
rect 16003 25304 16061 25305
rect 16003 25264 16012 25304
rect 16052 25264 16061 25304
rect 16003 25263 16061 25264
rect 17251 25304 17309 25305
rect 17251 25264 17260 25304
rect 17300 25264 17309 25304
rect 17251 25263 17309 25264
rect 17635 25304 17693 25305
rect 17635 25264 17644 25304
rect 17684 25264 17693 25304
rect 17635 25263 17693 25264
rect 18883 25304 18941 25305
rect 18883 25264 18892 25304
rect 18932 25264 18941 25304
rect 19371 25304 19413 25313
rect 18883 25263 18941 25264
rect 19275 25283 19317 25292
rect 19275 25243 19276 25283
rect 19316 25243 19317 25283
rect 19371 25264 19372 25304
rect 19412 25264 19413 25304
rect 19563 25304 19605 25313
rect 19371 25255 19413 25264
rect 19467 25283 19509 25292
rect 19275 25234 19317 25243
rect 19467 25243 19468 25283
rect 19508 25243 19509 25283
rect 19563 25264 19564 25304
rect 19604 25264 19605 25304
rect 19563 25255 19605 25264
rect 19755 25304 19797 25313
rect 19755 25264 19756 25304
rect 19796 25264 19797 25304
rect 19755 25255 19797 25264
rect 19851 25304 19893 25313
rect 19851 25264 19852 25304
rect 19892 25264 19893 25304
rect 19851 25255 19893 25264
rect 19467 25234 19509 25243
rect 3819 25220 3861 25229
rect 3819 25180 3820 25220
rect 3860 25180 3861 25220
rect 11787 25220 11829 25229
rect 3819 25171 3861 25180
rect 8715 25178 8757 25187
rect 1323 25136 1365 25145
rect 8715 25138 8716 25178
rect 8756 25138 8757 25178
rect 11787 25180 11788 25220
rect 11828 25180 11829 25220
rect 11787 25171 11829 25180
rect 15435 25220 15477 25229
rect 15435 25180 15436 25220
rect 15476 25180 15477 25220
rect 15435 25171 15477 25180
rect 1323 25096 1324 25136
rect 1364 25096 1365 25136
rect 1323 25087 1365 25096
rect 6115 25136 6173 25137
rect 6115 25096 6124 25136
rect 6164 25096 6173 25136
rect 8715 25129 8757 25138
rect 15619 25136 15677 25137
rect 6115 25095 6173 25096
rect 15619 25096 15628 25136
rect 15668 25096 15677 25136
rect 15619 25095 15677 25096
rect 20035 25136 20093 25137
rect 20035 25096 20044 25136
rect 20084 25096 20093 25136
rect 20035 25095 20093 25096
rect 1152 24968 20452 24992
rect 1152 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20452 24968
rect 1152 24904 20452 24928
rect 1419 24800 1461 24809
rect 1419 24760 1420 24800
rect 1460 24760 1461 24800
rect 1419 24751 1461 24760
rect 1699 24800 1757 24801
rect 1699 24760 1708 24800
rect 1748 24760 1757 24800
rect 1699 24759 1757 24760
rect 3435 24800 3477 24809
rect 3435 24760 3436 24800
rect 3476 24760 3477 24800
rect 3435 24751 3477 24760
rect 7563 24800 7605 24809
rect 7563 24760 7564 24800
rect 7604 24760 7605 24800
rect 7563 24751 7605 24760
rect 11403 24800 11445 24809
rect 11403 24760 11404 24800
rect 11444 24760 11445 24800
rect 11403 24751 11445 24760
rect 13035 24800 13077 24809
rect 13035 24760 13036 24800
rect 13076 24760 13077 24800
rect 13035 24751 13077 24760
rect 13323 24800 13365 24809
rect 13323 24760 13324 24800
rect 13364 24760 13365 24800
rect 13323 24751 13365 24760
rect 13795 24800 13853 24801
rect 13795 24760 13804 24800
rect 13844 24760 13853 24800
rect 13795 24759 13853 24760
rect 15435 24800 15477 24809
rect 15435 24760 15436 24800
rect 15476 24760 15477 24800
rect 15435 24751 15477 24760
rect 3723 24716 3765 24725
rect 3723 24676 3724 24716
rect 3764 24676 3765 24716
rect 3723 24667 3765 24676
rect 9579 24716 9621 24725
rect 9579 24676 9580 24716
rect 9620 24676 9621 24716
rect 9579 24667 9621 24676
rect 17739 24716 17781 24725
rect 17739 24676 17740 24716
rect 17780 24676 17781 24716
rect 17739 24667 17781 24676
rect 20235 24716 20277 24725
rect 20235 24676 20236 24716
rect 20276 24676 20277 24716
rect 20235 24667 20277 24676
rect 13899 24653 13941 24662
rect 1323 24632 1365 24641
rect 1323 24592 1324 24632
rect 1364 24592 1365 24632
rect 1323 24583 1365 24592
rect 1515 24632 1557 24641
rect 1515 24592 1516 24632
rect 1556 24592 1557 24632
rect 1515 24583 1557 24592
rect 1987 24632 2045 24633
rect 1987 24592 1996 24632
rect 2036 24592 2045 24632
rect 1987 24591 2045 24592
rect 3235 24632 3293 24633
rect 3235 24592 3244 24632
rect 3284 24592 3293 24632
rect 3235 24591 3293 24592
rect 3915 24627 3957 24636
rect 3915 24587 3916 24627
rect 3956 24587 3957 24627
rect 4387 24632 4445 24633
rect 4387 24592 4396 24632
rect 4436 24592 4445 24632
rect 4387 24591 4445 24592
rect 5355 24632 5397 24641
rect 5355 24592 5356 24632
rect 5396 24592 5397 24632
rect 3915 24578 3957 24587
rect 5355 24583 5397 24592
rect 5451 24632 5493 24641
rect 5451 24592 5452 24632
rect 5492 24592 5493 24632
rect 5451 24583 5493 24592
rect 6115 24632 6173 24633
rect 6115 24592 6124 24632
rect 6164 24592 6173 24632
rect 6115 24591 6173 24592
rect 7363 24632 7421 24633
rect 7363 24592 7372 24632
rect 7412 24592 7421 24632
rect 7363 24591 7421 24592
rect 7851 24632 7893 24641
rect 7851 24592 7852 24632
rect 7892 24592 7893 24632
rect 7851 24583 7893 24592
rect 7947 24632 7989 24641
rect 7947 24592 7948 24632
rect 7988 24592 7989 24632
rect 7947 24583 7989 24592
rect 8331 24632 8373 24641
rect 8331 24592 8332 24632
rect 8372 24592 8373 24632
rect 8331 24583 8373 24592
rect 8899 24632 8957 24633
rect 8899 24592 8908 24632
rect 8948 24592 8957 24632
rect 9955 24632 10013 24633
rect 8899 24591 8957 24592
rect 9387 24618 9429 24627
rect 9387 24578 9388 24618
rect 9428 24578 9429 24618
rect 9955 24592 9964 24632
rect 10004 24592 10013 24632
rect 9955 24591 10013 24592
rect 11203 24632 11261 24633
rect 11203 24592 11212 24632
rect 11252 24592 11261 24632
rect 11203 24591 11261 24592
rect 11587 24632 11645 24633
rect 11587 24592 11596 24632
rect 11636 24592 11645 24632
rect 11587 24591 11645 24592
rect 12835 24632 12893 24633
rect 12835 24592 12844 24632
rect 12884 24592 12893 24632
rect 12835 24591 12893 24592
rect 13227 24632 13269 24641
rect 13227 24592 13228 24632
rect 13268 24592 13269 24632
rect 13227 24583 13269 24592
rect 13419 24632 13461 24641
rect 13419 24592 13420 24632
rect 13460 24592 13461 24632
rect 13419 24583 13461 24592
rect 13515 24632 13557 24641
rect 13515 24592 13516 24632
rect 13556 24592 13557 24632
rect 13899 24613 13900 24653
rect 13940 24613 13941 24653
rect 13899 24604 13941 24613
rect 13995 24632 14037 24641
rect 13515 24583 13557 24592
rect 13995 24592 13996 24632
rect 14036 24592 14037 24632
rect 13995 24583 14037 24592
rect 14091 24632 14133 24641
rect 14091 24592 14092 24632
rect 14132 24592 14133 24632
rect 14091 24583 14133 24592
rect 14283 24632 14325 24641
rect 14283 24592 14284 24632
rect 14324 24592 14325 24632
rect 14283 24583 14325 24592
rect 14475 24632 14517 24641
rect 14475 24592 14476 24632
rect 14516 24592 14517 24632
rect 14475 24583 14517 24592
rect 14571 24632 14613 24641
rect 14571 24592 14572 24632
rect 14612 24592 14613 24632
rect 14571 24583 14613 24592
rect 14851 24632 14909 24633
rect 14851 24592 14860 24632
rect 14900 24592 14909 24632
rect 14851 24591 14909 24592
rect 16011 24632 16053 24641
rect 16011 24592 16012 24632
rect 16052 24592 16053 24632
rect 16011 24583 16053 24592
rect 16107 24632 16149 24641
rect 16107 24592 16108 24632
rect 16148 24592 16149 24632
rect 16107 24583 16149 24592
rect 16491 24632 16533 24641
rect 16491 24592 16492 24632
rect 16532 24592 16533 24632
rect 16491 24583 16533 24592
rect 17059 24632 17117 24633
rect 17059 24592 17068 24632
rect 17108 24592 17117 24632
rect 17059 24591 17117 24592
rect 17547 24627 17589 24636
rect 17547 24587 17548 24627
rect 17588 24587 17589 24627
rect 17547 24578 17589 24587
rect 17931 24632 17973 24641
rect 17931 24592 17932 24632
rect 17972 24592 17973 24632
rect 17931 24583 17973 24592
rect 18123 24632 18165 24641
rect 18123 24592 18124 24632
rect 18164 24592 18165 24632
rect 18123 24583 18165 24592
rect 18211 24632 18269 24633
rect 18211 24592 18220 24632
rect 18260 24592 18269 24632
rect 18603 24632 18645 24641
rect 18211 24591 18269 24592
rect 18507 24613 18549 24622
rect 9387 24569 9429 24578
rect 18507 24573 18508 24613
rect 18548 24573 18549 24613
rect 18603 24592 18604 24632
rect 18644 24592 18645 24632
rect 18603 24583 18645 24592
rect 18987 24632 19029 24641
rect 18987 24592 18988 24632
rect 19028 24592 19029 24632
rect 18987 24583 19029 24592
rect 19555 24632 19613 24633
rect 19555 24592 19564 24632
rect 19604 24592 19613 24632
rect 19555 24591 19613 24592
rect 20043 24618 20085 24627
rect 18507 24564 18549 24573
rect 20043 24578 20044 24618
rect 20084 24578 20085 24618
rect 20043 24569 20085 24578
rect 4875 24548 4917 24557
rect 4875 24508 4876 24548
rect 4916 24508 4917 24548
rect 4875 24499 4917 24508
rect 4971 24548 5013 24557
rect 4971 24508 4972 24548
rect 5012 24508 5013 24548
rect 4971 24499 5013 24508
rect 8427 24548 8469 24557
rect 8427 24508 8428 24548
rect 8468 24508 8469 24548
rect 8427 24499 8469 24508
rect 14763 24548 14805 24557
rect 14763 24508 14764 24548
rect 14804 24508 14805 24548
rect 14763 24499 14805 24508
rect 15235 24548 15293 24549
rect 15235 24508 15244 24548
rect 15284 24508 15293 24548
rect 15235 24507 15293 24508
rect 16587 24548 16629 24557
rect 16587 24508 16588 24548
rect 16628 24508 16629 24548
rect 16587 24499 16629 24508
rect 19083 24548 19125 24557
rect 19083 24508 19084 24548
rect 19124 24508 19125 24548
rect 19083 24499 19125 24508
rect 15627 24464 15669 24473
rect 15627 24424 15628 24464
rect 15668 24424 15669 24464
rect 15627 24415 15669 24424
rect 17931 24380 17973 24389
rect 17931 24340 17932 24380
rect 17972 24340 17973 24380
rect 17931 24331 17973 24340
rect 1152 24212 20352 24236
rect 1152 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 20352 24212
rect 1152 24148 20352 24172
rect 3619 24044 3677 24045
rect 3619 24004 3628 24044
rect 3668 24004 3677 24044
rect 3619 24003 3677 24004
rect 9387 24044 9429 24053
rect 9387 24004 9388 24044
rect 9428 24004 9429 24044
rect 9387 23995 9429 24004
rect 1515 23960 1557 23969
rect 1515 23920 1516 23960
rect 1556 23920 1557 23960
rect 1515 23911 1557 23920
rect 3435 23960 3477 23969
rect 3435 23920 3436 23960
rect 3476 23920 3477 23960
rect 3435 23911 3477 23920
rect 4587 23960 4629 23969
rect 4587 23920 4588 23960
rect 4628 23920 4629 23960
rect 4587 23911 4629 23920
rect 7467 23960 7509 23969
rect 7467 23920 7468 23960
rect 7508 23920 7509 23960
rect 7467 23911 7509 23920
rect 17355 23960 17397 23969
rect 17355 23920 17356 23960
rect 17396 23920 17397 23960
rect 17355 23911 17397 23920
rect 18123 23960 18165 23969
rect 18123 23920 18124 23960
rect 18164 23920 18165 23960
rect 18123 23911 18165 23920
rect 1803 23876 1845 23885
rect 1803 23836 1804 23876
rect 1844 23836 1845 23876
rect 1803 23827 1845 23836
rect 15907 23834 15965 23835
rect 1987 23792 2045 23793
rect 1987 23752 1996 23792
rect 2036 23752 2045 23792
rect 1987 23751 2045 23752
rect 3235 23792 3293 23793
rect 3235 23752 3244 23792
rect 3284 23752 3293 23792
rect 3235 23751 3293 23752
rect 4011 23792 4053 23801
rect 4011 23752 4012 23792
rect 4052 23752 4053 23792
rect 4011 23743 4053 23752
rect 4291 23792 4349 23793
rect 4291 23752 4300 23792
rect 4340 23752 4349 23792
rect 4291 23751 4349 23752
rect 4587 23792 4629 23801
rect 4587 23752 4588 23792
rect 4628 23752 4629 23792
rect 4587 23743 4629 23752
rect 4779 23792 4821 23801
rect 4779 23752 4780 23792
rect 4820 23752 4821 23792
rect 4779 23743 4821 23752
rect 4867 23792 4925 23793
rect 4867 23752 4876 23792
rect 4916 23752 4925 23792
rect 4867 23751 4925 23752
rect 5067 23792 5109 23801
rect 5067 23752 5068 23792
rect 5108 23752 5109 23792
rect 5067 23743 5109 23752
rect 5163 23792 5205 23801
rect 5163 23752 5164 23792
rect 5204 23752 5205 23792
rect 5163 23743 5205 23752
rect 6019 23792 6077 23793
rect 6019 23752 6028 23792
rect 6068 23752 6077 23792
rect 6019 23751 6077 23752
rect 7267 23792 7325 23793
rect 7267 23752 7276 23792
rect 7316 23752 7325 23792
rect 7267 23751 7325 23752
rect 7939 23792 7997 23793
rect 7939 23752 7948 23792
rect 7988 23752 7997 23792
rect 7939 23751 7997 23752
rect 9187 23792 9245 23793
rect 9187 23752 9196 23792
rect 9236 23752 9245 23792
rect 9187 23751 9245 23752
rect 9763 23792 9821 23793
rect 9763 23752 9772 23792
rect 9812 23752 9821 23792
rect 9763 23751 9821 23752
rect 11011 23792 11069 23793
rect 11011 23752 11020 23792
rect 11060 23752 11069 23792
rect 11011 23751 11069 23752
rect 11203 23792 11261 23793
rect 11203 23752 11212 23792
rect 11252 23752 11261 23792
rect 11203 23751 11261 23752
rect 11299 23792 11357 23793
rect 11299 23752 11308 23792
rect 11348 23752 11357 23792
rect 11299 23751 11357 23752
rect 11499 23792 11541 23801
rect 11499 23752 11500 23792
rect 11540 23752 11541 23792
rect 11499 23743 11541 23752
rect 11595 23792 11637 23801
rect 15907 23794 15916 23834
rect 15956 23794 15965 23834
rect 15907 23793 15965 23794
rect 11595 23752 11596 23792
rect 11636 23752 11637 23792
rect 11595 23743 11637 23752
rect 11688 23792 11746 23793
rect 11688 23752 11697 23792
rect 11737 23752 11746 23792
rect 11688 23751 11746 23752
rect 13219 23792 13277 23793
rect 13219 23752 13228 23792
rect 13268 23752 13277 23792
rect 13219 23751 13277 23752
rect 14467 23792 14525 23793
rect 14467 23752 14476 23792
rect 14516 23752 14525 23792
rect 14467 23751 14525 23752
rect 17155 23792 17213 23793
rect 17155 23752 17164 23792
rect 17204 23752 17213 23792
rect 17155 23751 17213 23752
rect 17547 23792 17589 23801
rect 17547 23752 17548 23792
rect 17588 23752 17589 23792
rect 17547 23743 17589 23752
rect 17739 23792 17781 23801
rect 17739 23752 17740 23792
rect 17780 23752 17781 23792
rect 17739 23743 17781 23752
rect 18307 23792 18365 23793
rect 18307 23752 18316 23792
rect 18356 23752 18365 23792
rect 18307 23751 18365 23752
rect 19555 23792 19613 23793
rect 19555 23752 19564 23792
rect 19604 23752 19613 23792
rect 19555 23751 19613 23752
rect 19947 23792 19989 23801
rect 19947 23752 19948 23792
rect 19988 23752 19989 23792
rect 19947 23743 19989 23752
rect 20043 23792 20085 23801
rect 20043 23752 20044 23792
rect 20084 23752 20085 23792
rect 20043 23743 20085 23752
rect 3915 23708 3957 23717
rect 3915 23668 3916 23708
rect 3956 23668 3957 23708
rect 3915 23659 3957 23668
rect 5347 23624 5405 23625
rect 5347 23584 5356 23624
rect 5396 23584 5405 23624
rect 5347 23583 5405 23584
rect 9579 23624 9621 23633
rect 9579 23584 9580 23624
rect 9620 23584 9621 23624
rect 9579 23575 9621 23584
rect 11683 23624 11741 23625
rect 11683 23584 11692 23624
rect 11732 23584 11741 23624
rect 11683 23583 11741 23584
rect 14667 23624 14709 23633
rect 14667 23584 14668 23624
rect 14708 23584 14709 23624
rect 14667 23575 14709 23584
rect 15619 23624 15677 23625
rect 15619 23584 15628 23624
rect 15668 23584 15677 23624
rect 15619 23583 15677 23584
rect 17643 23624 17685 23633
rect 17643 23584 17644 23624
rect 17684 23584 17685 23624
rect 17643 23575 17685 23584
rect 19747 23624 19805 23625
rect 19747 23584 19756 23624
rect 19796 23584 19805 23624
rect 19747 23583 19805 23584
rect 1152 23456 20452 23480
rect 1152 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20452 23456
rect 1152 23392 20452 23416
rect 4011 23288 4053 23297
rect 4011 23248 4012 23288
rect 4052 23248 4053 23288
rect 4011 23239 4053 23248
rect 9291 23288 9333 23297
rect 9291 23248 9292 23288
rect 9332 23248 9333 23288
rect 9291 23239 9333 23248
rect 9675 23288 9717 23297
rect 9675 23248 9676 23288
rect 9716 23248 9717 23288
rect 9675 23239 9717 23248
rect 14859 23288 14901 23297
rect 14859 23248 14860 23288
rect 14900 23248 14901 23288
rect 14859 23239 14901 23248
rect 18891 23288 18933 23297
rect 18891 23248 18892 23288
rect 18932 23248 18933 23288
rect 18891 23239 18933 23248
rect 20131 23288 20189 23289
rect 20131 23248 20140 23288
rect 20180 23248 20189 23288
rect 20131 23247 20189 23248
rect 3147 23204 3189 23213
rect 3147 23164 3148 23204
rect 3188 23164 3189 23204
rect 3147 23155 3189 23164
rect 3627 23204 3669 23213
rect 3627 23164 3628 23204
rect 3668 23164 3669 23204
rect 3627 23155 3669 23164
rect 5931 23204 5973 23213
rect 5931 23164 5932 23204
rect 5972 23164 5973 23204
rect 5931 23155 5973 23164
rect 7563 23204 7605 23213
rect 7563 23164 7564 23204
rect 7604 23164 7605 23204
rect 7563 23155 7605 23164
rect 12843 23204 12885 23213
rect 12843 23164 12844 23204
rect 12884 23164 12885 23204
rect 12843 23155 12885 23164
rect 1699 23120 1757 23121
rect 1699 23080 1708 23120
rect 1748 23080 1757 23120
rect 1699 23079 1757 23080
rect 2947 23120 3005 23121
rect 2947 23080 2956 23120
rect 2996 23080 3005 23120
rect 2947 23079 3005 23080
rect 3339 23120 3381 23129
rect 3339 23080 3340 23120
rect 3380 23080 3381 23120
rect 3339 23071 3381 23080
rect 3435 23120 3477 23129
rect 3435 23080 3436 23120
rect 3476 23080 3477 23120
rect 3435 23071 3477 23080
rect 3531 23120 3573 23129
rect 3531 23080 3532 23120
rect 3572 23080 3573 23120
rect 3531 23071 3573 23080
rect 3819 23120 3861 23129
rect 3819 23080 3820 23120
rect 3860 23080 3861 23120
rect 3819 23071 3861 23080
rect 4107 23120 4149 23129
rect 4107 23080 4108 23120
rect 4148 23080 4149 23120
rect 4107 23071 4149 23080
rect 4483 23120 4541 23121
rect 4483 23080 4492 23120
rect 4532 23080 4541 23120
rect 4483 23079 4541 23080
rect 5731 23120 5789 23121
rect 5731 23080 5740 23120
rect 5780 23080 5789 23120
rect 5731 23079 5789 23080
rect 6499 23120 6557 23121
rect 6499 23080 6508 23120
rect 6548 23080 6557 23120
rect 6499 23079 6557 23080
rect 6795 23120 6837 23129
rect 6795 23080 6796 23120
rect 6836 23080 6837 23120
rect 6795 23071 6837 23080
rect 6891 23120 6933 23129
rect 6891 23080 6892 23120
rect 6932 23080 6933 23120
rect 6891 23071 6933 23080
rect 7467 23120 7509 23129
rect 7467 23080 7468 23120
rect 7508 23080 7509 23120
rect 7467 23071 7509 23080
rect 7659 23120 7701 23129
rect 7659 23080 7660 23120
rect 7700 23080 7701 23120
rect 7659 23071 7701 23080
rect 7747 23120 7805 23121
rect 7747 23080 7756 23120
rect 7796 23080 7805 23120
rect 7747 23079 7805 23080
rect 7947 23120 7989 23129
rect 7947 23080 7948 23120
rect 7988 23080 7989 23120
rect 7947 23071 7989 23080
rect 8139 23120 8181 23129
rect 8139 23080 8140 23120
rect 8180 23080 8181 23120
rect 8139 23071 8181 23080
rect 8227 23120 8285 23121
rect 8227 23080 8236 23120
rect 8276 23080 8285 23120
rect 8227 23079 8285 23080
rect 8715 23120 8757 23129
rect 8715 23080 8716 23120
rect 8756 23080 8757 23120
rect 8715 23071 8757 23080
rect 8907 23120 8949 23129
rect 8907 23080 8908 23120
rect 8948 23080 8949 23120
rect 8907 23071 8949 23080
rect 9003 23120 9045 23129
rect 9003 23080 9004 23120
rect 9044 23080 9045 23120
rect 9003 23071 9045 23080
rect 9195 23120 9237 23129
rect 9195 23080 9196 23120
rect 9236 23080 9237 23120
rect 9195 23071 9237 23080
rect 9387 23120 9429 23129
rect 9387 23080 9388 23120
rect 9428 23080 9429 23120
rect 9387 23071 9429 23080
rect 9483 23120 9525 23129
rect 9483 23080 9484 23120
rect 9524 23080 9525 23120
rect 9483 23071 9525 23080
rect 9859 23120 9917 23121
rect 9859 23080 9868 23120
rect 9908 23080 9917 23120
rect 9859 23079 9917 23080
rect 11107 23120 11165 23121
rect 11107 23080 11116 23120
rect 11156 23080 11165 23120
rect 11107 23079 11165 23080
rect 11395 23120 11453 23121
rect 11395 23080 11404 23120
rect 11444 23080 11453 23120
rect 11395 23079 11453 23080
rect 12643 23120 12701 23121
rect 12643 23080 12652 23120
rect 12692 23080 12701 23120
rect 12643 23079 12701 23080
rect 13131 23120 13173 23129
rect 13131 23080 13132 23120
rect 13172 23080 13173 23120
rect 13131 23071 13173 23080
rect 13227 23120 13269 23129
rect 13227 23080 13228 23120
rect 13268 23080 13269 23120
rect 13227 23071 13269 23080
rect 13611 23120 13653 23129
rect 13611 23080 13612 23120
rect 13652 23080 13653 23120
rect 13611 23071 13653 23080
rect 14179 23120 14237 23121
rect 14179 23080 14188 23120
rect 14228 23080 14237 23120
rect 14179 23079 14237 23080
rect 14667 23115 14709 23124
rect 14667 23075 14668 23115
rect 14708 23075 14709 23115
rect 15907 23120 15965 23121
rect 15907 23080 15916 23120
rect 15956 23080 15965 23120
rect 15907 23079 15965 23080
rect 16011 23120 16053 23129
rect 16011 23080 16012 23120
rect 16052 23080 16053 23120
rect 14667 23066 14709 23075
rect 16011 23071 16053 23080
rect 16203 23120 16245 23129
rect 16203 23080 16204 23120
rect 16244 23080 16245 23120
rect 16203 23071 16245 23080
rect 16579 23120 16637 23121
rect 16579 23080 16588 23120
rect 16628 23080 16637 23120
rect 16579 23079 16637 23080
rect 16875 23120 16917 23129
rect 16875 23080 16876 23120
rect 16916 23080 16917 23120
rect 16875 23071 16917 23080
rect 16971 23120 17013 23129
rect 16971 23080 16972 23120
rect 17012 23080 17013 23120
rect 16971 23071 17013 23080
rect 17443 23120 17501 23121
rect 17443 23080 17452 23120
rect 17492 23080 17501 23120
rect 17443 23079 17501 23080
rect 18691 23120 18749 23121
rect 18691 23080 18700 23120
rect 18740 23080 18749 23120
rect 18691 23079 18749 23080
rect 19112 23120 19170 23121
rect 19112 23080 19121 23120
rect 19161 23080 19170 23120
rect 19112 23079 19170 23080
rect 19275 23120 19317 23129
rect 19275 23080 19276 23120
rect 19316 23080 19317 23120
rect 19275 23071 19317 23080
rect 19371 23120 19413 23129
rect 19371 23080 19372 23120
rect 19412 23080 19413 23120
rect 19371 23071 19413 23080
rect 19555 23120 19613 23121
rect 19555 23080 19564 23120
rect 19604 23080 19613 23120
rect 19555 23079 19613 23080
rect 19651 23120 19709 23121
rect 19651 23080 19660 23120
rect 19700 23080 19709 23120
rect 19651 23079 19709 23080
rect 19851 23120 19893 23129
rect 19851 23080 19852 23120
rect 19892 23080 19893 23120
rect 19851 23071 19893 23080
rect 19947 23120 19989 23129
rect 19947 23080 19948 23120
rect 19988 23080 19989 23120
rect 19947 23071 19989 23080
rect 13707 23036 13749 23045
rect 13707 22996 13708 23036
rect 13748 22996 13749 23036
rect 13707 22987 13749 22996
rect 15235 23036 15293 23037
rect 15235 22996 15244 23036
rect 15284 22996 15293 23036
rect 15235 22995 15293 22996
rect 7947 22952 7989 22961
rect 7947 22912 7948 22952
rect 7988 22912 7989 22952
rect 7947 22903 7989 22912
rect 8995 22952 9053 22953
rect 8995 22912 9004 22952
rect 9044 22912 9053 22952
rect 8995 22911 9053 22912
rect 15627 22952 15669 22961
rect 15627 22912 15628 22952
rect 15668 22912 15669 22952
rect 15627 22903 15669 22912
rect 17251 22952 17309 22953
rect 17251 22912 17260 22952
rect 17300 22912 17309 22952
rect 17251 22911 17309 22912
rect 7171 22868 7229 22869
rect 7171 22828 7180 22868
rect 7220 22828 7229 22868
rect 7171 22827 7229 22828
rect 15435 22868 15477 22877
rect 15435 22828 15436 22868
rect 15476 22828 15477 22868
rect 15435 22819 15477 22828
rect 16203 22868 16245 22877
rect 16203 22828 16204 22868
rect 16244 22828 16245 22868
rect 16203 22819 16245 22828
rect 19659 22868 19701 22877
rect 19659 22828 19660 22868
rect 19700 22828 19701 22868
rect 19659 22819 19701 22828
rect 1152 22700 20352 22724
rect 1152 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 20352 22700
rect 1152 22636 20352 22660
rect 2667 22532 2709 22541
rect 2667 22492 2668 22532
rect 2708 22492 2709 22532
rect 2667 22483 2709 22492
rect 9579 22532 9621 22541
rect 9579 22492 9580 22532
rect 9620 22492 9621 22532
rect 9579 22483 9621 22492
rect 18123 22532 18165 22541
rect 18123 22492 18124 22532
rect 18164 22492 18165 22532
rect 18123 22483 18165 22492
rect 20043 22532 20085 22541
rect 20043 22492 20044 22532
rect 20084 22492 20085 22532
rect 20043 22483 20085 22492
rect 5451 22448 5493 22457
rect 5451 22408 5452 22448
rect 5492 22408 5493 22448
rect 5451 22399 5493 22408
rect 12363 22448 12405 22457
rect 12363 22408 12364 22448
rect 12404 22408 12405 22448
rect 12363 22399 12405 22408
rect 13227 22364 13269 22373
rect 13227 22324 13228 22364
rect 13268 22324 13269 22364
rect 13227 22315 13269 22324
rect 3051 22299 3093 22308
rect 1219 22280 1277 22281
rect 1219 22240 1228 22280
rect 1268 22240 1277 22280
rect 1219 22239 1277 22240
rect 2467 22280 2525 22281
rect 2467 22240 2476 22280
rect 2516 22240 2525 22280
rect 3051 22259 3052 22299
rect 3092 22259 3093 22299
rect 4587 22294 4629 22303
rect 7371 22299 7413 22308
rect 3051 22250 3093 22259
rect 3147 22280 3189 22289
rect 2467 22239 2525 22240
rect 3147 22240 3148 22280
rect 3188 22240 3189 22280
rect 3147 22231 3189 22240
rect 3531 22280 3573 22289
rect 3531 22240 3532 22280
rect 3572 22240 3573 22280
rect 3531 22231 3573 22240
rect 3627 22280 3669 22289
rect 3627 22240 3628 22280
rect 3668 22240 3669 22280
rect 3627 22231 3669 22240
rect 4099 22280 4157 22281
rect 4099 22240 4108 22280
rect 4148 22240 4157 22280
rect 4587 22254 4588 22294
rect 4628 22254 4629 22294
rect 4587 22245 4629 22254
rect 5259 22280 5301 22289
rect 4099 22239 4157 22240
rect 5259 22240 5260 22280
rect 5300 22240 5301 22280
rect 5259 22231 5301 22240
rect 5451 22280 5493 22289
rect 5451 22240 5452 22280
rect 5492 22240 5493 22280
rect 5451 22231 5493 22240
rect 5835 22285 5877 22294
rect 5835 22245 5836 22285
rect 5876 22245 5877 22285
rect 5835 22236 5877 22245
rect 6307 22280 6365 22281
rect 6307 22240 6316 22280
rect 6356 22240 6365 22280
rect 6307 22239 6365 22240
rect 6795 22280 6837 22289
rect 6795 22240 6796 22280
rect 6836 22240 6837 22280
rect 6795 22231 6837 22240
rect 6891 22280 6933 22289
rect 6891 22240 6892 22280
rect 6932 22240 6933 22280
rect 6891 22231 6933 22240
rect 7275 22280 7317 22289
rect 7275 22240 7276 22280
rect 7316 22240 7317 22280
rect 7371 22259 7372 22299
rect 7412 22259 7413 22299
rect 12747 22299 12789 22308
rect 7371 22250 7413 22259
rect 7851 22280 7893 22289
rect 7275 22231 7317 22240
rect 7851 22240 7852 22280
rect 7892 22240 7893 22280
rect 7851 22231 7893 22240
rect 7947 22280 7989 22289
rect 7947 22240 7948 22280
rect 7988 22240 7989 22280
rect 7947 22231 7989 22240
rect 8131 22280 8189 22281
rect 8131 22240 8140 22280
rect 8180 22240 8189 22280
rect 8131 22239 8189 22240
rect 9379 22280 9437 22281
rect 9379 22240 9388 22280
rect 9428 22240 9437 22280
rect 9379 22239 9437 22240
rect 9763 22280 9821 22281
rect 9763 22240 9772 22280
rect 9812 22240 9821 22280
rect 9763 22239 9821 22240
rect 9859 22280 9917 22281
rect 9859 22240 9868 22280
rect 9908 22240 9917 22280
rect 9859 22239 9917 22240
rect 10059 22280 10101 22289
rect 10059 22240 10060 22280
rect 10100 22240 10101 22280
rect 10059 22231 10101 22240
rect 10155 22280 10197 22289
rect 10155 22240 10156 22280
rect 10196 22240 10197 22280
rect 10155 22231 10197 22240
rect 10248 22280 10306 22281
rect 10248 22240 10257 22280
rect 10297 22240 10306 22280
rect 10248 22239 10306 22240
rect 10915 22280 10973 22281
rect 10915 22240 10924 22280
rect 10964 22240 10973 22280
rect 10915 22239 10973 22240
rect 12163 22280 12221 22281
rect 12163 22240 12172 22280
rect 12212 22240 12221 22280
rect 12163 22239 12221 22240
rect 12651 22280 12693 22289
rect 12651 22240 12652 22280
rect 12692 22240 12693 22280
rect 12747 22259 12748 22299
rect 12788 22259 12789 22299
rect 12747 22250 12789 22259
rect 13131 22280 13173 22289
rect 14187 22285 14229 22294
rect 12651 22231 12693 22240
rect 13131 22240 13132 22280
rect 13172 22240 13173 22280
rect 13131 22231 13173 22240
rect 13699 22280 13757 22281
rect 13699 22240 13708 22280
rect 13748 22240 13757 22280
rect 13699 22239 13757 22240
rect 14187 22245 14188 22285
rect 14228 22245 14229 22285
rect 14187 22236 14229 22245
rect 14571 22280 14613 22289
rect 14571 22240 14572 22280
rect 14612 22240 14613 22280
rect 14571 22231 14613 22240
rect 14763 22280 14805 22289
rect 14763 22240 14764 22280
rect 14804 22240 14805 22280
rect 14763 22231 14805 22240
rect 14859 22280 14901 22289
rect 14859 22240 14860 22280
rect 14900 22240 14901 22280
rect 14859 22231 14901 22240
rect 15051 22280 15093 22289
rect 15051 22240 15052 22280
rect 15092 22240 15093 22280
rect 15051 22231 15093 22240
rect 15147 22280 15189 22289
rect 15147 22240 15148 22280
rect 15188 22240 15189 22280
rect 15147 22231 15189 22240
rect 15998 22280 16056 22281
rect 15998 22240 16007 22280
rect 16047 22240 16056 22280
rect 15998 22239 16056 22240
rect 16107 22280 16149 22289
rect 16107 22240 16108 22280
rect 16148 22240 16149 22280
rect 16107 22231 16149 22240
rect 16203 22280 16245 22289
rect 16203 22240 16204 22280
rect 16244 22240 16245 22280
rect 16203 22231 16245 22240
rect 16387 22280 16445 22281
rect 16387 22240 16396 22280
rect 16436 22240 16445 22280
rect 16387 22239 16445 22240
rect 16483 22280 16541 22281
rect 16483 22240 16492 22280
rect 16532 22240 16541 22280
rect 16483 22239 16541 22240
rect 16675 22280 16733 22281
rect 16675 22240 16684 22280
rect 16724 22240 16733 22280
rect 16675 22239 16733 22240
rect 17923 22280 17981 22281
rect 17923 22240 17932 22280
rect 17972 22240 17981 22280
rect 17923 22239 17981 22240
rect 18595 22280 18653 22281
rect 18595 22240 18604 22280
rect 18644 22240 18653 22280
rect 18595 22239 18653 22240
rect 19843 22280 19901 22281
rect 19843 22240 19852 22280
rect 19892 22240 19901 22280
rect 19843 22239 19901 22240
rect 4779 22196 4821 22205
rect 4779 22156 4780 22196
rect 4820 22156 4821 22196
rect 4779 22147 4821 22156
rect 5643 22196 5685 22205
rect 5643 22156 5644 22196
rect 5684 22156 5685 22196
rect 5643 22147 5685 22156
rect 7651 22112 7709 22113
rect 7651 22072 7660 22112
rect 7700 22072 7709 22112
rect 7651 22071 7709 22072
rect 10147 22112 10205 22113
rect 10147 22072 10156 22112
rect 10196 22072 10205 22112
rect 10147 22071 10205 22072
rect 14379 22112 14421 22121
rect 14379 22072 14380 22112
rect 14420 22072 14421 22112
rect 14379 22063 14421 22072
rect 14667 22112 14709 22121
rect 14667 22072 14668 22112
rect 14708 22072 14709 22112
rect 14667 22063 14709 22072
rect 15331 22112 15389 22113
rect 15331 22072 15340 22112
rect 15380 22072 15389 22112
rect 15331 22071 15389 22072
rect 15619 22112 15677 22113
rect 15619 22072 15628 22112
rect 15668 22072 15677 22112
rect 15619 22071 15677 22072
rect 16099 22112 16157 22113
rect 16099 22072 16108 22112
rect 16148 22072 16157 22112
rect 16099 22071 16157 22072
rect 18411 22112 18453 22121
rect 18411 22072 18412 22112
rect 18452 22072 18453 22112
rect 18411 22063 18453 22072
rect 1152 21944 20452 21968
rect 1152 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20452 21944
rect 1152 21880 20452 21904
rect 2955 21776 2997 21785
rect 2955 21736 2956 21776
rect 2996 21736 2997 21776
rect 2955 21727 2997 21736
rect 3427 21776 3485 21777
rect 3427 21736 3436 21776
rect 3476 21736 3485 21776
rect 3427 21735 3485 21736
rect 3907 21776 3965 21777
rect 3907 21736 3916 21776
rect 3956 21736 3965 21776
rect 3907 21735 3965 21736
rect 4675 21776 4733 21777
rect 4675 21736 4684 21776
rect 4724 21736 4733 21776
rect 4675 21735 4733 21736
rect 6891 21776 6933 21785
rect 6891 21736 6892 21776
rect 6932 21736 6933 21776
rect 6891 21727 6933 21736
rect 9483 21776 9525 21785
rect 9483 21736 9484 21776
rect 9524 21736 9525 21776
rect 9483 21727 9525 21736
rect 9955 21776 10013 21777
rect 9955 21736 9964 21776
rect 10004 21736 10013 21776
rect 9955 21735 10013 21736
rect 11299 21776 11357 21777
rect 11299 21736 11308 21776
rect 11348 21736 11357 21776
rect 11299 21735 11357 21736
rect 14659 21776 14717 21777
rect 14659 21736 14668 21776
rect 14708 21736 14717 21776
rect 14659 21735 14717 21736
rect 19083 21776 19125 21785
rect 19083 21736 19084 21776
rect 19124 21736 19125 21776
rect 19083 21727 19125 21736
rect 19267 21776 19325 21777
rect 19267 21736 19276 21776
rect 19316 21736 19325 21776
rect 19267 21735 19325 21736
rect 7563 21692 7605 21701
rect 7563 21652 7564 21692
rect 7604 21652 7605 21692
rect 7563 21643 7605 21652
rect 13995 21692 14037 21701
rect 13995 21652 13996 21692
rect 14036 21652 14037 21692
rect 13995 21643 14037 21652
rect 1507 21608 1565 21609
rect 1507 21568 1516 21608
rect 1556 21568 1565 21608
rect 1507 21567 1565 21568
rect 2755 21608 2813 21609
rect 2755 21568 2764 21608
rect 2804 21568 2813 21608
rect 2755 21567 2813 21568
rect 3627 21608 3669 21617
rect 3627 21568 3628 21608
rect 3668 21568 3669 21608
rect 3627 21559 3669 21568
rect 3723 21608 3765 21617
rect 3723 21568 3724 21608
rect 3764 21568 3765 21608
rect 3723 21559 3765 21568
rect 4011 21608 4053 21617
rect 4011 21568 4012 21608
rect 4052 21568 4053 21608
rect 4011 21559 4053 21568
rect 4107 21608 4149 21617
rect 4107 21568 4108 21608
rect 4148 21568 4149 21608
rect 4107 21559 4149 21568
rect 4203 21608 4245 21617
rect 4203 21568 4204 21608
rect 4244 21568 4245 21608
rect 4203 21559 4245 21568
rect 4395 21608 4437 21617
rect 4395 21568 4396 21608
rect 4436 21568 4437 21608
rect 4395 21559 4437 21568
rect 4491 21608 4533 21617
rect 4491 21568 4492 21608
rect 4532 21568 4533 21608
rect 4491 21559 4533 21568
rect 5443 21608 5501 21609
rect 5443 21568 5452 21608
rect 5492 21568 5501 21608
rect 5443 21567 5501 21568
rect 6691 21608 6749 21609
rect 6691 21568 6700 21608
rect 6740 21568 6749 21608
rect 6691 21567 6749 21568
rect 7171 21608 7229 21609
rect 7171 21568 7180 21608
rect 7220 21568 7229 21608
rect 7171 21567 7229 21568
rect 7467 21608 7509 21617
rect 7467 21568 7468 21608
rect 7508 21568 7509 21608
rect 7467 21559 7509 21568
rect 8035 21608 8093 21609
rect 8035 21568 8044 21608
rect 8084 21568 8093 21608
rect 8035 21567 8093 21568
rect 9283 21608 9341 21609
rect 9283 21568 9292 21608
rect 9332 21568 9341 21608
rect 9283 21567 9341 21568
rect 9675 21608 9717 21617
rect 9675 21568 9676 21608
rect 9716 21568 9717 21608
rect 9675 21559 9717 21568
rect 9771 21608 9813 21617
rect 9771 21568 9772 21608
rect 9812 21568 9813 21608
rect 9771 21559 9813 21568
rect 11019 21608 11061 21617
rect 11019 21568 11020 21608
rect 11060 21568 11061 21608
rect 11019 21559 11061 21568
rect 11115 21608 11157 21617
rect 11115 21568 11116 21608
rect 11156 21568 11157 21608
rect 11115 21559 11157 21568
rect 12547 21608 12605 21609
rect 12547 21568 12556 21608
rect 12596 21568 12605 21608
rect 12547 21567 12605 21568
rect 13795 21608 13853 21609
rect 13795 21568 13804 21608
rect 13844 21568 13853 21608
rect 13795 21567 13853 21568
rect 14467 21608 14525 21609
rect 14467 21568 14476 21608
rect 14516 21568 14525 21608
rect 14467 21567 14525 21568
rect 14563 21608 14621 21609
rect 14563 21568 14572 21608
rect 14612 21568 14621 21608
rect 14563 21567 14621 21568
rect 14763 21608 14805 21617
rect 14763 21568 14764 21608
rect 14804 21568 14805 21608
rect 14763 21559 14805 21568
rect 14859 21608 14901 21617
rect 14859 21568 14860 21608
rect 14900 21568 14901 21608
rect 14859 21559 14901 21568
rect 15006 21608 15064 21609
rect 15006 21568 15015 21608
rect 15055 21568 15064 21608
rect 15006 21567 15064 21568
rect 15243 21608 15285 21617
rect 15243 21568 15244 21608
rect 15284 21568 15285 21608
rect 15243 21559 15285 21568
rect 15331 21608 15389 21609
rect 15331 21568 15340 21608
rect 15380 21568 15389 21608
rect 15331 21567 15389 21568
rect 15523 21608 15581 21609
rect 15523 21568 15532 21608
rect 15572 21568 15581 21608
rect 15523 21567 15581 21568
rect 16771 21608 16829 21609
rect 16771 21568 16780 21608
rect 16820 21568 16829 21608
rect 16771 21567 16829 21568
rect 17163 21608 17205 21617
rect 17163 21568 17164 21608
rect 17204 21568 17205 21608
rect 17163 21559 17205 21568
rect 17259 21608 17301 21617
rect 17259 21568 17260 21608
rect 17300 21568 17301 21608
rect 17259 21559 17301 21568
rect 17451 21608 17493 21617
rect 17451 21568 17452 21608
rect 17492 21568 17493 21608
rect 17451 21559 17493 21568
rect 17635 21608 17693 21609
rect 17635 21568 17644 21608
rect 17684 21568 17693 21608
rect 17635 21567 17693 21568
rect 18883 21608 18941 21609
rect 18883 21568 18892 21608
rect 18932 21568 18941 21608
rect 18883 21567 18941 21568
rect 19467 21608 19509 21617
rect 19467 21568 19468 21608
rect 19508 21568 19509 21608
rect 19467 21559 19509 21568
rect 19563 21608 19605 21617
rect 19563 21568 19564 21608
rect 19604 21568 19605 21608
rect 19563 21559 19605 21568
rect 19851 21608 19893 21617
rect 19851 21568 19852 21608
rect 19892 21568 19893 21608
rect 19851 21559 19893 21568
rect 19947 21608 19989 21617
rect 19947 21568 19948 21608
rect 19988 21568 19989 21608
rect 19947 21559 19989 21568
rect 20139 21608 20181 21617
rect 20139 21568 20140 21608
rect 20180 21568 20181 21608
rect 20139 21559 20181 21568
rect 7843 21440 7901 21441
rect 7843 21400 7852 21440
rect 7892 21400 7901 21440
rect 7843 21399 7901 21400
rect 17155 21440 17213 21441
rect 17155 21400 17164 21440
rect 17204 21400 17213 21440
rect 17155 21399 17213 21400
rect 19843 21440 19901 21441
rect 19843 21400 19852 21440
rect 19892 21400 19901 21440
rect 19843 21399 19901 21400
rect 16971 21356 17013 21365
rect 16971 21316 16972 21356
rect 17012 21316 17013 21356
rect 16971 21307 17013 21316
rect 1152 21188 20352 21212
rect 1152 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 20352 21188
rect 1152 21124 20352 21148
rect 2667 21020 2709 21029
rect 2667 20980 2668 21020
rect 2708 20980 2709 21020
rect 2667 20971 2709 20980
rect 6891 21020 6933 21029
rect 6891 20980 6892 21020
rect 6932 20980 6933 21020
rect 6891 20971 6933 20980
rect 14859 21020 14901 21029
rect 14859 20980 14860 21020
rect 14900 20980 14901 21020
rect 14859 20971 14901 20980
rect 17067 21020 17109 21029
rect 17067 20980 17068 21020
rect 17108 20980 17109 21020
rect 17067 20971 17109 20980
rect 17451 21020 17493 21029
rect 17451 20980 17452 21020
rect 17492 20980 17493 21020
rect 17451 20971 17493 20980
rect 20235 21020 20277 21029
rect 20235 20980 20236 21020
rect 20276 20980 20277 21020
rect 20235 20971 20277 20980
rect 11019 20936 11061 20945
rect 11019 20896 11020 20936
rect 11060 20896 11061 20936
rect 11019 20887 11061 20896
rect 12931 20936 12989 20937
rect 12931 20896 12940 20936
rect 12980 20896 12989 20936
rect 12931 20895 12989 20896
rect 13131 20936 13173 20945
rect 13131 20896 13132 20936
rect 13172 20896 13173 20936
rect 13131 20887 13173 20896
rect 17643 20936 17685 20945
rect 17643 20896 17644 20936
rect 17684 20896 17685 20936
rect 17643 20887 17685 20896
rect 3435 20852 3477 20861
rect 3435 20812 3436 20852
rect 3476 20812 3477 20852
rect 3435 20803 3477 20812
rect 3531 20852 3573 20861
rect 3531 20812 3532 20852
rect 3572 20812 3573 20852
rect 3531 20803 3573 20812
rect 17251 20852 17309 20853
rect 17251 20812 17260 20852
rect 17300 20812 17309 20852
rect 17251 20811 17309 20812
rect 11752 20783 11794 20792
rect 1219 20768 1277 20769
rect 1219 20728 1228 20768
rect 1268 20728 1277 20768
rect 1219 20727 1277 20728
rect 2467 20768 2525 20769
rect 2467 20728 2476 20768
rect 2516 20728 2525 20768
rect 2467 20727 2525 20728
rect 2955 20768 2997 20777
rect 2955 20728 2956 20768
rect 2996 20728 2997 20768
rect 2955 20719 2997 20728
rect 3051 20768 3093 20777
rect 4491 20773 4533 20782
rect 3051 20728 3052 20768
rect 3092 20728 3093 20768
rect 3051 20719 3093 20728
rect 4003 20768 4061 20769
rect 4003 20728 4012 20768
rect 4052 20728 4061 20768
rect 4003 20727 4061 20728
rect 4491 20733 4492 20773
rect 4532 20733 4533 20773
rect 4491 20724 4533 20733
rect 5443 20768 5501 20769
rect 5443 20728 5452 20768
rect 5492 20728 5501 20768
rect 5443 20727 5501 20728
rect 6691 20768 6749 20769
rect 6691 20728 6700 20768
rect 6740 20728 6749 20768
rect 6691 20727 6749 20728
rect 7075 20768 7133 20769
rect 7075 20728 7084 20768
rect 7124 20728 7133 20768
rect 7075 20727 7133 20728
rect 8323 20768 8381 20769
rect 8323 20728 8332 20768
rect 8372 20728 8381 20768
rect 8323 20727 8381 20728
rect 9571 20768 9629 20769
rect 9571 20728 9580 20768
rect 9620 20728 9629 20768
rect 9571 20727 9629 20728
rect 10819 20768 10877 20769
rect 10819 20728 10828 20768
rect 10868 20728 10877 20768
rect 10819 20727 10877 20728
rect 11203 20768 11261 20769
rect 11203 20728 11212 20768
rect 11252 20728 11261 20768
rect 11203 20727 11261 20728
rect 11299 20768 11357 20769
rect 11299 20728 11308 20768
rect 11348 20728 11357 20768
rect 11299 20727 11357 20728
rect 11499 20768 11541 20777
rect 11499 20728 11500 20768
rect 11540 20728 11541 20768
rect 11499 20719 11541 20728
rect 11595 20768 11637 20777
rect 11595 20728 11596 20768
rect 11636 20728 11637 20768
rect 11752 20743 11753 20783
rect 11793 20743 11794 20783
rect 11752 20734 11794 20743
rect 11979 20768 12021 20777
rect 11595 20719 11637 20728
rect 11979 20728 11980 20768
rect 12020 20728 12021 20768
rect 11979 20719 12021 20728
rect 12075 20768 12117 20777
rect 12075 20728 12076 20768
rect 12116 20728 12117 20768
rect 12075 20719 12117 20728
rect 12651 20768 12693 20777
rect 12651 20728 12652 20768
rect 12692 20728 12693 20768
rect 12651 20719 12693 20728
rect 12843 20768 12885 20777
rect 12843 20728 12844 20768
rect 12884 20728 12885 20768
rect 12843 20719 12885 20728
rect 12939 20768 12981 20777
rect 12939 20728 12940 20768
rect 12980 20728 12981 20768
rect 12939 20719 12981 20728
rect 13411 20768 13469 20769
rect 13411 20728 13420 20768
rect 13460 20728 13469 20768
rect 13411 20727 13469 20728
rect 14659 20768 14717 20769
rect 14659 20728 14668 20768
rect 14708 20728 14717 20768
rect 14659 20727 14717 20728
rect 15339 20768 15381 20777
rect 15339 20728 15340 20768
rect 15380 20728 15381 20768
rect 15339 20719 15381 20728
rect 15435 20768 15477 20777
rect 15435 20728 15436 20768
rect 15476 20728 15477 20768
rect 15435 20719 15477 20728
rect 15619 20768 15677 20769
rect 15619 20728 15628 20768
rect 15668 20728 15677 20768
rect 15619 20727 15677 20728
rect 16867 20768 16925 20769
rect 16867 20728 16876 20768
rect 16916 20728 16925 20768
rect 16867 20727 16925 20728
rect 18014 20768 18072 20769
rect 18014 20728 18023 20768
rect 18063 20728 18072 20768
rect 18014 20727 18072 20728
rect 18123 20768 18165 20777
rect 18123 20728 18124 20768
rect 18164 20728 18165 20768
rect 18123 20719 18165 20728
rect 18219 20768 18261 20777
rect 18219 20728 18220 20768
rect 18260 20728 18261 20768
rect 18219 20719 18261 20728
rect 18403 20768 18461 20769
rect 18403 20728 18412 20768
rect 18452 20728 18461 20768
rect 18403 20727 18461 20728
rect 18499 20768 18557 20769
rect 18499 20728 18508 20768
rect 18548 20728 18557 20768
rect 18499 20727 18557 20728
rect 18787 20768 18845 20769
rect 18787 20728 18796 20768
rect 18836 20728 18845 20768
rect 18787 20727 18845 20728
rect 20035 20768 20093 20769
rect 20035 20728 20044 20768
rect 20084 20728 20093 20768
rect 20035 20727 20093 20728
rect 4683 20684 4725 20693
rect 4683 20644 4684 20684
rect 4724 20644 4725 20684
rect 4683 20635 4725 20644
rect 6891 20600 6933 20609
rect 6891 20560 6892 20600
rect 6932 20560 6933 20600
rect 6891 20551 6933 20560
rect 8523 20600 8565 20609
rect 8523 20560 8524 20600
rect 8564 20560 8565 20600
rect 8523 20551 8565 20560
rect 11395 20600 11453 20601
rect 11395 20560 11404 20600
rect 11444 20560 11453 20600
rect 11395 20559 11453 20560
rect 12259 20600 12317 20601
rect 12259 20560 12268 20600
rect 12308 20560 12317 20600
rect 12259 20559 12317 20560
rect 15139 20600 15197 20601
rect 15139 20560 15148 20600
rect 15188 20560 15197 20600
rect 15139 20559 15197 20560
rect 17739 20600 17781 20609
rect 17739 20560 17740 20600
rect 17780 20560 17781 20600
rect 17739 20551 17781 20560
rect 18019 20600 18077 20601
rect 18019 20560 18028 20600
rect 18068 20560 18077 20600
rect 18019 20559 18077 20560
rect 1152 20432 20452 20456
rect 1152 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20452 20432
rect 1152 20368 20452 20392
rect 8803 20264 8861 20265
rect 8803 20224 8812 20264
rect 8852 20224 8861 20264
rect 8803 20223 8861 20224
rect 9379 20264 9437 20265
rect 9379 20224 9388 20264
rect 9428 20224 9437 20264
rect 9379 20223 9437 20224
rect 11499 20264 11541 20273
rect 11499 20224 11500 20264
rect 11540 20224 11541 20264
rect 11499 20215 11541 20224
rect 13227 20264 13269 20273
rect 13227 20224 13228 20264
rect 13268 20224 13269 20264
rect 13227 20215 13269 20224
rect 14955 20264 14997 20273
rect 14955 20224 14956 20264
rect 14996 20224 14997 20264
rect 14955 20215 14997 20224
rect 18891 20264 18933 20273
rect 18891 20224 18892 20264
rect 18932 20224 18933 20264
rect 18891 20215 18933 20224
rect 2667 20180 2709 20189
rect 2667 20140 2668 20180
rect 2708 20140 2709 20180
rect 2667 20131 2709 20140
rect 6315 20180 6357 20189
rect 6315 20140 6316 20180
rect 6356 20140 6357 20180
rect 6315 20131 6357 20140
rect 7275 20180 7317 20189
rect 7275 20140 7276 20180
rect 7316 20140 7317 20180
rect 7275 20131 7317 20140
rect 11115 20180 11157 20189
rect 11115 20140 11116 20180
rect 11156 20140 11157 20180
rect 11115 20131 11157 20140
rect 1219 20096 1277 20097
rect 1219 20056 1228 20096
rect 1268 20056 1277 20096
rect 1219 20055 1277 20056
rect 2467 20096 2525 20097
rect 2467 20056 2476 20096
rect 2516 20056 2525 20096
rect 2467 20055 2525 20056
rect 2851 20096 2909 20097
rect 2851 20056 2860 20096
rect 2900 20056 2909 20096
rect 2851 20055 2909 20056
rect 4099 20096 4157 20097
rect 4099 20056 4108 20096
rect 4148 20056 4157 20096
rect 4099 20055 4157 20056
rect 4587 20096 4629 20105
rect 4587 20056 4588 20096
rect 4628 20056 4629 20096
rect 4587 20047 4629 20056
rect 4683 20096 4725 20105
rect 4683 20056 4684 20096
rect 4724 20056 4725 20096
rect 4683 20047 4725 20056
rect 5163 20096 5205 20105
rect 5163 20056 5164 20096
rect 5204 20056 5205 20096
rect 5163 20047 5205 20056
rect 5635 20096 5693 20097
rect 5635 20056 5644 20096
rect 5684 20056 5693 20096
rect 5635 20055 5693 20056
rect 6123 20091 6165 20100
rect 6123 20051 6124 20091
rect 6164 20051 6165 20091
rect 7171 20096 7229 20097
rect 7171 20056 7180 20096
rect 7220 20056 7229 20096
rect 7171 20055 7229 20056
rect 7851 20096 7893 20105
rect 7851 20056 7852 20096
rect 7892 20056 7893 20096
rect 6123 20042 6165 20051
rect 7851 20047 7893 20056
rect 8043 20096 8085 20105
rect 8043 20056 8044 20096
rect 8084 20056 8085 20096
rect 8043 20047 8085 20056
rect 8139 20096 8181 20105
rect 8139 20056 8140 20096
rect 8180 20056 8181 20096
rect 8139 20047 8181 20056
rect 8323 20096 8381 20097
rect 8323 20056 8332 20096
rect 8372 20056 8381 20096
rect 8323 20055 8381 20056
rect 8419 20096 8477 20097
rect 8419 20056 8428 20096
rect 8468 20056 8477 20096
rect 8715 20096 8757 20105
rect 8419 20055 8477 20056
rect 8571 20081 8613 20090
rect 8571 20041 8572 20081
rect 8612 20041 8613 20081
rect 8715 20056 8716 20096
rect 8756 20056 8757 20096
rect 9099 20096 9141 20105
rect 8715 20047 8757 20056
rect 8872 20081 8914 20090
rect 8571 20032 8613 20041
rect 8872 20041 8873 20081
rect 8913 20041 8914 20081
rect 9099 20056 9100 20096
rect 9140 20056 9141 20096
rect 9099 20047 9141 20056
rect 9195 20096 9237 20105
rect 9195 20056 9196 20096
rect 9236 20056 9237 20096
rect 9195 20047 9237 20056
rect 9667 20096 9725 20097
rect 9667 20056 9676 20096
rect 9716 20056 9725 20096
rect 9667 20055 9725 20056
rect 10915 20096 10973 20097
rect 10915 20056 10924 20096
rect 10964 20056 10973 20096
rect 10915 20055 10973 20056
rect 11307 20096 11349 20105
rect 11307 20056 11308 20096
rect 11348 20056 11349 20096
rect 11307 20047 11349 20056
rect 11403 20096 11445 20105
rect 11403 20056 11404 20096
rect 11444 20056 11445 20096
rect 11403 20047 11445 20056
rect 11595 20096 11637 20105
rect 11595 20056 11596 20096
rect 11636 20056 11637 20096
rect 11595 20047 11637 20056
rect 11779 20096 11837 20097
rect 11779 20056 11788 20096
rect 11828 20056 11837 20096
rect 11779 20055 11837 20056
rect 13027 20096 13085 20097
rect 13027 20056 13036 20096
rect 13076 20056 13085 20096
rect 13027 20055 13085 20056
rect 13507 20096 13565 20097
rect 13507 20056 13516 20096
rect 13556 20056 13565 20096
rect 13507 20055 13565 20056
rect 14755 20096 14813 20097
rect 14755 20056 14764 20096
rect 14804 20056 14813 20096
rect 14755 20055 14813 20056
rect 15811 20096 15869 20097
rect 15811 20056 15820 20096
rect 15860 20056 15869 20096
rect 15811 20055 15869 20056
rect 17059 20096 17117 20097
rect 17059 20056 17068 20096
rect 17108 20056 17117 20096
rect 17059 20055 17117 20056
rect 17443 20096 17501 20097
rect 17443 20056 17452 20096
rect 17492 20056 17501 20096
rect 17443 20055 17501 20056
rect 18691 20096 18749 20097
rect 18691 20056 18700 20096
rect 18740 20056 18749 20096
rect 18691 20055 18749 20056
rect 19166 20096 19224 20097
rect 19166 20056 19175 20096
rect 19215 20056 19224 20096
rect 19166 20055 19224 20056
rect 19275 20096 19317 20105
rect 19275 20056 19276 20096
rect 19316 20056 19317 20096
rect 19275 20047 19317 20056
rect 19371 20096 19413 20105
rect 19371 20056 19372 20096
rect 19412 20056 19413 20096
rect 19371 20047 19413 20056
rect 19555 20096 19613 20097
rect 19555 20056 19564 20096
rect 19604 20056 19613 20096
rect 19555 20055 19613 20056
rect 19651 20096 19709 20097
rect 19651 20056 19660 20096
rect 19700 20056 19709 20096
rect 19651 20055 19709 20056
rect 19851 20096 19893 20105
rect 19851 20056 19852 20096
rect 19892 20056 19893 20096
rect 19851 20047 19893 20056
rect 19947 20096 19989 20105
rect 19947 20056 19948 20096
rect 19988 20056 19989 20096
rect 19947 20047 19989 20056
rect 20043 20096 20085 20105
rect 20043 20056 20044 20096
rect 20084 20056 20085 20096
rect 20043 20047 20085 20056
rect 20139 20091 20181 20100
rect 20139 20051 20140 20091
rect 20180 20051 20181 20091
rect 20139 20042 20181 20051
rect 8872 20032 8914 20041
rect 5067 20012 5109 20021
rect 5067 19972 5068 20012
rect 5108 19972 5109 20012
rect 5067 19963 5109 19972
rect 4299 19928 4341 19937
rect 4299 19888 4300 19928
rect 4340 19888 4341 19928
rect 4299 19879 4341 19888
rect 8131 19928 8189 19929
rect 8131 19888 8140 19928
rect 8180 19888 8189 19928
rect 8131 19887 8189 19888
rect 17259 19928 17301 19937
rect 17259 19888 17260 19928
rect 17300 19888 17301 19928
rect 17259 19879 17301 19888
rect 19659 19844 19701 19853
rect 19659 19804 19660 19844
rect 19700 19804 19701 19844
rect 19659 19795 19701 19804
rect 1152 19676 20352 19700
rect 1152 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 20352 19676
rect 1152 19612 20352 19636
rect 2667 19508 2709 19517
rect 2667 19468 2668 19508
rect 2708 19468 2709 19508
rect 2667 19459 2709 19468
rect 4491 19508 4533 19517
rect 4491 19468 4492 19508
rect 4532 19468 4533 19508
rect 4491 19459 4533 19468
rect 6219 19508 6261 19517
rect 6219 19468 6220 19508
rect 6260 19468 6261 19508
rect 6219 19459 6261 19468
rect 8235 19508 8277 19517
rect 8235 19468 8236 19508
rect 8276 19468 8277 19508
rect 8235 19459 8277 19468
rect 10251 19508 10293 19517
rect 10251 19468 10252 19508
rect 10292 19468 10293 19508
rect 10251 19459 10293 19468
rect 13131 19508 13173 19517
rect 13131 19468 13132 19508
rect 13172 19468 13173 19508
rect 13131 19459 13173 19468
rect 17259 19508 17301 19517
rect 17259 19468 17260 19508
rect 17300 19468 17301 19508
rect 17259 19459 17301 19468
rect 17547 19424 17589 19433
rect 17547 19384 17548 19424
rect 17588 19384 17589 19424
rect 17547 19375 17589 19384
rect 19747 19424 19805 19425
rect 19747 19384 19756 19424
rect 19796 19384 19805 19424
rect 19747 19383 19805 19384
rect 10051 19298 10109 19299
rect 10051 19258 10060 19298
rect 10100 19258 10109 19298
rect 11080 19271 11122 19280
rect 10051 19257 10109 19258
rect 1219 19256 1277 19257
rect 1219 19216 1228 19256
rect 1268 19216 1277 19256
rect 1219 19215 1277 19216
rect 2467 19256 2525 19257
rect 2467 19216 2476 19256
rect 2516 19216 2525 19256
rect 2467 19215 2525 19216
rect 3043 19256 3101 19257
rect 3043 19216 3052 19256
rect 3092 19216 3101 19256
rect 3043 19215 3101 19216
rect 4291 19256 4349 19257
rect 4291 19216 4300 19256
rect 4340 19216 4349 19256
rect 4291 19215 4349 19216
rect 4771 19256 4829 19257
rect 4771 19216 4780 19256
rect 4820 19216 4829 19256
rect 4771 19215 4829 19216
rect 6019 19256 6077 19257
rect 6019 19216 6028 19256
rect 6068 19216 6077 19256
rect 6019 19215 6077 19216
rect 6787 19256 6845 19257
rect 6787 19216 6796 19256
rect 6836 19216 6845 19256
rect 6787 19215 6845 19216
rect 8035 19256 8093 19257
rect 8035 19216 8044 19256
rect 8084 19216 8093 19256
rect 8035 19215 8093 19216
rect 8803 19256 8861 19257
rect 8803 19216 8812 19256
rect 8852 19216 8861 19256
rect 8803 19215 8861 19216
rect 10531 19256 10589 19257
rect 10531 19216 10540 19256
rect 10580 19216 10589 19256
rect 10531 19215 10589 19216
rect 10627 19256 10685 19257
rect 10627 19216 10636 19256
rect 10676 19216 10685 19256
rect 10627 19215 10685 19216
rect 10827 19256 10869 19265
rect 10827 19216 10828 19256
rect 10868 19216 10869 19256
rect 10827 19207 10869 19216
rect 10923 19256 10965 19265
rect 10923 19216 10924 19256
rect 10964 19216 10965 19256
rect 11080 19231 11081 19271
rect 11121 19231 11122 19271
rect 11080 19222 11122 19231
rect 11683 19256 11741 19257
rect 10923 19207 10965 19216
rect 11683 19216 11692 19256
rect 11732 19216 11741 19256
rect 11683 19215 11741 19216
rect 12931 19256 12989 19257
rect 12931 19216 12940 19256
rect 12980 19216 12989 19256
rect 12931 19215 12989 19216
rect 13315 19256 13373 19257
rect 13315 19216 13324 19256
rect 13364 19216 13373 19256
rect 13315 19215 13373 19216
rect 13411 19256 13469 19257
rect 13411 19216 13420 19256
rect 13460 19216 13469 19256
rect 13411 19215 13469 19216
rect 13611 19256 13653 19265
rect 13611 19216 13612 19256
rect 13652 19216 13653 19256
rect 13611 19207 13653 19216
rect 13707 19256 13749 19265
rect 13707 19216 13708 19256
rect 13748 19216 13749 19256
rect 13707 19207 13749 19216
rect 13800 19256 13858 19257
rect 13800 19216 13809 19256
rect 13849 19216 13858 19256
rect 13800 19215 13858 19216
rect 14091 19256 14133 19265
rect 14091 19216 14092 19256
rect 14132 19216 14133 19256
rect 14091 19207 14133 19216
rect 14187 19256 14229 19265
rect 14187 19216 14188 19256
rect 14228 19216 14229 19256
rect 14187 19207 14229 19216
rect 15811 19256 15869 19257
rect 15811 19216 15820 19256
rect 15860 19216 15869 19256
rect 15811 19215 15869 19216
rect 17059 19256 17117 19257
rect 17059 19216 17068 19256
rect 17108 19216 17117 19256
rect 17059 19215 17117 19216
rect 17827 19256 17885 19257
rect 17827 19216 17836 19256
rect 17876 19216 17885 19256
rect 17827 19215 17885 19216
rect 19075 19256 19133 19257
rect 19075 19216 19084 19256
rect 19124 19216 19133 19256
rect 19075 19215 19133 19216
rect 19659 19256 19701 19265
rect 19659 19216 19660 19256
rect 19700 19216 19701 19256
rect 19659 19207 19701 19216
rect 19755 19256 19797 19265
rect 19755 19216 19756 19256
rect 19796 19216 19797 19256
rect 19755 19207 19797 19216
rect 19947 19256 19989 19265
rect 19947 19216 19948 19256
rect 19988 19216 19989 19256
rect 19947 19207 19989 19216
rect 19275 19172 19317 19181
rect 19275 19132 19276 19172
rect 19316 19132 19317 19172
rect 19275 19123 19317 19132
rect 10723 19088 10781 19089
rect 10723 19048 10732 19088
rect 10772 19048 10781 19088
rect 10723 19047 10781 19048
rect 13131 19088 13173 19097
rect 13131 19048 13132 19088
rect 13172 19048 13173 19088
rect 13131 19039 13173 19048
rect 13699 19088 13757 19089
rect 13699 19048 13708 19088
rect 13748 19048 13757 19088
rect 13699 19047 13757 19048
rect 14371 19088 14429 19089
rect 14371 19048 14380 19088
rect 14420 19048 14429 19088
rect 14371 19047 14429 19048
rect 17259 19088 17301 19097
rect 17259 19048 17260 19088
rect 17300 19048 17301 19088
rect 17259 19039 17301 19048
rect 17635 19088 17693 19089
rect 17635 19048 17644 19088
rect 17684 19048 17693 19088
rect 17635 19047 17693 19048
rect 1152 18920 20452 18944
rect 1152 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20452 18920
rect 1152 18856 20452 18880
rect 19363 18794 19421 18795
rect 2667 18752 2709 18761
rect 2667 18712 2668 18752
rect 2708 18712 2709 18752
rect 2667 18703 2709 18712
rect 6115 18752 6173 18753
rect 6115 18712 6124 18752
rect 6164 18712 6173 18752
rect 6115 18711 6173 18712
rect 8235 18752 8277 18761
rect 8235 18712 8236 18752
rect 8276 18712 8277 18752
rect 8235 18703 8277 18712
rect 10819 18752 10877 18753
rect 10819 18712 10828 18752
rect 10868 18712 10877 18752
rect 10819 18711 10877 18712
rect 14667 18752 14709 18761
rect 19363 18754 19372 18794
rect 19412 18754 19421 18794
rect 19363 18753 19421 18754
rect 14667 18712 14668 18752
rect 14708 18712 14709 18752
rect 14667 18703 14709 18712
rect 16963 18752 17021 18753
rect 16963 18712 16972 18752
rect 17012 18712 17021 18752
rect 16963 18711 17021 18712
rect 20235 18752 20277 18761
rect 20235 18712 20236 18752
rect 20276 18712 20277 18752
rect 20235 18703 20277 18712
rect 5067 18668 5109 18677
rect 5067 18628 5068 18668
rect 5108 18628 5109 18668
rect 5067 18619 5109 18628
rect 10155 18668 10197 18677
rect 10155 18628 10156 18668
rect 10196 18628 10197 18668
rect 10155 18619 10197 18628
rect 16683 18668 16725 18677
rect 16683 18628 16684 18668
rect 16724 18628 16725 18668
rect 16683 18619 16725 18628
rect 18891 18668 18933 18677
rect 18891 18628 18892 18668
rect 18932 18628 18933 18668
rect 18891 18619 18933 18628
rect 1219 18584 1277 18585
rect 1219 18544 1228 18584
rect 1268 18544 1277 18584
rect 1219 18543 1277 18544
rect 2467 18584 2525 18585
rect 2467 18544 2476 18584
rect 2516 18544 2525 18584
rect 2467 18543 2525 18544
rect 3331 18584 3389 18585
rect 3331 18544 3340 18584
rect 3380 18544 3389 18584
rect 3331 18543 3389 18544
rect 4579 18584 4637 18585
rect 4579 18544 4588 18584
rect 4628 18544 4637 18584
rect 4579 18543 4637 18544
rect 4971 18584 5013 18593
rect 4971 18544 4972 18584
rect 5012 18544 5013 18584
rect 4971 18535 5013 18544
rect 5163 18584 5205 18593
rect 5163 18544 5164 18584
rect 5204 18544 5205 18584
rect 5163 18535 5205 18544
rect 5355 18584 5397 18593
rect 5355 18544 5356 18584
rect 5396 18544 5397 18584
rect 5355 18535 5397 18544
rect 5643 18584 5685 18593
rect 5643 18544 5644 18584
rect 5684 18544 5685 18584
rect 5643 18535 5685 18544
rect 5835 18584 5877 18593
rect 5835 18544 5836 18584
rect 5876 18544 5877 18584
rect 5835 18535 5877 18544
rect 5931 18584 5973 18593
rect 5931 18544 5932 18584
rect 5972 18544 5973 18584
rect 5931 18535 5973 18544
rect 6307 18584 6365 18585
rect 6307 18544 6316 18584
rect 6356 18544 6365 18584
rect 6307 18543 6365 18544
rect 6500 18583 6542 18592
rect 6500 18543 6501 18583
rect 6541 18543 6542 18583
rect 6787 18584 6845 18585
rect 6787 18544 6796 18584
rect 6836 18544 6845 18584
rect 6787 18543 6845 18544
rect 8035 18584 8093 18585
rect 8035 18544 8044 18584
rect 8084 18544 8093 18584
rect 8035 18543 8093 18544
rect 8707 18584 8765 18585
rect 8707 18544 8716 18584
rect 8756 18544 8765 18584
rect 8707 18543 8765 18544
rect 9955 18584 10013 18585
rect 9955 18544 9964 18584
rect 10004 18544 10013 18584
rect 9955 18543 10013 18544
rect 10539 18584 10581 18593
rect 10539 18544 10540 18584
rect 10580 18544 10581 18584
rect 6500 18534 6542 18543
rect 10539 18535 10581 18544
rect 10635 18584 10677 18593
rect 10635 18544 10636 18584
rect 10676 18544 10677 18584
rect 10635 18535 10677 18544
rect 11395 18584 11453 18585
rect 11395 18544 11404 18584
rect 11444 18544 11453 18584
rect 11395 18543 11453 18544
rect 12643 18584 12701 18585
rect 12643 18544 12652 18584
rect 12692 18544 12701 18584
rect 12643 18543 12701 18544
rect 13219 18584 13277 18585
rect 13219 18544 13228 18584
rect 13268 18544 13277 18584
rect 13219 18543 13277 18544
rect 14467 18584 14525 18585
rect 14467 18544 14476 18584
rect 14516 18544 14525 18584
rect 14467 18543 14525 18544
rect 14955 18584 14997 18593
rect 14955 18544 14956 18584
rect 14996 18544 14997 18584
rect 14955 18535 14997 18544
rect 15051 18584 15093 18593
rect 15051 18544 15052 18584
rect 15092 18544 15093 18584
rect 15051 18535 15093 18544
rect 15531 18584 15573 18593
rect 15531 18544 15532 18584
rect 15572 18544 15573 18584
rect 15531 18535 15573 18544
rect 16003 18584 16061 18585
rect 16003 18544 16012 18584
rect 16052 18544 16061 18584
rect 17163 18584 17205 18593
rect 16003 18543 16061 18544
rect 16491 18570 16533 18579
rect 16491 18530 16492 18570
rect 16532 18530 16533 18570
rect 17163 18544 17164 18584
rect 17204 18544 17205 18584
rect 17163 18535 17205 18544
rect 17259 18584 17301 18593
rect 17259 18544 17260 18584
rect 17300 18544 17301 18584
rect 17259 18535 17301 18544
rect 18691 18584 18749 18585
rect 18691 18544 18700 18584
rect 18740 18544 18749 18584
rect 18691 18543 18749 18544
rect 19083 18584 19125 18593
rect 19083 18544 19084 18584
rect 19124 18544 19125 18584
rect 17443 18542 17501 18543
rect 16491 18521 16533 18530
rect 15435 18500 15477 18509
rect 17443 18502 17452 18542
rect 17492 18502 17501 18542
rect 19083 18535 19125 18544
rect 19179 18584 19221 18593
rect 19179 18544 19180 18584
rect 19220 18544 19221 18584
rect 19179 18535 19221 18544
rect 19563 18584 19605 18593
rect 19563 18544 19564 18584
rect 19604 18544 19605 18584
rect 19563 18535 19605 18544
rect 19659 18584 19701 18593
rect 19659 18544 19660 18584
rect 19700 18544 19701 18584
rect 19659 18535 19701 18544
rect 19851 18584 19893 18593
rect 19851 18544 19852 18584
rect 19892 18544 19893 18584
rect 19851 18535 19893 18544
rect 17443 18501 17501 18502
rect 15435 18460 15436 18500
rect 15476 18460 15477 18500
rect 15435 18451 15477 18460
rect 20035 18500 20093 18501
rect 20035 18460 20044 18500
rect 20084 18460 20093 18500
rect 20035 18459 20093 18460
rect 3051 18416 3093 18425
rect 3051 18376 3052 18416
rect 3092 18376 3093 18416
rect 3051 18367 3093 18376
rect 5643 18416 5685 18425
rect 5643 18376 5644 18416
rect 5684 18376 5685 18416
rect 5643 18367 5685 18376
rect 19555 18416 19613 18417
rect 19555 18376 19564 18416
rect 19604 18376 19613 18416
rect 19555 18375 19613 18376
rect 4779 18332 4821 18341
rect 4779 18292 4780 18332
rect 4820 18292 4821 18332
rect 4779 18283 4821 18292
rect 6411 18332 6453 18341
rect 6411 18292 6412 18332
rect 6452 18292 6453 18332
rect 6411 18283 6453 18292
rect 12843 18332 12885 18341
rect 12843 18292 12844 18332
rect 12884 18292 12885 18332
rect 12843 18283 12885 18292
rect 1152 18164 20352 18188
rect 1152 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 20352 18164
rect 1152 18100 20352 18124
rect 2091 17996 2133 18005
rect 2091 17956 2092 17996
rect 2132 17956 2133 17996
rect 2091 17947 2133 17956
rect 16779 17996 16821 18005
rect 16779 17956 16780 17996
rect 16820 17956 16821 17996
rect 16779 17947 16821 17956
rect 17163 17996 17205 18005
rect 17163 17956 17164 17996
rect 17204 17956 17205 17996
rect 17163 17947 17205 17956
rect 18795 17996 18837 18005
rect 18795 17956 18796 17996
rect 18836 17956 18837 17996
rect 18795 17947 18837 17956
rect 10435 17912 10493 17913
rect 10435 17872 10444 17912
rect 10484 17872 10493 17912
rect 10435 17871 10493 17872
rect 12843 17912 12885 17921
rect 12843 17872 12844 17912
rect 12884 17872 12885 17912
rect 12843 17863 12885 17872
rect 13795 17912 13853 17913
rect 13795 17872 13804 17912
rect 13844 17872 13853 17912
rect 13795 17871 13853 17872
rect 2859 17828 2901 17837
rect 2859 17788 2860 17828
rect 2900 17788 2901 17828
rect 2859 17779 2901 17788
rect 2955 17828 2997 17837
rect 2955 17788 2956 17828
rect 2996 17788 2997 17828
rect 2955 17779 2997 17788
rect 16195 17828 16253 17829
rect 16195 17788 16204 17828
rect 16244 17788 16253 17828
rect 16195 17787 16253 17788
rect 16579 17828 16637 17829
rect 16579 17788 16588 17828
rect 16628 17788 16637 17828
rect 16579 17787 16637 17788
rect 16963 17828 17021 17829
rect 16963 17788 16972 17828
rect 17012 17788 17021 17828
rect 16963 17787 17021 17788
rect 12643 17786 12701 17787
rect 1899 17757 1941 17766
rect 8619 17758 8661 17767
rect 1795 17744 1853 17745
rect 1795 17704 1804 17744
rect 1844 17704 1853 17744
rect 1899 17717 1900 17757
rect 1940 17717 1941 17757
rect 1899 17708 1941 17717
rect 2083 17744 2141 17745
rect 1795 17703 1853 17704
rect 2083 17704 2092 17744
rect 2132 17704 2141 17744
rect 2083 17703 2141 17704
rect 2379 17744 2421 17753
rect 2379 17704 2380 17744
rect 2420 17704 2421 17744
rect 2379 17695 2421 17704
rect 2475 17744 2517 17753
rect 3915 17749 3957 17758
rect 2475 17704 2476 17744
rect 2516 17704 2517 17744
rect 2475 17695 2517 17704
rect 3427 17744 3485 17745
rect 3427 17704 3436 17744
rect 3476 17704 3485 17744
rect 3427 17703 3485 17704
rect 3915 17709 3916 17749
rect 3956 17709 3957 17749
rect 3915 17700 3957 17709
rect 4395 17744 4437 17753
rect 4395 17704 4396 17744
rect 4436 17704 4437 17744
rect 4395 17695 4437 17704
rect 4587 17744 4629 17753
rect 4587 17704 4588 17744
rect 4628 17704 4629 17744
rect 4587 17695 4629 17704
rect 4683 17744 4725 17753
rect 4683 17704 4684 17744
rect 4724 17704 4725 17744
rect 4683 17695 4725 17704
rect 5067 17744 5109 17753
rect 5067 17704 5068 17744
rect 5108 17704 5109 17744
rect 5067 17695 5109 17704
rect 5163 17744 5205 17753
rect 5163 17704 5164 17744
rect 5204 17704 5205 17744
rect 5163 17695 5205 17704
rect 5347 17744 5405 17745
rect 5347 17704 5356 17744
rect 5396 17704 5405 17744
rect 5347 17703 5405 17704
rect 6595 17744 6653 17745
rect 6595 17704 6604 17744
rect 6644 17704 6653 17744
rect 6595 17703 6653 17704
rect 7083 17744 7125 17753
rect 7083 17704 7084 17744
rect 7124 17704 7125 17744
rect 7083 17695 7125 17704
rect 7179 17744 7221 17753
rect 7179 17704 7180 17744
rect 7220 17704 7221 17744
rect 7179 17695 7221 17704
rect 7563 17744 7605 17753
rect 7563 17704 7564 17744
rect 7604 17704 7605 17744
rect 7563 17695 7605 17704
rect 7659 17744 7701 17753
rect 7659 17704 7660 17744
rect 7700 17704 7701 17744
rect 7659 17695 7701 17704
rect 8131 17744 8189 17745
rect 8131 17704 8140 17744
rect 8180 17704 8189 17744
rect 8619 17718 8620 17758
rect 8660 17718 8661 17758
rect 8619 17709 8661 17718
rect 9195 17749 9237 17758
rect 9195 17709 9196 17749
rect 9236 17709 9237 17749
rect 8131 17703 8189 17704
rect 9195 17700 9237 17709
rect 9387 17744 9429 17753
rect 9387 17704 9388 17744
rect 9428 17704 9429 17744
rect 9387 17695 9429 17704
rect 9483 17744 9525 17753
rect 9483 17704 9484 17744
rect 9524 17704 9525 17744
rect 9483 17695 9525 17704
rect 9675 17744 9717 17753
rect 9675 17704 9676 17744
rect 9716 17704 9717 17744
rect 9675 17695 9717 17704
rect 9771 17744 9813 17753
rect 9771 17704 9772 17744
rect 9812 17704 9813 17744
rect 9771 17695 9813 17704
rect 10155 17744 10197 17753
rect 10155 17704 10156 17744
rect 10196 17704 10197 17744
rect 10155 17695 10197 17704
rect 10347 17744 10389 17753
rect 10347 17704 10348 17744
rect 10388 17704 10389 17744
rect 10347 17695 10389 17704
rect 10443 17744 10485 17753
rect 10443 17704 10444 17744
rect 10484 17704 10485 17744
rect 10443 17695 10485 17704
rect 10627 17744 10685 17745
rect 10627 17704 10636 17744
rect 10676 17704 10685 17744
rect 10627 17703 10685 17704
rect 10723 17744 10781 17745
rect 10723 17704 10732 17744
rect 10772 17704 10781 17744
rect 10723 17703 10781 17704
rect 10923 17744 10965 17753
rect 10923 17704 10924 17744
rect 10964 17704 10965 17744
rect 10923 17695 10965 17704
rect 11019 17744 11061 17753
rect 12643 17746 12652 17786
rect 12692 17746 12701 17786
rect 13323 17759 13365 17768
rect 12643 17745 12701 17746
rect 13075 17755 13133 17756
rect 11019 17704 11020 17744
rect 11060 17704 11061 17744
rect 11019 17695 11061 17704
rect 11112 17744 11170 17745
rect 11112 17704 11121 17744
rect 11161 17704 11170 17744
rect 11112 17703 11170 17704
rect 11395 17744 11453 17745
rect 11395 17704 11404 17744
rect 11444 17704 11453 17744
rect 13075 17715 13084 17755
rect 13124 17715 13133 17755
rect 13075 17714 13133 17715
rect 13227 17744 13269 17753
rect 11395 17703 11453 17704
rect 13227 17704 13228 17744
rect 13268 17704 13269 17744
rect 13323 17719 13324 17759
rect 13364 17719 13365 17759
rect 13323 17710 13365 17719
rect 13507 17744 13565 17745
rect 13227 17695 13269 17704
rect 13507 17704 13516 17744
rect 13556 17704 13565 17744
rect 13507 17703 13565 17704
rect 13603 17744 13661 17745
rect 13603 17704 13612 17744
rect 13652 17704 13661 17744
rect 13603 17703 13661 17704
rect 13803 17744 13845 17753
rect 13803 17704 13804 17744
rect 13844 17704 13845 17744
rect 13803 17695 13845 17704
rect 13899 17744 13941 17753
rect 13899 17704 13900 17744
rect 13940 17704 13941 17744
rect 13899 17695 13941 17704
rect 14091 17744 14133 17753
rect 14091 17704 14092 17744
rect 14132 17704 14133 17744
rect 14091 17695 14133 17704
rect 14275 17744 14333 17745
rect 14275 17704 14284 17744
rect 14324 17704 14333 17744
rect 14275 17703 14333 17704
rect 15523 17744 15581 17745
rect 15523 17704 15532 17744
rect 15572 17704 15581 17744
rect 15523 17703 15581 17704
rect 17347 17744 17405 17745
rect 17347 17704 17356 17744
rect 17396 17704 17405 17744
rect 17347 17703 17405 17704
rect 18595 17744 18653 17745
rect 18595 17704 18604 17744
rect 18644 17704 18653 17744
rect 18595 17703 18653 17704
rect 19070 17744 19128 17745
rect 19070 17704 19079 17744
rect 19119 17704 19128 17744
rect 19070 17703 19128 17704
rect 19179 17744 19221 17753
rect 19179 17704 19180 17744
rect 19220 17704 19221 17744
rect 19179 17695 19221 17704
rect 19275 17744 19317 17753
rect 19275 17704 19276 17744
rect 19316 17704 19317 17744
rect 19275 17695 19317 17704
rect 19459 17744 19517 17745
rect 19459 17704 19468 17744
rect 19508 17704 19517 17744
rect 19459 17703 19517 17704
rect 19555 17744 19613 17745
rect 19555 17704 19564 17744
rect 19604 17704 19613 17744
rect 19555 17703 19613 17704
rect 19755 17744 19797 17753
rect 19755 17704 19756 17744
rect 19796 17704 19797 17744
rect 19755 17695 19797 17704
rect 19851 17744 19893 17753
rect 19851 17704 19852 17744
rect 19892 17704 19893 17744
rect 19851 17695 19893 17704
rect 4107 17660 4149 17669
rect 4107 17620 4108 17660
rect 4148 17620 4149 17660
rect 4107 17611 4149 17620
rect 6795 17660 6837 17669
rect 6795 17620 6796 17660
rect 6836 17620 6837 17660
rect 6795 17611 6837 17620
rect 9291 17660 9333 17669
rect 9291 17620 9292 17660
rect 9332 17620 9333 17660
rect 9291 17611 9333 17620
rect 4491 17576 4533 17585
rect 4491 17536 4492 17576
rect 4532 17536 4533 17576
rect 4491 17527 4533 17536
rect 4867 17576 4925 17577
rect 4867 17536 4876 17576
rect 4916 17536 4925 17576
rect 9955 17576 10013 17577
rect 4867 17535 4925 17536
rect 8811 17534 8853 17543
rect 9955 17536 9964 17576
rect 10004 17536 10013 17576
rect 9955 17535 10013 17536
rect 11107 17576 11165 17577
rect 11107 17536 11116 17576
rect 11156 17536 11165 17576
rect 11107 17535 11165 17536
rect 13123 17576 13181 17577
rect 13123 17536 13132 17576
rect 13172 17536 13181 17576
rect 13123 17535 13181 17536
rect 15723 17576 15765 17585
rect 15723 17536 15724 17576
rect 15764 17536 15765 17576
rect 8811 17494 8812 17534
rect 8852 17494 8853 17534
rect 15723 17527 15765 17536
rect 16395 17576 16437 17585
rect 16395 17536 16396 17576
rect 16436 17536 16437 17576
rect 16395 17527 16437 17536
rect 19075 17576 19133 17577
rect 19075 17536 19084 17576
rect 19124 17536 19133 17576
rect 19075 17535 19133 17536
rect 20035 17576 20093 17577
rect 20035 17536 20044 17576
rect 20084 17536 20093 17576
rect 20035 17535 20093 17536
rect 8811 17485 8853 17494
rect 1152 17408 20452 17432
rect 1152 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20452 17408
rect 1152 17344 20452 17368
rect 3523 17240 3581 17241
rect 3523 17200 3532 17240
rect 3572 17200 3581 17240
rect 3523 17199 3581 17200
rect 3915 17240 3957 17249
rect 3915 17200 3916 17240
rect 3956 17200 3957 17240
rect 3915 17191 3957 17200
rect 9483 17240 9525 17249
rect 9483 17200 9484 17240
rect 9524 17200 9525 17240
rect 9483 17191 9525 17200
rect 16587 17240 16629 17249
rect 16587 17200 16588 17240
rect 16628 17200 16629 17240
rect 16587 17191 16629 17200
rect 17163 17240 17205 17249
rect 17163 17200 17164 17240
rect 17204 17200 17205 17240
rect 17163 17191 17205 17200
rect 19083 17240 19125 17249
rect 19083 17200 19084 17240
rect 19124 17200 19125 17240
rect 19083 17191 19125 17200
rect 19851 17240 19893 17249
rect 19851 17200 19852 17240
rect 19892 17200 19893 17240
rect 19851 17191 19893 17200
rect 20235 17240 20277 17249
rect 20235 17200 20236 17240
rect 20276 17200 20277 17240
rect 20235 17191 20277 17200
rect 7275 17156 7317 17165
rect 7275 17116 7276 17156
rect 7316 17116 7317 17156
rect 7275 17107 7317 17116
rect 9291 17156 9333 17165
rect 9291 17116 9292 17156
rect 9332 17116 9333 17156
rect 9291 17107 9333 17116
rect 12747 17156 12789 17165
rect 12747 17116 12748 17156
rect 12788 17116 12789 17156
rect 12747 17107 12789 17116
rect 14763 17156 14805 17165
rect 14763 17116 14764 17156
rect 14804 17116 14805 17156
rect 14763 17107 14805 17116
rect 13131 17092 13173 17101
rect 1219 17072 1277 17073
rect 1219 17032 1228 17072
rect 1268 17032 1277 17072
rect 1219 17031 1277 17032
rect 2467 17072 2525 17073
rect 2467 17032 2476 17072
rect 2516 17032 2525 17072
rect 2467 17031 2525 17032
rect 2947 17072 3005 17073
rect 2947 17032 2956 17072
rect 2996 17032 3005 17072
rect 2947 17031 3005 17032
rect 3230 17072 3288 17073
rect 3230 17032 3239 17072
rect 3279 17032 3288 17072
rect 3230 17031 3288 17032
rect 3339 17072 3381 17081
rect 3339 17032 3340 17072
rect 3380 17032 3381 17072
rect 3339 17023 3381 17032
rect 3435 17072 3477 17081
rect 3435 17032 3436 17072
rect 3476 17032 3477 17072
rect 3435 17023 3477 17032
rect 3619 17072 3677 17073
rect 3619 17032 3628 17072
rect 3668 17032 3677 17072
rect 3619 17031 3677 17032
rect 3715 17072 3773 17073
rect 3715 17032 3724 17072
rect 3764 17032 3773 17072
rect 3715 17031 3773 17032
rect 4099 17072 4157 17073
rect 4099 17032 4108 17072
rect 4148 17032 4157 17072
rect 4099 17031 4157 17032
rect 5347 17072 5405 17073
rect 5347 17032 5356 17072
rect 5396 17032 5405 17072
rect 5347 17031 5405 17032
rect 5827 17072 5885 17073
rect 5827 17032 5836 17072
rect 5876 17032 5885 17072
rect 5827 17031 5885 17032
rect 7075 17072 7133 17073
rect 7075 17032 7084 17072
rect 7124 17032 7133 17072
rect 7075 17031 7133 17032
rect 7563 17072 7605 17081
rect 7563 17032 7564 17072
rect 7604 17032 7605 17072
rect 7563 17023 7605 17032
rect 7659 17072 7701 17081
rect 7659 17032 7660 17072
rect 7700 17032 7701 17072
rect 7659 17023 7701 17032
rect 8611 17072 8669 17073
rect 8611 17032 8620 17072
rect 8660 17032 8669 17072
rect 9667 17072 9725 17073
rect 8611 17031 8669 17032
rect 9099 17058 9141 17067
rect 9099 17018 9100 17058
rect 9140 17018 9141 17058
rect 9667 17032 9676 17072
rect 9716 17032 9725 17072
rect 9667 17031 9725 17032
rect 10915 17072 10973 17073
rect 10915 17032 10924 17072
rect 10964 17032 10973 17072
rect 10915 17031 10973 17032
rect 11299 17072 11357 17073
rect 11299 17032 11308 17072
rect 11348 17032 11357 17072
rect 11299 17031 11357 17032
rect 12547 17072 12605 17073
rect 12547 17032 12556 17072
rect 12596 17032 12605 17072
rect 12547 17031 12605 17032
rect 13035 17072 13077 17081
rect 13035 17032 13036 17072
rect 13076 17032 13077 17072
rect 13131 17052 13132 17092
rect 13172 17052 13173 17092
rect 13131 17043 13173 17052
rect 14083 17072 14141 17073
rect 13035 17023 13077 17032
rect 14083 17032 14092 17072
rect 14132 17032 14141 17072
rect 15139 17072 15197 17073
rect 14083 17031 14141 17032
rect 14619 17030 14661 17039
rect 15139 17032 15148 17072
rect 15188 17032 15197 17072
rect 15139 17031 15197 17032
rect 16387 17072 16445 17073
rect 16387 17032 16396 17072
rect 16436 17032 16445 17072
rect 16387 17031 16445 17032
rect 17635 17072 17693 17073
rect 17635 17032 17644 17072
rect 17684 17032 17693 17072
rect 17635 17031 17693 17032
rect 18883 17072 18941 17073
rect 18883 17032 18892 17072
rect 18932 17032 18941 17072
rect 18883 17031 18941 17032
rect 9099 17009 9141 17018
rect 8043 16988 8085 16997
rect 8043 16948 8044 16988
rect 8084 16948 8085 16988
rect 8043 16939 8085 16948
rect 8139 16988 8181 16997
rect 8139 16948 8140 16988
rect 8180 16948 8181 16988
rect 8139 16939 8181 16948
rect 13515 16988 13557 16997
rect 13515 16948 13516 16988
rect 13556 16948 13557 16988
rect 13515 16939 13557 16948
rect 13611 16988 13653 16997
rect 13611 16948 13612 16988
rect 13652 16948 13653 16988
rect 14619 16990 14620 17030
rect 14660 16990 14661 17030
rect 14619 16981 14661 16990
rect 16963 16988 17021 16989
rect 13611 16939 13653 16948
rect 16963 16948 16972 16988
rect 17012 16948 17021 16988
rect 16963 16947 17021 16948
rect 19267 16988 19325 16989
rect 19267 16948 19276 16988
rect 19316 16948 19325 16988
rect 19267 16947 19325 16948
rect 19651 16988 19709 16989
rect 19651 16948 19660 16988
rect 19700 16948 19709 16988
rect 19651 16947 19709 16948
rect 20035 16988 20093 16989
rect 20035 16948 20044 16988
rect 20084 16948 20093 16988
rect 20035 16947 20093 16948
rect 2667 16904 2709 16913
rect 2667 16864 2668 16904
rect 2708 16864 2709 16904
rect 2667 16855 2709 16864
rect 2859 16904 2901 16913
rect 2859 16864 2860 16904
rect 2900 16864 2901 16904
rect 2859 16855 2901 16864
rect 19467 16820 19509 16829
rect 19467 16780 19468 16820
rect 19508 16780 19509 16820
rect 19467 16771 19509 16780
rect 1152 16652 20352 16676
rect 1152 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 20352 16652
rect 1152 16588 20352 16612
rect 5251 16484 5309 16485
rect 5251 16444 5260 16484
rect 5300 16444 5309 16484
rect 5251 16443 5309 16444
rect 9099 16484 9141 16493
rect 9099 16444 9100 16484
rect 9140 16444 9141 16484
rect 9099 16435 9141 16444
rect 9387 16484 9429 16493
rect 9387 16444 9388 16484
rect 9428 16444 9429 16484
rect 9387 16435 9429 16444
rect 14859 16484 14901 16493
rect 14859 16444 14860 16484
rect 14900 16444 14901 16484
rect 14859 16435 14901 16444
rect 15435 16400 15477 16409
rect 15435 16360 15436 16400
rect 15476 16360 15477 16400
rect 15435 16351 15477 16360
rect 17451 16400 17493 16409
rect 17451 16360 17452 16400
rect 17492 16360 17493 16400
rect 17451 16351 17493 16360
rect 17835 16400 17877 16409
rect 17835 16360 17836 16400
rect 17876 16360 17877 16400
rect 17835 16351 17877 16360
rect 15235 16316 15293 16317
rect 15235 16276 15244 16316
rect 15284 16276 15293 16316
rect 15235 16275 15293 16276
rect 17251 16316 17309 16317
rect 17251 16276 17260 16316
rect 17300 16276 17309 16316
rect 17251 16275 17309 16276
rect 17635 16316 17693 16317
rect 17635 16276 17644 16316
rect 17684 16276 17693 16316
rect 17635 16275 17693 16276
rect 2275 16232 2333 16233
rect 2275 16192 2284 16232
rect 2324 16192 2333 16232
rect 2275 16191 2333 16192
rect 3523 16232 3581 16233
rect 3523 16192 3532 16232
rect 3572 16192 3581 16232
rect 3523 16191 3581 16192
rect 4107 16232 4149 16241
rect 4107 16192 4108 16232
rect 4148 16192 4149 16232
rect 4107 16183 4149 16192
rect 4203 16232 4245 16241
rect 4203 16192 4204 16232
rect 4244 16192 4245 16232
rect 4203 16183 4245 16192
rect 4579 16232 4637 16233
rect 4579 16192 4588 16232
rect 4628 16192 4637 16232
rect 4579 16191 4637 16192
rect 4875 16232 4917 16241
rect 4875 16192 4876 16232
rect 4916 16192 4917 16232
rect 4875 16183 4917 16192
rect 5539 16232 5597 16233
rect 5539 16192 5548 16232
rect 5588 16192 5597 16232
rect 5539 16191 5597 16192
rect 6787 16232 6845 16233
rect 6787 16192 6796 16232
rect 6836 16192 6845 16232
rect 6787 16191 6845 16192
rect 7651 16232 7709 16233
rect 7651 16192 7660 16232
rect 7700 16192 7709 16232
rect 7651 16191 7709 16192
rect 8899 16232 8957 16233
rect 8899 16192 8908 16232
rect 8948 16192 8957 16232
rect 8899 16191 8957 16192
rect 9571 16232 9629 16233
rect 9571 16192 9580 16232
rect 9620 16192 9629 16232
rect 9571 16191 9629 16192
rect 10819 16232 10877 16233
rect 10819 16192 10828 16232
rect 10868 16192 10877 16232
rect 10819 16191 10877 16192
rect 12843 16232 12885 16241
rect 12843 16192 12844 16232
rect 12884 16192 12885 16232
rect 12843 16183 12885 16192
rect 12939 16232 12981 16241
rect 12939 16192 12940 16232
rect 12980 16192 12981 16232
rect 12939 16183 12981 16192
rect 13411 16232 13469 16233
rect 13411 16192 13420 16232
rect 13460 16192 13469 16232
rect 13411 16191 13469 16192
rect 14659 16232 14717 16233
rect 14659 16192 14668 16232
rect 14708 16192 14717 16232
rect 14659 16191 14717 16192
rect 15619 16232 15677 16233
rect 15619 16192 15628 16232
rect 15668 16192 15677 16232
rect 15619 16191 15677 16192
rect 16867 16232 16925 16233
rect 16867 16192 16876 16232
rect 16916 16192 16925 16232
rect 16867 16191 16925 16192
rect 18027 16232 18069 16241
rect 18027 16192 18028 16232
rect 18068 16192 18069 16232
rect 18027 16183 18069 16192
rect 18219 16232 18261 16241
rect 18219 16192 18220 16232
rect 18260 16192 18261 16232
rect 18219 16183 18261 16192
rect 18514 16237 18556 16246
rect 18514 16197 18515 16237
rect 18555 16197 18556 16237
rect 18514 16188 18556 16197
rect 18699 16232 18741 16241
rect 18699 16192 18700 16232
rect 18740 16192 18741 16232
rect 18699 16183 18741 16192
rect 18795 16232 18837 16241
rect 18795 16192 18796 16232
rect 18836 16192 18837 16232
rect 18795 16183 18837 16192
rect 18979 16232 19037 16233
rect 18979 16192 18988 16232
rect 19028 16192 19037 16232
rect 18979 16191 19037 16192
rect 19075 16232 19133 16233
rect 19075 16192 19084 16232
rect 19124 16192 19133 16232
rect 19075 16191 19133 16192
rect 19275 16232 19317 16241
rect 19275 16192 19276 16232
rect 19316 16192 19317 16232
rect 19275 16183 19317 16192
rect 19371 16232 19413 16241
rect 19371 16192 19372 16232
rect 19412 16192 19413 16232
rect 19371 16183 19413 16192
rect 19518 16232 19576 16233
rect 19518 16192 19527 16232
rect 19567 16192 19576 16232
rect 19518 16191 19576 16192
rect 19755 16232 19797 16241
rect 19755 16192 19756 16232
rect 19796 16192 19797 16232
rect 19755 16183 19797 16192
rect 19851 16232 19893 16241
rect 19851 16192 19852 16232
rect 19892 16192 19893 16232
rect 19851 16183 19893 16192
rect 3723 16148 3765 16157
rect 3723 16108 3724 16148
rect 3764 16108 3765 16148
rect 3723 16099 3765 16108
rect 4971 16148 5013 16157
rect 4971 16108 4972 16148
rect 5012 16108 5013 16148
rect 4971 16099 5013 16108
rect 3907 16064 3965 16065
rect 3907 16024 3916 16064
rect 3956 16024 3965 16064
rect 3907 16023 3965 16024
rect 6987 16064 7029 16073
rect 6987 16024 6988 16064
rect 7028 16024 7029 16064
rect 6987 16015 7029 16024
rect 13123 16064 13181 16065
rect 13123 16024 13132 16064
rect 13172 16024 13181 16064
rect 13123 16023 13181 16024
rect 17067 16064 17109 16073
rect 17067 16024 17068 16064
rect 17108 16024 17109 16064
rect 17067 16015 17109 16024
rect 18123 16064 18165 16073
rect 18123 16024 18124 16064
rect 18164 16024 18165 16064
rect 18123 16015 18165 16024
rect 18603 16064 18645 16073
rect 18603 16024 18604 16064
rect 18644 16024 18645 16064
rect 18603 16015 18645 16024
rect 19171 16064 19229 16065
rect 19171 16024 19180 16064
rect 19220 16024 19229 16064
rect 19171 16023 19229 16024
rect 20035 16064 20093 16065
rect 20035 16024 20044 16064
rect 20084 16024 20093 16064
rect 20035 16023 20093 16024
rect 1152 15896 20452 15920
rect 1152 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20452 15896
rect 1152 15832 20452 15856
rect 3051 15728 3093 15737
rect 3051 15688 3052 15728
rect 3092 15688 3093 15728
rect 3051 15679 3093 15688
rect 3627 15728 3669 15737
rect 3627 15688 3628 15728
rect 3668 15688 3669 15728
rect 3627 15679 3669 15688
rect 16971 15728 17013 15737
rect 16971 15688 16972 15728
rect 17012 15688 17013 15728
rect 16971 15679 17013 15688
rect 19083 15728 19125 15737
rect 19083 15688 19084 15728
rect 19124 15688 19125 15728
rect 19083 15679 19125 15688
rect 19467 15728 19509 15737
rect 19467 15688 19468 15728
rect 19508 15688 19509 15728
rect 19467 15679 19509 15688
rect 19851 15728 19893 15737
rect 19851 15688 19852 15728
rect 19892 15688 19893 15728
rect 19851 15679 19893 15688
rect 20235 15728 20277 15737
rect 20235 15688 20236 15728
rect 20276 15688 20277 15728
rect 20235 15679 20277 15688
rect 5643 15644 5685 15653
rect 5643 15604 5644 15644
rect 5684 15604 5685 15644
rect 5643 15595 5685 15604
rect 8619 15644 8661 15653
rect 8619 15604 8620 15644
rect 8660 15604 8661 15644
rect 8619 15595 8661 15604
rect 1603 15560 1661 15561
rect 1603 15520 1612 15560
rect 1652 15520 1661 15560
rect 1603 15519 1661 15520
rect 2851 15560 2909 15561
rect 2851 15520 2860 15560
rect 2900 15520 2909 15560
rect 2851 15519 2909 15520
rect 3915 15560 3957 15569
rect 3915 15520 3916 15560
rect 3956 15520 3957 15560
rect 3915 15511 3957 15520
rect 4011 15560 4053 15569
rect 4011 15520 4012 15560
rect 4052 15520 4053 15560
rect 4011 15511 4053 15520
rect 4491 15560 4533 15569
rect 4491 15520 4492 15560
rect 4532 15520 4533 15560
rect 4491 15511 4533 15520
rect 4963 15560 5021 15561
rect 4963 15520 4972 15560
rect 5012 15520 5021 15560
rect 6891 15560 6933 15569
rect 4963 15519 5021 15520
rect 5451 15546 5493 15555
rect 5451 15506 5452 15546
rect 5492 15506 5493 15546
rect 6891 15520 6892 15560
rect 6932 15520 6933 15560
rect 6891 15511 6933 15520
rect 6987 15560 7029 15569
rect 6987 15520 6988 15560
rect 7028 15520 7029 15560
rect 6987 15511 7029 15520
rect 7939 15560 7997 15561
rect 7939 15520 7948 15560
rect 7988 15520 7997 15560
rect 8899 15560 8957 15561
rect 7939 15519 7997 15520
rect 8427 15546 8469 15555
rect 5451 15497 5493 15506
rect 8427 15506 8428 15546
rect 8468 15506 8469 15546
rect 8899 15520 8908 15560
rect 8948 15520 8957 15560
rect 8899 15519 8957 15520
rect 10147 15560 10205 15561
rect 10147 15520 10156 15560
rect 10196 15520 10205 15560
rect 10147 15519 10205 15520
rect 10531 15560 10589 15561
rect 10531 15520 10540 15560
rect 10580 15520 10589 15560
rect 10531 15519 10589 15520
rect 10731 15560 10773 15569
rect 10731 15520 10732 15560
rect 10772 15520 10773 15560
rect 10731 15511 10773 15520
rect 11587 15560 11645 15561
rect 11587 15520 11596 15560
rect 11636 15520 11645 15560
rect 11587 15519 11645 15520
rect 12835 15560 12893 15561
rect 12835 15520 12844 15560
rect 12884 15520 12893 15560
rect 12835 15519 12893 15520
rect 13699 15560 13757 15561
rect 13699 15520 13708 15560
rect 13748 15520 13757 15560
rect 13699 15519 13757 15520
rect 14947 15560 15005 15561
rect 14947 15520 14956 15560
rect 14996 15520 15005 15560
rect 14947 15519 15005 15520
rect 15523 15560 15581 15561
rect 15523 15520 15532 15560
rect 15572 15520 15581 15560
rect 15523 15519 15581 15520
rect 16771 15560 16829 15561
rect 16771 15520 16780 15560
rect 16820 15520 16829 15560
rect 16771 15519 16829 15520
rect 17155 15560 17213 15561
rect 17155 15520 17164 15560
rect 17204 15520 17213 15560
rect 17155 15519 17213 15520
rect 17259 15560 17301 15569
rect 17259 15520 17260 15560
rect 17300 15520 17301 15560
rect 17259 15511 17301 15520
rect 17451 15560 17493 15569
rect 17451 15520 17452 15560
rect 17492 15520 17493 15560
rect 17451 15511 17493 15520
rect 17635 15560 17693 15561
rect 17635 15520 17644 15560
rect 17684 15520 17693 15560
rect 17635 15519 17693 15520
rect 18883 15560 18941 15561
rect 18883 15520 18892 15560
rect 18932 15520 18941 15560
rect 18883 15519 18941 15520
rect 8427 15497 8469 15506
rect 3427 15476 3485 15477
rect 3427 15436 3436 15476
rect 3476 15436 3485 15476
rect 3427 15435 3485 15436
rect 4395 15476 4437 15485
rect 4395 15436 4396 15476
rect 4436 15436 4437 15476
rect 4395 15427 4437 15436
rect 7371 15476 7413 15485
rect 7371 15436 7372 15476
rect 7412 15436 7413 15476
rect 7371 15427 7413 15436
rect 7467 15476 7509 15485
rect 7467 15436 7468 15476
rect 7508 15436 7509 15476
rect 7467 15427 7509 15436
rect 19267 15476 19325 15477
rect 19267 15436 19276 15476
rect 19316 15436 19325 15476
rect 19267 15435 19325 15436
rect 19651 15476 19709 15477
rect 19651 15436 19660 15476
rect 19700 15436 19709 15476
rect 19651 15435 19709 15436
rect 20035 15476 20093 15477
rect 20035 15436 20044 15476
rect 20084 15436 20093 15476
rect 20035 15435 20093 15436
rect 13419 15392 13461 15401
rect 13419 15352 13420 15392
rect 13460 15352 13461 15392
rect 13419 15343 13461 15352
rect 10347 15308 10389 15317
rect 10347 15268 10348 15308
rect 10388 15268 10389 15308
rect 10347 15259 10389 15268
rect 10635 15308 10677 15317
rect 10635 15268 10636 15308
rect 10676 15268 10677 15308
rect 10635 15259 10677 15268
rect 13035 15308 13077 15317
rect 13035 15268 13036 15308
rect 13076 15268 13077 15308
rect 13035 15259 13077 15268
rect 15147 15308 15189 15317
rect 15147 15268 15148 15308
rect 15188 15268 15189 15308
rect 15147 15259 15189 15268
rect 17451 15308 17493 15317
rect 17451 15268 17452 15308
rect 17492 15268 17493 15308
rect 17451 15259 17493 15268
rect 1152 15140 20352 15164
rect 1152 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 20352 15140
rect 1152 15076 20352 15100
rect 2667 14972 2709 14981
rect 2667 14932 2668 14972
rect 2708 14932 2709 14972
rect 2667 14923 2709 14932
rect 5451 14972 5493 14981
rect 5451 14932 5452 14972
rect 5492 14932 5493 14972
rect 5451 14923 5493 14932
rect 8139 14972 8181 14981
rect 8139 14932 8140 14972
rect 8180 14932 8181 14972
rect 8139 14923 8181 14932
rect 17259 14972 17301 14981
rect 17259 14932 17260 14972
rect 17300 14932 17301 14972
rect 17259 14923 17301 14932
rect 19179 14972 19221 14981
rect 19179 14932 19180 14972
rect 19220 14932 19221 14972
rect 19179 14923 19221 14932
rect 20043 14972 20085 14981
rect 20043 14932 20044 14972
rect 20084 14932 20085 14972
rect 20043 14923 20085 14932
rect 3627 14888 3669 14897
rect 3627 14848 3628 14888
rect 3668 14848 3669 14888
rect 3627 14839 3669 14848
rect 9187 14888 9245 14889
rect 9187 14848 9196 14888
rect 9236 14848 9245 14888
rect 9187 14847 9245 14848
rect 9579 14888 9621 14897
rect 9579 14848 9580 14888
rect 9620 14848 9621 14888
rect 9579 14839 9621 14848
rect 19843 14804 19901 14805
rect 19843 14764 19852 14804
rect 19892 14764 19901 14804
rect 19843 14763 19901 14764
rect 1219 14720 1277 14721
rect 1219 14680 1228 14720
rect 1268 14680 1277 14720
rect 1219 14679 1277 14680
rect 2467 14720 2525 14721
rect 2467 14680 2476 14720
rect 2516 14680 2525 14720
rect 2467 14679 2525 14680
rect 3051 14720 3093 14729
rect 3051 14680 3052 14720
rect 3092 14680 3093 14720
rect 3051 14671 3093 14680
rect 3339 14720 3381 14729
rect 3339 14680 3340 14720
rect 3380 14680 3381 14720
rect 3339 14671 3381 14680
rect 3531 14720 3573 14729
rect 3531 14680 3532 14720
rect 3572 14680 3573 14720
rect 3531 14671 3573 14680
rect 3723 14720 3765 14729
rect 3723 14680 3724 14720
rect 3764 14680 3765 14720
rect 3723 14671 3765 14680
rect 3819 14720 3861 14729
rect 3819 14680 3820 14720
rect 3860 14680 3861 14720
rect 3819 14671 3861 14680
rect 4003 14720 4061 14721
rect 4003 14680 4012 14720
rect 4052 14680 4061 14720
rect 4003 14679 4061 14680
rect 5251 14720 5309 14721
rect 5251 14680 5260 14720
rect 5300 14680 5309 14720
rect 5251 14679 5309 14680
rect 5643 14720 5685 14729
rect 5643 14680 5644 14720
rect 5684 14680 5685 14720
rect 5643 14671 5685 14680
rect 5835 14720 5877 14729
rect 5835 14680 5836 14720
rect 5876 14680 5877 14720
rect 5835 14671 5877 14680
rect 5931 14720 5973 14729
rect 5931 14680 5932 14720
rect 5972 14680 5973 14720
rect 5931 14671 5973 14680
rect 6691 14720 6749 14721
rect 6691 14680 6700 14720
rect 6740 14680 6749 14720
rect 6691 14679 6749 14680
rect 7939 14720 7997 14721
rect 7939 14680 7948 14720
rect 7988 14680 7997 14720
rect 7939 14679 7997 14680
rect 8515 14720 8573 14721
rect 8515 14680 8524 14720
rect 8564 14680 8573 14720
rect 8515 14679 8573 14680
rect 8811 14720 8853 14729
rect 8811 14680 8812 14720
rect 8852 14680 8853 14720
rect 8811 14671 8853 14680
rect 9387 14720 9429 14729
rect 9387 14680 9388 14720
rect 9428 14680 9429 14720
rect 9387 14671 9429 14680
rect 9579 14720 9621 14729
rect 9579 14680 9580 14720
rect 9620 14680 9621 14720
rect 9579 14671 9621 14680
rect 9771 14720 9813 14729
rect 9771 14680 9772 14720
rect 9812 14680 9813 14720
rect 9771 14671 9813 14680
rect 10059 14720 10101 14729
rect 10059 14680 10060 14720
rect 10100 14680 10101 14720
rect 10059 14671 10101 14680
rect 10347 14720 10389 14729
rect 10347 14680 10348 14720
rect 10388 14680 10389 14720
rect 10347 14671 10389 14680
rect 10443 14720 10485 14729
rect 10443 14680 10444 14720
rect 10484 14680 10485 14720
rect 10443 14671 10485 14680
rect 10827 14720 10869 14729
rect 10827 14680 10828 14720
rect 10868 14680 10869 14720
rect 10827 14671 10869 14680
rect 10923 14720 10965 14729
rect 11883 14725 11925 14734
rect 15003 14729 15045 14738
rect 10923 14680 10924 14720
rect 10964 14680 10965 14720
rect 10923 14671 10965 14680
rect 11395 14720 11453 14721
rect 11395 14680 11404 14720
rect 11444 14680 11453 14720
rect 11395 14679 11453 14680
rect 11883 14685 11884 14725
rect 11924 14685 11925 14725
rect 11883 14676 11925 14685
rect 13419 14720 13461 14729
rect 13419 14680 13420 14720
rect 13460 14680 13461 14720
rect 13419 14671 13461 14680
rect 13515 14720 13557 14729
rect 13515 14680 13516 14720
rect 13556 14680 13557 14720
rect 13515 14671 13557 14680
rect 13899 14720 13941 14729
rect 13899 14680 13900 14720
rect 13940 14680 13941 14720
rect 13899 14671 13941 14680
rect 13995 14720 14037 14729
rect 13995 14680 13996 14720
rect 14036 14680 14037 14720
rect 13995 14671 14037 14680
rect 14467 14720 14525 14721
rect 14467 14680 14476 14720
rect 14516 14680 14525 14720
rect 15003 14689 15004 14729
rect 15044 14689 15045 14729
rect 15003 14680 15045 14689
rect 15523 14720 15581 14721
rect 15523 14680 15532 14720
rect 15572 14680 15581 14720
rect 14467 14679 14525 14680
rect 15523 14679 15581 14680
rect 16771 14720 16829 14721
rect 16771 14680 16780 14720
rect 16820 14680 16829 14720
rect 16771 14679 16829 14680
rect 16963 14720 17021 14721
rect 16963 14680 16972 14720
rect 17012 14680 17021 14720
rect 16963 14679 17021 14680
rect 17067 14720 17109 14729
rect 17067 14680 17068 14720
rect 17108 14680 17109 14720
rect 17067 14671 17109 14680
rect 17259 14720 17301 14729
rect 17259 14680 17260 14720
rect 17300 14680 17301 14720
rect 17259 14671 17301 14680
rect 17451 14720 17493 14729
rect 17451 14680 17452 14720
rect 17492 14680 17493 14720
rect 17451 14671 17493 14680
rect 17539 14720 17597 14721
rect 17539 14680 17548 14720
rect 17588 14680 17597 14720
rect 17539 14679 17597 14680
rect 17731 14720 17789 14721
rect 17731 14680 17740 14720
rect 17780 14680 17789 14720
rect 17731 14679 17789 14680
rect 18979 14720 19037 14721
rect 18979 14680 18988 14720
rect 19028 14680 19037 14720
rect 18979 14679 19037 14680
rect 19371 14720 19413 14729
rect 19371 14680 19372 14720
rect 19412 14680 19413 14720
rect 19371 14671 19413 14680
rect 19467 14720 19509 14729
rect 19467 14680 19468 14720
rect 19508 14680 19509 14720
rect 19467 14671 19509 14680
rect 19659 14720 19701 14729
rect 19659 14680 19660 14720
rect 19700 14680 19701 14720
rect 19659 14671 19701 14680
rect 3243 14636 3285 14645
rect 3243 14596 3244 14636
rect 3284 14596 3285 14636
rect 3243 14587 3285 14596
rect 8907 14636 8949 14645
rect 8907 14596 8908 14636
rect 8948 14596 8949 14636
rect 8907 14587 8949 14596
rect 12075 14636 12117 14645
rect 12075 14596 12076 14636
rect 12116 14596 12117 14636
rect 12075 14587 12117 14596
rect 15339 14636 15381 14645
rect 15339 14596 15340 14636
rect 15380 14596 15381 14636
rect 15339 14587 15381 14596
rect 5739 14552 5781 14561
rect 5739 14512 5740 14552
rect 5780 14512 5781 14552
rect 5739 14503 5781 14512
rect 9963 14552 10005 14561
rect 9963 14512 9964 14552
rect 10004 14512 10005 14552
rect 9963 14503 10005 14512
rect 15147 14552 15189 14561
rect 15147 14512 15148 14552
rect 15188 14512 15189 14552
rect 15147 14503 15189 14512
rect 19563 14552 19605 14561
rect 19563 14512 19564 14552
rect 19604 14512 19605 14552
rect 19563 14503 19605 14512
rect 1152 14384 20452 14408
rect 1152 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20452 14384
rect 1152 14320 20452 14344
rect 3147 14216 3189 14225
rect 3147 14176 3148 14216
rect 3188 14176 3189 14216
rect 3147 14167 3189 14176
rect 5347 14216 5405 14217
rect 5347 14176 5356 14216
rect 5396 14176 5405 14216
rect 5347 14175 5405 14176
rect 5827 14216 5885 14217
rect 5827 14176 5836 14216
rect 5876 14176 5885 14216
rect 5827 14175 5885 14176
rect 8043 14216 8085 14225
rect 8043 14176 8044 14216
rect 8084 14176 8085 14216
rect 8043 14167 8085 14176
rect 8235 14216 8277 14225
rect 8235 14176 8236 14216
rect 8276 14176 8277 14216
rect 8235 14167 8277 14176
rect 11403 14216 11445 14225
rect 11403 14176 11404 14216
rect 11444 14176 11445 14216
rect 11403 14167 11445 14176
rect 13035 14216 13077 14225
rect 13035 14176 13036 14216
rect 13076 14176 13077 14216
rect 13035 14167 13077 14176
rect 17547 14216 17589 14225
rect 17547 14176 17548 14216
rect 17588 14176 17589 14216
rect 17547 14167 17589 14176
rect 18019 14216 18077 14217
rect 18019 14176 18028 14216
rect 18068 14176 18077 14216
rect 18019 14175 18077 14176
rect 20235 14216 20277 14225
rect 20235 14176 20236 14216
rect 20276 14176 20277 14216
rect 20235 14167 20277 14176
rect 15147 14132 15189 14141
rect 15147 14092 15148 14132
rect 15188 14092 15189 14132
rect 15147 14083 15189 14092
rect 1699 14048 1757 14049
rect 1699 14008 1708 14048
rect 1748 14008 1757 14048
rect 1699 14007 1757 14008
rect 2947 14048 3005 14049
rect 2947 14008 2956 14048
rect 2996 14008 3005 14048
rect 2947 14007 3005 14008
rect 3531 14048 3573 14057
rect 3531 14008 3532 14048
rect 3572 14008 3573 14048
rect 3531 13999 3573 14008
rect 3627 14048 3669 14057
rect 3627 14008 3628 14048
rect 3668 14008 3669 14048
rect 3627 13999 3669 14008
rect 3723 14048 3765 14057
rect 3723 14008 3724 14048
rect 3764 14008 3765 14048
rect 3723 13999 3765 14008
rect 3819 14048 3861 14057
rect 3819 14008 3820 14048
rect 3860 14008 3861 14048
rect 3819 13999 3861 14008
rect 4003 14048 4061 14049
rect 4003 14008 4012 14048
rect 4052 14008 4061 14048
rect 4003 14007 4061 14008
rect 4395 14048 4437 14057
rect 4395 14008 4396 14048
rect 4436 14008 4437 14048
rect 4395 13999 4437 14008
rect 4867 14048 4925 14049
rect 4867 14008 4876 14048
rect 4916 14008 4925 14048
rect 4867 14007 4925 14008
rect 4963 14048 5021 14049
rect 4963 14008 4972 14048
rect 5012 14008 5021 14048
rect 4963 14007 5021 14008
rect 5163 14048 5205 14057
rect 5163 14008 5164 14048
rect 5204 14008 5205 14048
rect 5163 13999 5205 14008
rect 5259 14048 5301 14057
rect 5259 14008 5260 14048
rect 5300 14008 5301 14048
rect 6027 14048 6069 14057
rect 5259 13999 5301 14008
rect 5416 14033 5458 14042
rect 5416 13993 5417 14033
rect 5457 13993 5458 14033
rect 6027 14008 6028 14048
rect 6068 14008 6069 14048
rect 6027 13999 6069 14008
rect 6123 14048 6165 14057
rect 6123 14008 6124 14048
rect 6164 14008 6165 14048
rect 6123 13999 6165 14008
rect 6403 14048 6461 14049
rect 6403 14008 6412 14048
rect 6452 14008 6461 14048
rect 6403 14007 6461 14008
rect 6595 14048 6653 14049
rect 6595 14008 6604 14048
rect 6644 14008 6653 14048
rect 6595 14007 6653 14008
rect 7843 14048 7901 14049
rect 7843 14008 7852 14048
rect 7892 14008 7901 14048
rect 7843 14007 7901 14008
rect 8419 14048 8477 14049
rect 8419 14008 8428 14048
rect 8468 14008 8477 14048
rect 8419 14007 8477 14008
rect 9667 14048 9725 14049
rect 9667 14008 9676 14048
rect 9716 14008 9725 14048
rect 9667 14007 9725 14008
rect 9955 14048 10013 14049
rect 9955 14008 9964 14048
rect 10004 14008 10013 14048
rect 9955 14007 10013 14008
rect 11203 14048 11261 14049
rect 11203 14008 11212 14048
rect 11252 14008 11261 14048
rect 11203 14007 11261 14008
rect 11587 14048 11645 14049
rect 11587 14008 11596 14048
rect 11636 14008 11645 14048
rect 11587 14007 11645 14008
rect 12835 14048 12893 14049
rect 12835 14008 12844 14048
rect 12884 14008 12893 14048
rect 12835 14007 12893 14008
rect 13419 14048 13461 14057
rect 13419 14008 13420 14048
rect 13460 14008 13461 14048
rect 13419 13999 13461 14008
rect 13515 14048 13557 14057
rect 13515 14008 13516 14048
rect 13556 14008 13557 14048
rect 13515 13999 13557 14008
rect 14467 14048 14525 14049
rect 14467 14008 14476 14048
rect 14516 14008 14525 14048
rect 14467 14007 14525 14008
rect 14955 14043 14997 14052
rect 14955 14003 14956 14043
rect 14996 14003 14997 14043
rect 14955 13994 14997 14003
rect 15819 14048 15861 14057
rect 15819 14008 15820 14048
rect 15860 14008 15861 14048
rect 15819 13999 15861 14008
rect 15915 14048 15957 14057
rect 15915 14008 15916 14048
rect 15956 14008 15957 14048
rect 15915 13999 15957 14008
rect 16867 14048 16925 14049
rect 16867 14008 16876 14048
rect 16916 14008 16925 14048
rect 16867 14007 16925 14008
rect 17355 14043 17397 14052
rect 17355 14003 17356 14043
rect 17396 14003 17397 14043
rect 17355 13994 17397 14003
rect 17739 14048 17781 14057
rect 17739 14008 17740 14048
rect 17780 14008 17781 14048
rect 17739 13999 17781 14008
rect 17835 14048 17877 14057
rect 17835 14008 17836 14048
rect 17876 14008 17877 14048
rect 17835 13999 17877 14008
rect 18403 14048 18461 14049
rect 18403 14008 18412 14048
rect 18452 14008 18461 14048
rect 18403 14007 18461 14008
rect 19651 14048 19709 14049
rect 19651 14008 19660 14048
rect 19700 14008 19709 14048
rect 19651 14007 19709 14008
rect 5416 13984 5458 13993
rect 4107 13964 4149 13973
rect 4107 13924 4108 13964
rect 4148 13924 4149 13964
rect 4107 13915 4149 13924
rect 4299 13964 4341 13973
rect 4299 13924 4300 13964
rect 4340 13924 4341 13964
rect 4299 13915 4341 13924
rect 6315 13964 6357 13973
rect 6315 13924 6316 13964
rect 6356 13924 6357 13964
rect 6315 13915 6357 13924
rect 13899 13964 13941 13973
rect 13899 13924 13900 13964
rect 13940 13924 13941 13964
rect 13899 13915 13941 13924
rect 13995 13964 14037 13973
rect 13995 13924 13996 13964
rect 14036 13924 14037 13964
rect 13995 13915 14037 13924
rect 16299 13964 16341 13973
rect 16299 13924 16300 13964
rect 16340 13924 16341 13964
rect 16299 13915 16341 13924
rect 16395 13964 16437 13973
rect 16395 13924 16396 13964
rect 16436 13924 16437 13964
rect 16395 13915 16437 13924
rect 20035 13964 20093 13965
rect 20035 13924 20044 13964
rect 20084 13924 20093 13964
rect 20035 13923 20093 13924
rect 4203 13880 4245 13889
rect 4203 13840 4204 13880
rect 4244 13840 4245 13880
rect 4203 13831 4245 13840
rect 4683 13880 4725 13889
rect 4683 13840 4684 13880
rect 4724 13840 4725 13880
rect 4683 13831 4725 13840
rect 8043 13796 8085 13805
rect 8043 13756 8044 13796
rect 8084 13756 8085 13796
rect 8043 13747 8085 13756
rect 8235 13796 8277 13805
rect 8235 13756 8236 13796
rect 8276 13756 8277 13796
rect 8235 13747 8277 13756
rect 19851 13796 19893 13805
rect 19851 13756 19852 13796
rect 19892 13756 19893 13796
rect 19851 13747 19893 13756
rect 1152 13628 20352 13652
rect 1152 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 20352 13628
rect 1152 13564 20352 13588
rect 3147 13460 3189 13469
rect 3147 13420 3148 13460
rect 3188 13420 3189 13460
rect 3147 13411 3189 13420
rect 7179 13460 7221 13469
rect 7179 13420 7180 13460
rect 7220 13420 7221 13460
rect 7179 13411 7221 13420
rect 15907 13460 15965 13461
rect 15907 13420 15916 13460
rect 15956 13420 15965 13460
rect 15907 13419 15965 13420
rect 16867 13460 16925 13461
rect 16867 13420 16876 13460
rect 16916 13420 16925 13460
rect 16867 13419 16925 13420
rect 20235 13460 20277 13469
rect 20235 13420 20236 13460
rect 20276 13420 20277 13460
rect 20235 13411 20277 13420
rect 3619 13376 3677 13377
rect 3619 13336 3628 13376
rect 3668 13336 3677 13376
rect 3619 13335 3677 13336
rect 4683 13376 4725 13385
rect 4683 13336 4684 13376
rect 4724 13336 4725 13376
rect 4683 13327 4725 13336
rect 11595 13376 11637 13385
rect 11595 13336 11596 13376
rect 11636 13336 11637 13376
rect 11595 13327 11637 13336
rect 19075 13376 19133 13377
rect 19075 13336 19084 13376
rect 19124 13336 19133 13376
rect 19075 13335 19133 13336
rect 20035 13292 20093 13293
rect 20035 13252 20044 13292
rect 20084 13252 20093 13292
rect 20035 13251 20093 13252
rect 6699 13222 6741 13231
rect 1699 13208 1757 13209
rect 1699 13168 1708 13208
rect 1748 13168 1757 13208
rect 1699 13167 1757 13168
rect 2947 13208 3005 13209
rect 2947 13168 2956 13208
rect 2996 13168 3005 13208
rect 2947 13167 3005 13168
rect 3915 13208 3957 13217
rect 3915 13168 3916 13208
rect 3956 13168 3957 13208
rect 3915 13159 3957 13168
rect 4011 13208 4053 13217
rect 4011 13168 4012 13208
rect 4052 13168 4053 13208
rect 4011 13159 4053 13168
rect 4291 13208 4349 13209
rect 4291 13168 4300 13208
rect 4340 13168 4349 13208
rect 4291 13167 4349 13168
rect 5163 13208 5205 13217
rect 5163 13168 5164 13208
rect 5204 13168 5205 13208
rect 5163 13159 5205 13168
rect 5259 13208 5301 13217
rect 5259 13168 5260 13208
rect 5300 13168 5301 13208
rect 5259 13159 5301 13168
rect 5643 13208 5685 13217
rect 5643 13168 5644 13208
rect 5684 13168 5685 13208
rect 5643 13159 5685 13168
rect 5739 13208 5781 13217
rect 5739 13168 5740 13208
rect 5780 13168 5781 13208
rect 5739 13159 5781 13168
rect 6211 13208 6269 13209
rect 6211 13168 6220 13208
rect 6260 13168 6269 13208
rect 6699 13182 6700 13222
rect 6740 13182 6741 13222
rect 7563 13208 7605 13217
rect 6699 13173 6741 13182
rect 7075 13197 7133 13198
rect 6211 13167 6269 13168
rect 7075 13157 7084 13197
rect 7124 13157 7133 13197
rect 7563 13168 7564 13208
rect 7604 13168 7605 13208
rect 7563 13159 7605 13168
rect 7659 13208 7701 13217
rect 7659 13168 7660 13208
rect 7700 13168 7701 13208
rect 7659 13159 7701 13168
rect 7843 13208 7901 13209
rect 7843 13168 7852 13208
rect 7892 13168 7901 13208
rect 7843 13167 7901 13168
rect 7947 13208 7989 13217
rect 7947 13168 7948 13208
rect 7988 13168 7989 13208
rect 7947 13159 7989 13168
rect 8131 13208 8189 13209
rect 8131 13168 8140 13208
rect 8180 13168 8189 13208
rect 8131 13167 8189 13168
rect 8323 13208 8381 13209
rect 8323 13168 8332 13208
rect 8372 13168 8381 13208
rect 8323 13167 8381 13168
rect 9571 13208 9629 13209
rect 9571 13168 9580 13208
rect 9620 13168 9629 13208
rect 9571 13167 9629 13168
rect 9955 13208 10013 13209
rect 9955 13168 9964 13208
rect 10004 13168 10013 13208
rect 9955 13167 10013 13168
rect 11203 13208 11261 13209
rect 11203 13168 11212 13208
rect 11252 13168 11261 13208
rect 11203 13167 11261 13168
rect 12939 13208 12981 13217
rect 12939 13168 12940 13208
rect 12980 13168 12981 13208
rect 12939 13159 12981 13168
rect 13035 13208 13077 13217
rect 13035 13168 13036 13208
rect 13076 13168 13077 13208
rect 13035 13159 13077 13168
rect 13419 13208 13461 13217
rect 13419 13168 13420 13208
rect 13460 13168 13461 13208
rect 13419 13159 13461 13168
rect 13515 13208 13557 13217
rect 14475 13213 14517 13222
rect 13515 13168 13516 13208
rect 13556 13168 13557 13208
rect 13515 13159 13557 13168
rect 13987 13208 14045 13209
rect 13987 13168 13996 13208
rect 14036 13168 14045 13208
rect 13987 13167 14045 13168
rect 14475 13173 14476 13213
rect 14516 13173 14517 13213
rect 14475 13164 14517 13173
rect 15235 13208 15293 13209
rect 15235 13168 15244 13208
rect 15284 13168 15293 13208
rect 15235 13167 15293 13168
rect 15531 13208 15573 13217
rect 15531 13168 15532 13208
rect 15572 13168 15573 13208
rect 15531 13159 15573 13168
rect 15627 13208 15669 13217
rect 15627 13168 15628 13208
rect 15668 13168 15669 13208
rect 15627 13159 15669 13168
rect 16195 13208 16253 13209
rect 16195 13168 16204 13208
rect 16244 13168 16253 13208
rect 16195 13167 16253 13168
rect 16491 13208 16533 13217
rect 16491 13168 16492 13208
rect 16532 13168 16533 13208
rect 16491 13159 16533 13168
rect 16587 13208 16629 13217
rect 16587 13168 16588 13208
rect 16628 13168 16629 13208
rect 16587 13159 16629 13168
rect 17347 13208 17405 13209
rect 17347 13168 17356 13208
rect 17396 13168 17405 13208
rect 17347 13167 17405 13168
rect 18595 13208 18653 13209
rect 18595 13168 18604 13208
rect 18644 13168 18653 13208
rect 18595 13167 18653 13168
rect 19371 13208 19413 13217
rect 19371 13168 19372 13208
rect 19412 13168 19413 13208
rect 19371 13159 19413 13168
rect 19467 13208 19509 13217
rect 19467 13168 19468 13208
rect 19508 13168 19509 13208
rect 19467 13159 19509 13168
rect 19747 13208 19805 13209
rect 19747 13168 19756 13208
rect 19796 13168 19805 13208
rect 19747 13167 19805 13168
rect 7075 13156 7133 13157
rect 6891 13124 6933 13133
rect 6891 13084 6892 13124
rect 6932 13084 6933 13124
rect 6891 13075 6933 13084
rect 11403 13124 11445 13133
rect 11403 13084 11404 13124
rect 11444 13084 11445 13124
rect 11403 13075 11445 13084
rect 14667 13124 14709 13133
rect 14667 13084 14668 13124
rect 14708 13084 14709 13124
rect 14667 13075 14709 13084
rect 3147 13040 3189 13049
rect 3147 13000 3148 13040
rect 3188 13000 3189 13040
rect 3147 12991 3189 13000
rect 7363 13040 7421 13041
rect 7363 13000 7372 13040
rect 7412 13000 7421 13040
rect 7363 12999 7421 13000
rect 8139 13040 8181 13049
rect 8139 13000 8140 13040
rect 8180 13000 8181 13040
rect 8139 12991 8181 13000
rect 9771 13040 9813 13049
rect 9771 13000 9772 13040
rect 9812 13000 9813 13040
rect 9771 12991 9813 13000
rect 18795 13040 18837 13049
rect 18795 13000 18796 13040
rect 18836 13000 18837 13040
rect 18795 12991 18837 13000
rect 1152 12872 20452 12896
rect 1152 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20452 12872
rect 1152 12808 20452 12832
rect 10531 12704 10589 12705
rect 10531 12664 10540 12704
rect 10580 12664 10589 12704
rect 10531 12663 10589 12664
rect 14475 12704 14517 12713
rect 14475 12664 14476 12704
rect 14516 12664 14517 12704
rect 14475 12655 14517 12664
rect 17355 12704 17397 12713
rect 17355 12664 17356 12704
rect 17396 12664 17397 12704
rect 17355 12655 17397 12664
rect 17923 12704 17981 12705
rect 17923 12664 17932 12704
rect 17972 12664 17981 12704
rect 17923 12663 17981 12664
rect 3627 12620 3669 12629
rect 3627 12580 3628 12620
rect 3668 12580 3669 12620
rect 3627 12571 3669 12580
rect 4875 12620 4917 12629
rect 4875 12580 4876 12620
rect 4916 12580 4917 12620
rect 4875 12571 4917 12580
rect 6987 12620 7029 12629
rect 6987 12580 6988 12620
rect 7028 12580 7029 12620
rect 6987 12571 7029 12580
rect 9003 12620 9045 12629
rect 9003 12580 9004 12620
rect 9044 12580 9045 12620
rect 9003 12571 9045 12580
rect 12555 12620 12597 12629
rect 12555 12580 12556 12620
rect 12596 12580 12597 12620
rect 12555 12571 12597 12580
rect 15339 12620 15381 12629
rect 15339 12580 15340 12620
rect 15380 12580 15381 12620
rect 15339 12571 15381 12580
rect 20235 12620 20277 12629
rect 20235 12580 20236 12620
rect 20276 12580 20277 12620
rect 20235 12571 20277 12580
rect 1227 12536 1269 12545
rect 1227 12496 1228 12536
rect 1268 12496 1269 12536
rect 1227 12487 1269 12496
rect 1419 12536 1461 12545
rect 1419 12496 1420 12536
rect 1460 12496 1461 12536
rect 1419 12487 1461 12496
rect 1515 12536 1557 12545
rect 1515 12496 1516 12536
rect 1556 12496 1557 12536
rect 1515 12487 1557 12496
rect 1699 12536 1757 12537
rect 1699 12496 1708 12536
rect 1748 12496 1757 12536
rect 1699 12495 1757 12496
rect 2947 12536 3005 12537
rect 2947 12496 2956 12536
rect 2996 12496 3005 12536
rect 2947 12495 3005 12496
rect 3339 12536 3381 12545
rect 3339 12496 3340 12536
rect 3380 12496 3381 12536
rect 3339 12487 3381 12496
rect 3435 12536 3477 12545
rect 3435 12496 3436 12536
rect 3476 12496 3477 12536
rect 3435 12487 3477 12496
rect 3531 12536 3573 12545
rect 3531 12496 3532 12536
rect 3572 12496 3573 12536
rect 3531 12487 3573 12496
rect 3819 12536 3861 12545
rect 3819 12496 3820 12536
rect 3860 12496 3861 12536
rect 3819 12487 3861 12496
rect 3915 12536 3957 12545
rect 3915 12496 3916 12536
rect 3956 12496 3957 12536
rect 3915 12487 3957 12496
rect 4011 12536 4053 12545
rect 4011 12496 4012 12536
rect 4052 12496 4053 12536
rect 4011 12487 4053 12496
rect 4107 12536 4149 12545
rect 4107 12496 4108 12536
rect 4148 12496 4149 12536
rect 4107 12487 4149 12496
rect 4971 12536 5013 12545
rect 4971 12496 4972 12536
rect 5012 12496 5013 12536
rect 4971 12487 5013 12496
rect 5251 12536 5309 12537
rect 5251 12496 5260 12536
rect 5300 12496 5309 12536
rect 5251 12495 5309 12496
rect 5635 12536 5693 12537
rect 5635 12496 5644 12536
rect 5684 12496 5693 12536
rect 5635 12495 5693 12496
rect 5739 12536 5781 12545
rect 5739 12496 5740 12536
rect 5780 12496 5781 12536
rect 5739 12487 5781 12496
rect 5931 12536 5973 12545
rect 5931 12496 5932 12536
rect 5972 12496 5973 12536
rect 5931 12487 5973 12496
rect 6123 12536 6165 12545
rect 6123 12496 6124 12536
rect 6164 12496 6165 12536
rect 6123 12487 6165 12496
rect 6411 12536 6453 12545
rect 6411 12496 6412 12536
rect 6452 12496 6453 12536
rect 6411 12487 6453 12496
rect 7275 12536 7317 12545
rect 7275 12496 7276 12536
rect 7316 12496 7317 12536
rect 7275 12487 7317 12496
rect 7371 12536 7413 12545
rect 7371 12496 7372 12536
rect 7412 12496 7413 12536
rect 7371 12487 7413 12496
rect 7851 12536 7893 12545
rect 7851 12496 7852 12536
rect 7892 12496 7893 12536
rect 7851 12487 7893 12496
rect 8323 12536 8381 12537
rect 8323 12496 8332 12536
rect 8372 12496 8381 12536
rect 10251 12536 10293 12545
rect 8323 12495 8381 12496
rect 8811 12522 8853 12531
rect 8811 12482 8812 12522
rect 8852 12482 8853 12522
rect 10251 12496 10252 12536
rect 10292 12496 10293 12536
rect 10251 12487 10293 12496
rect 10347 12536 10389 12545
rect 10347 12496 10348 12536
rect 10388 12496 10389 12536
rect 10347 12487 10389 12496
rect 10827 12536 10869 12545
rect 10827 12496 10828 12536
rect 10868 12496 10869 12536
rect 10827 12487 10869 12496
rect 10923 12536 10965 12545
rect 10923 12496 10924 12536
rect 10964 12496 10965 12536
rect 10923 12487 10965 12496
rect 11403 12536 11445 12545
rect 11403 12496 11404 12536
rect 11444 12496 11445 12536
rect 11403 12487 11445 12496
rect 11875 12536 11933 12537
rect 11875 12496 11884 12536
rect 11924 12496 11933 12536
rect 13027 12536 13085 12537
rect 11875 12495 11933 12496
rect 12363 12522 12405 12531
rect 8811 12473 8853 12482
rect 12363 12482 12364 12522
rect 12404 12482 12405 12522
rect 13027 12496 13036 12536
rect 13076 12496 13085 12536
rect 13027 12495 13085 12496
rect 14275 12536 14333 12537
rect 14275 12496 14284 12536
rect 14324 12496 14333 12536
rect 14275 12495 14333 12496
rect 14851 12536 14909 12537
rect 14851 12496 14860 12536
rect 14900 12496 14909 12536
rect 14851 12495 14909 12496
rect 14955 12536 14997 12545
rect 14955 12496 14956 12536
rect 14996 12496 14997 12536
rect 14955 12487 14997 12496
rect 15147 12536 15189 12545
rect 15147 12496 15148 12536
rect 15188 12496 15189 12536
rect 16003 12536 16061 12537
rect 15147 12487 15189 12496
rect 15531 12522 15573 12531
rect 12363 12473 12405 12482
rect 15531 12482 15532 12522
rect 15572 12482 15573 12522
rect 16003 12496 16012 12536
rect 16052 12496 16061 12536
rect 16003 12495 16061 12496
rect 16491 12536 16533 12545
rect 16491 12496 16492 12536
rect 16532 12496 16533 12536
rect 16491 12487 16533 12496
rect 16971 12536 17013 12545
rect 16971 12496 16972 12536
rect 17012 12496 17013 12536
rect 16971 12487 17013 12496
rect 17067 12536 17109 12545
rect 17067 12496 17068 12536
rect 17108 12496 17109 12536
rect 17067 12487 17109 12496
rect 17643 12536 17685 12545
rect 17643 12496 17644 12536
rect 17684 12496 17685 12536
rect 17643 12487 17685 12496
rect 17739 12536 17781 12545
rect 17739 12496 17740 12536
rect 17780 12496 17781 12536
rect 17739 12487 17781 12496
rect 18507 12536 18549 12545
rect 18507 12496 18508 12536
rect 18548 12496 18549 12536
rect 18507 12487 18549 12496
rect 18603 12536 18645 12545
rect 18603 12496 18604 12536
rect 18644 12496 18645 12536
rect 18603 12487 18645 12496
rect 19555 12536 19613 12537
rect 19555 12496 19564 12536
rect 19604 12496 19613 12536
rect 19555 12495 19613 12496
rect 20043 12531 20085 12540
rect 20043 12491 20044 12531
rect 20084 12491 20085 12531
rect 20043 12482 20085 12491
rect 15531 12473 15573 12482
rect 7755 12452 7797 12461
rect 7755 12412 7756 12452
rect 7796 12412 7797 12452
rect 7755 12403 7797 12412
rect 11307 12452 11349 12461
rect 11307 12412 11308 12452
rect 11348 12412 11349 12452
rect 11307 12403 11349 12412
rect 16587 12452 16629 12461
rect 16587 12412 16588 12452
rect 16628 12412 16629 12452
rect 16587 12403 16629 12412
rect 18987 12452 19029 12461
rect 18987 12412 18988 12452
rect 19028 12412 19029 12452
rect 18987 12403 19029 12412
rect 19083 12452 19125 12461
rect 19083 12412 19084 12452
rect 19124 12412 19125 12452
rect 19083 12403 19125 12412
rect 1411 12368 1469 12369
rect 1411 12328 1420 12368
rect 1460 12328 1469 12368
rect 1411 12327 1469 12328
rect 4579 12368 4637 12369
rect 4579 12328 4588 12368
rect 4628 12328 4637 12368
rect 4579 12327 4637 12328
rect 5931 12368 5973 12377
rect 5931 12328 5932 12368
rect 5972 12328 5973 12368
rect 5931 12319 5973 12328
rect 6603 12368 6645 12377
rect 6603 12328 6604 12368
rect 6644 12328 6645 12368
rect 6603 12319 6645 12328
rect 9195 12368 9237 12377
rect 9195 12328 9196 12368
rect 9236 12328 9237 12368
rect 9195 12319 9237 12328
rect 15147 12368 15189 12377
rect 15147 12328 15148 12368
rect 15188 12328 15189 12368
rect 15147 12319 15189 12328
rect 3147 12284 3189 12293
rect 3147 12244 3148 12284
rect 3188 12244 3189 12284
rect 3147 12235 3189 12244
rect 6123 12284 6165 12293
rect 6123 12244 6124 12284
rect 6164 12244 6165 12284
rect 6123 12235 6165 12244
rect 1152 12116 20352 12140
rect 1152 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 20352 12116
rect 1152 12052 20352 12076
rect 3147 11948 3189 11957
rect 3147 11908 3148 11948
rect 3188 11908 3189 11948
rect 3147 11899 3189 11908
rect 6411 11948 6453 11957
rect 6411 11908 6412 11948
rect 6452 11908 6453 11948
rect 6411 11899 6453 11908
rect 6891 11948 6933 11957
rect 6891 11908 6892 11948
rect 6932 11908 6933 11948
rect 6891 11899 6933 11908
rect 9003 11948 9045 11957
rect 9003 11908 9004 11948
rect 9044 11908 9045 11948
rect 9003 11899 9045 11908
rect 10635 11948 10677 11957
rect 10635 11908 10636 11948
rect 10676 11908 10677 11948
rect 10635 11899 10677 11908
rect 12267 11948 12309 11957
rect 12267 11908 12268 11948
rect 12308 11908 12309 11948
rect 12267 11899 12309 11908
rect 17931 11948 17973 11957
rect 17931 11908 17932 11948
rect 17972 11908 17973 11948
rect 17931 11899 17973 11908
rect 20139 11948 20181 11957
rect 20139 11908 20140 11948
rect 20180 11908 20181 11948
rect 20139 11899 20181 11908
rect 3435 11864 3477 11873
rect 3435 11824 3436 11864
rect 3476 11824 3477 11864
rect 3435 11815 3477 11824
rect 3715 11864 3773 11865
rect 3715 11824 3724 11864
rect 3764 11824 3773 11864
rect 3715 11823 3773 11824
rect 4299 11864 4341 11873
rect 4299 11824 4300 11864
rect 4340 11824 4341 11864
rect 4299 11815 4341 11824
rect 4683 11864 4725 11873
rect 4683 11824 4684 11864
rect 4724 11824 4725 11864
rect 4683 11815 4725 11824
rect 1227 11696 1269 11705
rect 1227 11656 1228 11696
rect 1268 11656 1269 11696
rect 1227 11647 1269 11656
rect 1419 11696 1461 11705
rect 1419 11656 1420 11696
rect 1460 11656 1461 11696
rect 1419 11647 1461 11656
rect 1515 11696 1557 11705
rect 1515 11656 1516 11696
rect 1556 11656 1557 11696
rect 1515 11647 1557 11656
rect 1699 11696 1757 11697
rect 1699 11656 1708 11696
rect 1748 11656 1757 11696
rect 1699 11655 1757 11656
rect 2947 11696 3005 11697
rect 2947 11656 2956 11696
rect 2996 11656 3005 11696
rect 2947 11655 3005 11656
rect 3331 11696 3389 11697
rect 3331 11656 3340 11696
rect 3380 11656 3389 11696
rect 3331 11655 3389 11656
rect 3627 11696 3669 11705
rect 3627 11656 3628 11696
rect 3668 11656 3669 11696
rect 3627 11647 3669 11656
rect 3723 11696 3765 11705
rect 3723 11656 3724 11696
rect 3764 11656 3765 11696
rect 3723 11647 3765 11656
rect 3915 11696 3957 11705
rect 3915 11656 3916 11696
rect 3956 11656 3957 11696
rect 3915 11647 3957 11656
rect 4107 11696 4149 11705
rect 4107 11656 4108 11696
rect 4148 11656 4149 11696
rect 4107 11647 4149 11656
rect 4203 11696 4245 11705
rect 4203 11656 4204 11696
rect 4244 11656 4245 11696
rect 4203 11647 4245 11656
rect 4395 11696 4437 11705
rect 4395 11656 4396 11696
rect 4436 11656 4437 11696
rect 4395 11647 4437 11656
rect 4963 11696 5021 11697
rect 4963 11656 4972 11696
rect 5012 11656 5021 11696
rect 4963 11655 5021 11656
rect 6211 11696 6269 11697
rect 6211 11656 6220 11696
rect 6260 11656 6269 11696
rect 6211 11655 6269 11656
rect 6603 11696 6645 11705
rect 6603 11656 6604 11696
rect 6644 11656 6645 11696
rect 6603 11647 6645 11656
rect 6891 11696 6933 11705
rect 6891 11656 6892 11696
rect 6932 11656 6933 11696
rect 6891 11647 6933 11656
rect 7083 11696 7125 11705
rect 7083 11656 7084 11696
rect 7124 11656 7125 11696
rect 7083 11647 7125 11656
rect 7555 11696 7613 11697
rect 7555 11656 7564 11696
rect 7604 11656 7613 11696
rect 7555 11655 7613 11656
rect 8803 11696 8861 11697
rect 8803 11656 8812 11696
rect 8852 11656 8861 11696
rect 8803 11655 8861 11656
rect 10059 11696 10101 11705
rect 10059 11656 10060 11696
rect 10100 11656 10101 11696
rect 10059 11647 10101 11656
rect 10155 11696 10197 11705
rect 10155 11656 10156 11696
rect 10196 11656 10197 11696
rect 10155 11647 10197 11656
rect 10347 11696 10389 11705
rect 10347 11656 10348 11696
rect 10388 11656 10389 11696
rect 10347 11647 10389 11656
rect 10635 11696 10677 11705
rect 10635 11656 10636 11696
rect 10676 11656 10677 11696
rect 10635 11647 10677 11656
rect 10819 11696 10877 11697
rect 10819 11656 10828 11696
rect 10868 11656 10877 11696
rect 10819 11655 10877 11656
rect 12067 11696 12125 11697
rect 12067 11656 12076 11696
rect 12116 11656 12125 11696
rect 12067 11655 12125 11656
rect 13891 11696 13949 11697
rect 13891 11656 13900 11696
rect 13940 11656 13949 11696
rect 13891 11655 13949 11656
rect 15139 11696 15197 11697
rect 15139 11656 15148 11696
rect 15188 11656 15197 11696
rect 15139 11655 15197 11656
rect 15715 11696 15773 11697
rect 15715 11656 15724 11696
rect 15764 11656 15773 11696
rect 15715 11655 15773 11656
rect 16963 11696 17021 11697
rect 16963 11656 16972 11696
rect 17012 11656 17021 11696
rect 16963 11655 17021 11656
rect 17163 11696 17205 11705
rect 17163 11656 17164 11696
rect 17204 11656 17205 11696
rect 17163 11647 17205 11656
rect 17259 11696 17301 11705
rect 17259 11656 17260 11696
rect 17300 11656 17301 11696
rect 17259 11647 17301 11656
rect 17355 11696 17397 11705
rect 17355 11656 17356 11696
rect 17396 11656 17397 11696
rect 17355 11647 17397 11656
rect 17931 11696 17973 11705
rect 17931 11656 17932 11696
rect 17972 11656 17973 11696
rect 17931 11647 17973 11656
rect 18219 11696 18261 11705
rect 18219 11656 18220 11696
rect 18260 11656 18261 11696
rect 18219 11647 18261 11656
rect 18691 11696 18749 11697
rect 18691 11656 18700 11696
rect 18740 11656 18749 11696
rect 18691 11655 18749 11656
rect 19939 11696 19997 11697
rect 19939 11656 19948 11696
rect 19988 11656 19997 11696
rect 19939 11655 19997 11656
rect 9195 11612 9237 11621
rect 9195 11572 9196 11612
rect 9236 11572 9237 11612
rect 9195 11563 9237 11572
rect 15339 11612 15381 11621
rect 15339 11572 15340 11612
rect 15380 11572 15381 11612
rect 15339 11563 15381 11572
rect 1323 11528 1365 11537
rect 1323 11488 1324 11528
rect 1364 11488 1365 11528
rect 1323 11479 1365 11488
rect 6699 11528 6741 11537
rect 6699 11488 6700 11528
rect 6740 11488 6741 11528
rect 6699 11479 6741 11488
rect 9859 11528 9917 11529
rect 9859 11488 9868 11528
rect 9908 11488 9917 11528
rect 9859 11487 9917 11488
rect 15531 11528 15573 11537
rect 15531 11488 15532 11528
rect 15572 11488 15573 11528
rect 15531 11479 15573 11488
rect 17443 11528 17501 11529
rect 17443 11488 17452 11528
rect 17492 11488 17501 11528
rect 17443 11487 17501 11488
rect 1152 11360 20452 11384
rect 1152 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20452 11360
rect 1152 11296 20452 11320
rect 13035 11234 13077 11243
rect 2667 11192 2709 11201
rect 13035 11194 13036 11234
rect 13076 11194 13077 11234
rect 2667 11152 2668 11192
rect 2708 11152 2709 11192
rect 2667 11143 2709 11152
rect 4675 11192 4733 11193
rect 4675 11152 4684 11192
rect 4724 11152 4733 11192
rect 4675 11151 4733 11152
rect 6115 11192 6173 11193
rect 6115 11152 6124 11192
rect 6164 11152 6173 11192
rect 13035 11185 13077 11194
rect 16963 11192 17021 11193
rect 6115 11151 6173 11152
rect 16963 11152 16972 11192
rect 17012 11152 17021 11192
rect 16963 11151 17021 11152
rect 17731 11192 17789 11193
rect 17731 11152 17740 11192
rect 17780 11152 17789 11192
rect 17731 11151 17789 11152
rect 8619 11108 8661 11117
rect 8619 11068 8620 11108
rect 8660 11068 8661 11108
rect 8619 11059 8661 11068
rect 11019 11108 11061 11117
rect 11019 11068 11020 11108
rect 11060 11068 11061 11108
rect 11019 11059 11061 11068
rect 15051 11108 15093 11117
rect 15051 11068 15052 11108
rect 15092 11068 15093 11108
rect 15051 11059 15093 11068
rect 20139 11108 20181 11117
rect 20139 11068 20140 11108
rect 20180 11068 20181 11108
rect 20139 11059 20181 11068
rect 1219 11024 1277 11025
rect 1219 10984 1228 11024
rect 1268 10984 1277 11024
rect 1219 10983 1277 10984
rect 2467 11024 2525 11025
rect 2467 10984 2476 11024
rect 2516 10984 2525 11024
rect 2467 10983 2525 10984
rect 2851 11024 2909 11025
rect 2851 10984 2860 11024
rect 2900 10984 2909 11024
rect 2851 10983 2909 10984
rect 4099 11024 4157 11025
rect 4099 10984 4108 11024
rect 4148 10984 4157 11024
rect 4099 10983 4157 10984
rect 5163 11024 5205 11033
rect 5163 10984 5164 11024
rect 5204 10984 5205 11024
rect 5163 10975 5205 10984
rect 5451 11024 5493 11033
rect 5451 10984 5452 11024
rect 5492 10984 5493 11024
rect 5451 10975 5493 10984
rect 5643 11024 5685 11033
rect 5643 10984 5644 11024
rect 5684 10984 5685 11024
rect 5643 10975 5685 10984
rect 5835 11024 5877 11033
rect 5835 10984 5836 11024
rect 5876 10984 5877 11024
rect 5835 10975 5877 10984
rect 5923 11024 5981 11025
rect 5923 10984 5932 11024
rect 5972 10984 5981 11024
rect 5923 10983 5981 10984
rect 6315 11024 6357 11033
rect 6315 10984 6316 11024
rect 6356 10984 6357 11024
rect 6315 10975 6357 10984
rect 6411 11024 6453 11033
rect 6411 10984 6412 11024
rect 6452 10984 6453 11024
rect 6411 10975 6453 10984
rect 6691 11024 6749 11025
rect 6691 10984 6700 11024
rect 6740 10984 6749 11024
rect 6691 10983 6749 10984
rect 7171 11024 7229 11025
rect 7171 10984 7180 11024
rect 7220 10984 7229 11024
rect 7171 10983 7229 10984
rect 8419 11024 8477 11025
rect 8419 10984 8428 11024
rect 8468 10984 8477 11024
rect 8419 10983 8477 10984
rect 9195 11024 9237 11033
rect 9195 10984 9196 11024
rect 9236 10984 9237 11024
rect 9195 10975 9237 10984
rect 9379 11024 9437 11025
rect 9379 10984 9388 11024
rect 9428 10984 9437 11024
rect 9379 10983 9437 10984
rect 9571 11024 9629 11025
rect 9571 10984 9580 11024
rect 9620 10984 9629 11024
rect 9571 10983 9629 10984
rect 10819 11024 10877 11025
rect 10819 10984 10828 11024
rect 10868 10984 10877 11024
rect 10819 10983 10877 10984
rect 11307 11024 11349 11033
rect 11307 10984 11308 11024
rect 11348 10984 11349 11024
rect 11307 10975 11349 10984
rect 11403 11024 11445 11033
rect 11403 10984 11404 11024
rect 11444 10984 11445 11024
rect 11403 10975 11445 10984
rect 11883 11024 11925 11033
rect 11883 10984 11884 11024
rect 11924 10984 11925 11024
rect 11883 10975 11925 10984
rect 12355 11024 12413 11025
rect 12355 10984 12364 11024
rect 12404 10984 12413 11024
rect 13323 11024 13365 11033
rect 12355 10983 12413 10984
rect 12843 11010 12885 11019
rect 12843 10970 12844 11010
rect 12884 10970 12885 11010
rect 13323 10984 13324 11024
rect 13364 10984 13365 11024
rect 13323 10975 13365 10984
rect 13419 11024 13461 11033
rect 13419 10984 13420 11024
rect 13460 10984 13461 11024
rect 13419 10975 13461 10984
rect 13803 11024 13845 11033
rect 13803 10984 13804 11024
rect 13844 10984 13845 11024
rect 13803 10975 13845 10984
rect 14371 11024 14429 11025
rect 14371 10984 14380 11024
rect 14420 10984 14429 11024
rect 15435 11024 15477 11033
rect 14371 10983 14429 10984
rect 14859 11010 14901 11019
rect 12843 10961 12885 10970
rect 14859 10970 14860 11010
rect 14900 10970 14901 11010
rect 15435 10984 15436 11024
rect 15476 10984 15477 11024
rect 15435 10975 15477 10984
rect 15627 11024 15669 11033
rect 15627 10984 15628 11024
rect 15668 10984 15669 11024
rect 15627 10975 15669 10984
rect 15907 11024 15965 11025
rect 15907 10984 15916 11024
rect 15956 10984 15965 11024
rect 15907 10983 15965 10984
rect 16203 11024 16245 11033
rect 16203 10984 16204 11024
rect 16244 10984 16245 11024
rect 16203 10975 16245 10984
rect 16299 11024 16341 11033
rect 16299 10984 16300 11024
rect 16340 10984 16341 11024
rect 16299 10975 16341 10984
rect 16771 11024 16829 11025
rect 16771 10984 16780 11024
rect 16820 10984 16829 11024
rect 16771 10983 16829 10984
rect 16875 11024 16917 11033
rect 16875 10984 16876 11024
rect 16916 10984 16917 11024
rect 16875 10975 16917 10984
rect 17067 11024 17109 11033
rect 17067 10984 17068 11024
rect 17108 10984 17109 11024
rect 17067 10975 17109 10984
rect 17259 11024 17301 11033
rect 17259 10984 17260 11024
rect 17300 10984 17301 11024
rect 17259 10975 17301 10984
rect 17355 11024 17397 11033
rect 17355 10984 17356 11024
rect 17396 10984 17397 11024
rect 17355 10975 17397 10984
rect 17451 11024 17493 11033
rect 17451 10984 17452 11024
rect 17492 10984 17493 11024
rect 17451 10975 17493 10984
rect 17547 11024 17589 11033
rect 17547 10984 17548 11024
rect 17588 10984 17589 11024
rect 17547 10975 17589 10984
rect 17931 11024 17973 11033
rect 17931 10984 17932 11024
rect 17972 10984 17973 11024
rect 17931 10975 17973 10984
rect 18027 11024 18069 11033
rect 18027 10984 18028 11024
rect 18068 10984 18069 11024
rect 18027 10975 18069 10984
rect 18411 11024 18453 11033
rect 18411 10984 18412 11024
rect 18452 10984 18453 11024
rect 18411 10975 18453 10984
rect 18507 11024 18549 11033
rect 18507 10984 18508 11024
rect 18548 10984 18549 11024
rect 18507 10975 18549 10984
rect 18891 11024 18933 11033
rect 18891 10984 18892 11024
rect 18932 10984 18933 11024
rect 18891 10975 18933 10984
rect 19459 11024 19517 11025
rect 19459 10984 19468 11024
rect 19508 10984 19517 11024
rect 19459 10983 19517 10984
rect 19995 10982 20037 10991
rect 14859 10961 14901 10970
rect 11787 10940 11829 10949
rect 11787 10900 11788 10940
rect 11828 10900 11829 10940
rect 11787 10891 11829 10900
rect 13899 10940 13941 10949
rect 13899 10900 13900 10940
rect 13940 10900 13941 10940
rect 13899 10891 13941 10900
rect 18987 10940 19029 10949
rect 18987 10900 18988 10940
rect 19028 10900 19029 10940
rect 19995 10942 19996 10982
rect 20036 10942 20037 10982
rect 19995 10933 20037 10942
rect 18987 10891 19029 10900
rect 5451 10856 5493 10865
rect 5451 10816 5452 10856
rect 5492 10816 5493 10856
rect 5451 10807 5493 10816
rect 6891 10856 6933 10865
rect 6891 10816 6892 10856
rect 6932 10816 6933 10856
rect 6891 10807 6933 10816
rect 15435 10856 15477 10865
rect 15435 10816 15436 10856
rect 15476 10816 15477 10856
rect 15435 10807 15477 10816
rect 16579 10856 16637 10857
rect 16579 10816 16588 10856
rect 16628 10816 16637 10856
rect 16579 10815 16637 10816
rect 4299 10772 4341 10781
rect 4299 10732 4300 10772
rect 4340 10732 4341 10772
rect 4299 10723 4341 10732
rect 5643 10772 5685 10781
rect 5643 10732 5644 10772
rect 5684 10732 5685 10772
rect 5643 10723 5685 10732
rect 6603 10772 6645 10781
rect 6603 10732 6604 10772
rect 6644 10732 6645 10772
rect 6603 10723 6645 10732
rect 9291 10772 9333 10781
rect 9291 10732 9292 10772
rect 9332 10732 9333 10772
rect 9291 10723 9333 10732
rect 1152 10604 20352 10628
rect 1152 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 20352 10604
rect 1152 10540 20352 10564
rect 2667 10436 2709 10445
rect 2667 10396 2668 10436
rect 2708 10396 2709 10436
rect 2667 10387 2709 10396
rect 3435 10436 3477 10445
rect 3435 10396 3436 10436
rect 3476 10396 3477 10436
rect 3435 10387 3477 10396
rect 12843 10436 12885 10445
rect 12843 10396 12844 10436
rect 12884 10396 12885 10436
rect 12843 10387 12885 10396
rect 14763 10436 14805 10445
rect 14763 10396 14764 10436
rect 14804 10396 14805 10436
rect 14763 10387 14805 10396
rect 17163 10436 17205 10445
rect 17163 10396 17164 10436
rect 17204 10396 17205 10436
rect 17163 10387 17205 10396
rect 3819 10352 3861 10361
rect 3819 10312 3820 10352
rect 3860 10312 3861 10352
rect 3819 10303 3861 10312
rect 4587 10352 4629 10361
rect 4587 10312 4588 10352
rect 4628 10312 4629 10352
rect 4587 10303 4629 10312
rect 6979 10352 7037 10353
rect 6979 10312 6988 10352
rect 7028 10312 7037 10352
rect 6979 10311 7037 10312
rect 9195 10352 9237 10361
rect 9195 10312 9196 10352
rect 9236 10312 9237 10352
rect 9195 10303 9237 10312
rect 10819 10352 10877 10353
rect 10819 10312 10828 10352
rect 10868 10312 10877 10352
rect 10819 10311 10877 10312
rect 3723 10268 3765 10277
rect 3723 10228 3724 10268
rect 3764 10228 3765 10268
rect 3723 10219 3765 10228
rect 3915 10268 3957 10277
rect 3915 10228 3916 10268
rect 3956 10228 3957 10268
rect 3915 10219 3957 10228
rect 18315 10268 18357 10277
rect 18315 10228 18316 10268
rect 18356 10228 18357 10268
rect 18315 10219 18357 10228
rect 1219 10184 1277 10185
rect 1219 10144 1228 10184
rect 1268 10144 1277 10184
rect 1219 10143 1277 10144
rect 2467 10184 2525 10185
rect 2467 10144 2476 10184
rect 2516 10144 2525 10184
rect 2467 10143 2525 10144
rect 2851 10184 2909 10185
rect 2851 10144 2860 10184
rect 2900 10144 2909 10184
rect 2851 10143 2909 10144
rect 3147 10184 3189 10193
rect 3147 10144 3148 10184
rect 3188 10144 3189 10184
rect 3147 10135 3189 10144
rect 3435 10184 3477 10193
rect 3435 10144 3436 10184
rect 3476 10144 3477 10184
rect 3435 10135 3477 10144
rect 3619 10184 3677 10185
rect 3619 10144 3628 10184
rect 3668 10144 3677 10184
rect 3619 10143 3677 10144
rect 4011 10184 4053 10193
rect 4011 10144 4012 10184
rect 4052 10144 4053 10184
rect 4011 10135 4053 10144
rect 4203 10184 4245 10193
rect 4203 10144 4204 10184
rect 4244 10144 4245 10184
rect 4203 10135 4245 10144
rect 4387 10184 4445 10185
rect 4387 10144 4396 10184
rect 4436 10144 4445 10184
rect 4387 10143 4445 10144
rect 4587 10184 4629 10193
rect 4587 10144 4588 10184
rect 4628 10144 4629 10184
rect 4587 10135 4629 10144
rect 4779 10184 4821 10193
rect 4779 10144 4780 10184
rect 4820 10144 4821 10184
rect 4779 10135 4821 10144
rect 4867 10184 4925 10185
rect 4867 10144 4876 10184
rect 4916 10144 4925 10184
rect 4867 10143 4925 10144
rect 5150 10184 5208 10185
rect 5150 10144 5159 10184
rect 5199 10144 5208 10184
rect 5150 10143 5208 10144
rect 5259 10184 5301 10193
rect 5259 10144 5260 10184
rect 5300 10144 5301 10184
rect 5259 10135 5301 10144
rect 5355 10184 5397 10193
rect 5355 10144 5356 10184
rect 5396 10144 5397 10184
rect 5355 10135 5397 10144
rect 5539 10184 5597 10185
rect 5539 10144 5548 10184
rect 5588 10144 5597 10184
rect 5539 10143 5597 10144
rect 5635 10184 5693 10185
rect 5635 10144 5644 10184
rect 5684 10144 5693 10184
rect 5635 10143 5693 10144
rect 6027 10184 6069 10193
rect 6027 10144 6028 10184
rect 6068 10144 6069 10184
rect 6027 10135 6069 10144
rect 6315 10184 6357 10193
rect 6315 10144 6316 10184
rect 6356 10144 6357 10184
rect 6315 10135 6357 10144
rect 6987 10184 7029 10193
rect 6987 10144 6988 10184
rect 7028 10144 7029 10184
rect 6987 10135 7029 10144
rect 7083 10184 7125 10193
rect 7083 10144 7084 10184
rect 7124 10144 7125 10184
rect 7083 10135 7125 10144
rect 7275 10184 7317 10193
rect 7275 10144 7276 10184
rect 7316 10144 7317 10184
rect 7275 10135 7317 10144
rect 7555 10184 7613 10185
rect 7555 10144 7564 10184
rect 7604 10144 7613 10184
rect 7555 10143 7613 10144
rect 8803 10184 8861 10185
rect 8803 10144 8812 10184
rect 8852 10144 8861 10184
rect 8803 10143 8861 10144
rect 9475 10184 9533 10185
rect 9475 10144 9484 10184
rect 9524 10144 9533 10184
rect 9475 10143 9533 10144
rect 9579 10184 9621 10193
rect 9579 10144 9580 10184
rect 9620 10144 9621 10184
rect 9579 10135 9621 10144
rect 9763 10184 9821 10185
rect 9763 10144 9772 10184
rect 9812 10144 9821 10184
rect 9763 10143 9821 10144
rect 10147 10184 10205 10185
rect 10147 10144 10156 10184
rect 10196 10144 10205 10184
rect 10147 10143 10205 10144
rect 10443 10184 10485 10193
rect 10443 10144 10444 10184
rect 10484 10144 10485 10184
rect 10443 10135 10485 10144
rect 10539 10184 10581 10193
rect 10539 10144 10540 10184
rect 10580 10144 10581 10184
rect 10539 10135 10581 10144
rect 11019 10184 11061 10193
rect 11019 10144 11020 10184
rect 11060 10144 11061 10184
rect 11019 10135 11061 10144
rect 11211 10184 11253 10193
rect 11211 10144 11212 10184
rect 11252 10144 11253 10184
rect 11211 10135 11253 10144
rect 11395 10184 11453 10185
rect 11395 10144 11404 10184
rect 11444 10144 11453 10184
rect 11395 10143 11453 10144
rect 12643 10184 12701 10185
rect 12643 10144 12652 10184
rect 12692 10144 12701 10184
rect 12643 10143 12701 10144
rect 13315 10184 13373 10185
rect 13315 10144 13324 10184
rect 13364 10144 13373 10184
rect 13315 10143 13373 10144
rect 14563 10184 14621 10185
rect 14563 10144 14572 10184
rect 14612 10144 14621 10184
rect 14563 10143 14621 10144
rect 14955 10184 14997 10193
rect 14955 10144 14956 10184
rect 14996 10144 14997 10184
rect 14955 10135 14997 10144
rect 15051 10184 15093 10193
rect 15051 10144 15052 10184
rect 15092 10144 15093 10184
rect 15051 10135 15093 10144
rect 15715 10184 15773 10185
rect 15715 10144 15724 10184
rect 15764 10144 15773 10184
rect 15715 10143 15773 10144
rect 16963 10184 17021 10185
rect 16963 10144 16972 10184
rect 17012 10144 17021 10184
rect 16963 10143 17021 10144
rect 17739 10184 17781 10193
rect 17739 10144 17740 10184
rect 17780 10144 17781 10184
rect 17739 10135 17781 10144
rect 17835 10184 17877 10193
rect 17835 10144 17836 10184
rect 17876 10144 17877 10184
rect 17835 10135 17877 10144
rect 17931 10184 17973 10193
rect 17931 10144 17932 10184
rect 17972 10144 17973 10184
rect 17931 10135 17973 10144
rect 18027 10184 18069 10193
rect 18027 10144 18028 10184
rect 18068 10144 18069 10184
rect 18027 10135 18069 10144
rect 18219 10184 18261 10193
rect 18219 10144 18220 10184
rect 18260 10144 18261 10184
rect 18691 10184 18749 10185
rect 18219 10135 18261 10144
rect 18500 10169 18558 10170
rect 18500 10129 18509 10169
rect 18549 10129 18558 10169
rect 18691 10144 18700 10184
rect 18740 10144 18749 10184
rect 18691 10143 18749 10144
rect 19939 10184 19997 10185
rect 19939 10144 19948 10184
rect 19988 10144 19997 10184
rect 19939 10143 19997 10144
rect 18500 10128 18558 10129
rect 2955 10100 2997 10109
rect 2955 10060 2956 10100
rect 2996 10060 2997 10100
rect 2955 10051 2997 10060
rect 4299 10100 4341 10109
rect 4299 10060 4300 10100
rect 4340 10060 4341 10100
rect 4299 10051 4341 10060
rect 9003 10100 9045 10109
rect 9003 10060 9004 10100
rect 9044 10060 9045 10100
rect 9003 10051 9045 10060
rect 11115 10100 11157 10109
rect 11115 10060 11116 10100
rect 11156 10060 11157 10100
rect 11115 10051 11157 10060
rect 20139 10100 20181 10109
rect 20139 10060 20140 10100
rect 20180 10060 20181 10100
rect 20139 10051 20181 10060
rect 5347 10016 5405 10017
rect 5347 9976 5356 10016
rect 5396 9976 5405 10016
rect 5347 9975 5405 9976
rect 6123 10016 6165 10025
rect 6123 9976 6124 10016
rect 6164 9976 6165 10016
rect 6123 9967 6165 9976
rect 6699 10016 6741 10025
rect 6699 9976 6700 10016
rect 6740 9976 6741 10016
rect 6699 9967 6741 9976
rect 9771 10016 9813 10025
rect 9771 9976 9772 10016
rect 9812 9976 9813 10016
rect 9771 9967 9813 9976
rect 15235 10016 15293 10017
rect 15235 9976 15244 10016
rect 15284 9976 15293 10016
rect 15235 9975 15293 9976
rect 17347 10016 17405 10017
rect 17347 9976 17356 10016
rect 17396 9976 17405 10016
rect 17347 9975 17405 9976
rect 1152 9848 20452 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20452 9848
rect 1152 9784 20452 9808
rect 4683 9722 4725 9731
rect 3051 9680 3093 9689
rect 3051 9640 3052 9680
rect 3092 9640 3093 9680
rect 4683 9682 4684 9722
rect 4724 9682 4725 9722
rect 4683 9673 4725 9682
rect 5643 9680 5685 9689
rect 3051 9631 3093 9640
rect 5643 9640 5644 9680
rect 5684 9640 5685 9680
rect 5643 9631 5685 9640
rect 6691 9680 6749 9681
rect 6691 9640 6700 9680
rect 6740 9640 6749 9680
rect 6691 9639 6749 9640
rect 8715 9680 8757 9689
rect 8715 9640 8716 9680
rect 8756 9640 8757 9680
rect 8715 9631 8757 9640
rect 9195 9680 9237 9689
rect 9195 9640 9196 9680
rect 9236 9640 9237 9680
rect 9195 9631 9237 9640
rect 13131 9680 13173 9689
rect 13131 9640 13132 9680
rect 13172 9640 13173 9680
rect 13131 9631 13173 9640
rect 14467 9680 14525 9681
rect 14467 9640 14476 9680
rect 14516 9640 14525 9680
rect 14467 9639 14525 9640
rect 16779 9680 16821 9689
rect 16779 9640 16780 9680
rect 16820 9640 16821 9680
rect 16779 9631 16821 9640
rect 19083 9680 19125 9689
rect 19083 9640 19084 9680
rect 19124 9640 19125 9680
rect 19083 9631 19125 9640
rect 1603 9512 1661 9513
rect 1603 9472 1612 9512
rect 1652 9472 1661 9512
rect 1603 9471 1661 9472
rect 2851 9512 2909 9513
rect 2851 9472 2860 9512
rect 2900 9472 2909 9512
rect 2851 9471 2909 9472
rect 3715 9511 3757 9520
rect 3715 9471 3716 9511
rect 3756 9471 3757 9511
rect 4003 9512 4061 9513
rect 4003 9472 4012 9512
rect 4052 9472 4061 9512
rect 4003 9471 4061 9472
rect 4299 9512 4341 9521
rect 4299 9472 4300 9512
rect 4340 9472 4341 9512
rect 3715 9462 3757 9471
rect 4299 9463 4341 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4875 9512 4917 9521
rect 4875 9472 4876 9512
rect 4916 9472 4917 9512
rect 4875 9463 4917 9472
rect 4971 9512 5013 9521
rect 4971 9472 4972 9512
rect 5012 9472 5013 9512
rect 4971 9463 5013 9472
rect 5067 9512 5109 9521
rect 5067 9472 5068 9512
rect 5108 9472 5109 9512
rect 5067 9463 5109 9472
rect 5163 9512 5205 9521
rect 5163 9472 5164 9512
rect 5204 9472 5205 9512
rect 5163 9463 5205 9472
rect 5547 9512 5589 9521
rect 5547 9472 5548 9512
rect 5588 9472 5589 9512
rect 5547 9463 5589 9472
rect 5835 9512 5877 9521
rect 5835 9472 5836 9512
rect 5876 9472 5877 9512
rect 5835 9463 5877 9472
rect 6027 9512 6069 9521
rect 6027 9472 6028 9512
rect 6068 9472 6069 9512
rect 6307 9512 6365 9513
rect 6027 9463 6069 9472
rect 6211 9498 6269 9499
rect 6211 9458 6220 9498
rect 6260 9458 6269 9498
rect 6307 9472 6316 9512
rect 6356 9472 6365 9512
rect 6307 9471 6365 9472
rect 6987 9512 7029 9521
rect 6987 9472 6988 9512
rect 7028 9472 7029 9512
rect 6987 9463 7029 9472
rect 7083 9512 7125 9521
rect 7083 9472 7084 9512
rect 7124 9472 7125 9512
rect 7563 9512 7605 9521
rect 7083 9463 7125 9472
rect 7467 9470 7509 9479
rect 6211 9457 6269 9458
rect 7467 9430 7468 9470
rect 7508 9430 7509 9470
rect 7563 9472 7564 9512
rect 7604 9472 7605 9512
rect 7563 9463 7605 9472
rect 8035 9512 8093 9513
rect 8035 9472 8044 9512
rect 8084 9472 8093 9512
rect 9667 9512 9725 9513
rect 8035 9471 8093 9472
rect 8523 9498 8565 9507
rect 8523 9458 8524 9498
rect 8564 9458 8565 9498
rect 9667 9472 9676 9512
rect 9716 9472 9725 9512
rect 9667 9471 9725 9472
rect 10915 9512 10973 9513
rect 10915 9472 10924 9512
rect 10964 9472 10973 9512
rect 10915 9471 10973 9472
rect 11683 9512 11741 9513
rect 11683 9472 11692 9512
rect 11732 9472 11741 9512
rect 11683 9471 11741 9472
rect 12931 9512 12989 9513
rect 12931 9472 12940 9512
rect 12980 9472 12989 9512
rect 12931 9471 12989 9472
rect 13611 9512 13653 9521
rect 13611 9472 13612 9512
rect 13652 9472 13653 9512
rect 13611 9463 13653 9472
rect 13707 9512 13749 9521
rect 13707 9472 13708 9512
rect 13748 9472 13749 9512
rect 13707 9463 13749 9472
rect 13803 9512 13845 9521
rect 13803 9472 13804 9512
rect 13844 9472 13845 9512
rect 13803 9463 13845 9472
rect 13899 9512 13941 9521
rect 13899 9472 13900 9512
rect 13940 9472 13941 9512
rect 13899 9463 13941 9472
rect 14275 9512 14333 9513
rect 14275 9472 14284 9512
rect 14324 9472 14333 9512
rect 14275 9471 14333 9472
rect 14371 9512 14429 9513
rect 14371 9472 14380 9512
rect 14420 9472 14429 9512
rect 14371 9471 14429 9472
rect 14571 9512 14613 9521
rect 14571 9472 14572 9512
rect 14612 9472 14613 9512
rect 14571 9463 14613 9472
rect 14667 9512 14709 9521
rect 14667 9472 14668 9512
rect 14708 9472 14709 9512
rect 14667 9463 14709 9472
rect 14814 9512 14872 9513
rect 14814 9472 14823 9512
rect 14863 9472 14872 9512
rect 14814 9471 14872 9472
rect 15331 9512 15389 9513
rect 15331 9472 15340 9512
rect 15380 9472 15389 9512
rect 15331 9471 15389 9472
rect 16579 9512 16637 9513
rect 16579 9472 16588 9512
rect 16628 9472 16637 9512
rect 16579 9471 16637 9472
rect 17635 9512 17693 9513
rect 17635 9472 17644 9512
rect 17684 9472 17693 9512
rect 17635 9471 17693 9472
rect 18883 9512 18941 9513
rect 18883 9472 18892 9512
rect 18932 9472 18941 9512
rect 18883 9471 18941 9472
rect 19358 9512 19416 9513
rect 19358 9472 19367 9512
rect 19407 9472 19416 9512
rect 19358 9471 19416 9472
rect 19467 9512 19509 9521
rect 19467 9472 19468 9512
rect 19508 9472 19509 9512
rect 19467 9463 19509 9472
rect 19563 9512 19605 9521
rect 19563 9472 19564 9512
rect 19604 9472 19605 9512
rect 19563 9463 19605 9472
rect 19747 9512 19805 9513
rect 19747 9472 19756 9512
rect 19796 9472 19805 9512
rect 19747 9471 19805 9472
rect 19843 9512 19901 9513
rect 19843 9472 19852 9512
rect 19892 9472 19901 9512
rect 19843 9471 19901 9472
rect 20043 9512 20085 9521
rect 20043 9472 20044 9512
rect 20084 9472 20085 9512
rect 20043 9463 20085 9472
rect 20235 9512 20277 9521
rect 20235 9472 20236 9512
rect 20276 9472 20277 9512
rect 20235 9463 20277 9472
rect 8523 9449 8565 9458
rect 7467 9421 7509 9430
rect 20139 9428 20181 9437
rect 20139 9388 20140 9428
rect 20180 9388 20181 9428
rect 20139 9379 20181 9388
rect 3627 9344 3669 9353
rect 3627 9304 3628 9344
rect 3668 9304 3669 9344
rect 3627 9295 3669 9304
rect 6027 9344 6069 9353
rect 6027 9304 6028 9344
rect 6068 9304 6069 9344
rect 6027 9295 6069 9304
rect 15051 9344 15093 9353
rect 15051 9304 15052 9344
rect 15092 9304 15093 9344
rect 15051 9295 15093 9304
rect 17355 9344 17397 9353
rect 17355 9304 17356 9344
rect 17396 9304 17397 9344
rect 17355 9295 17397 9304
rect 3051 9260 3093 9269
rect 3051 9220 3052 9260
rect 3092 9220 3093 9260
rect 3051 9211 3093 9220
rect 11115 9260 11157 9269
rect 11115 9220 11116 9260
rect 11156 9220 11157 9260
rect 11115 9211 11157 9220
rect 19083 9260 19125 9269
rect 19083 9220 19084 9260
rect 19124 9220 19125 9260
rect 19083 9211 19125 9220
rect 19851 9260 19893 9269
rect 19851 9220 19852 9260
rect 19892 9220 19893 9260
rect 19851 9211 19893 9220
rect 1152 9092 20352 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 20352 9092
rect 1152 9028 20352 9052
rect 3915 8924 3957 8933
rect 3915 8884 3916 8924
rect 3956 8884 3957 8924
rect 3915 8875 3957 8884
rect 6315 8924 6357 8933
rect 6315 8884 6316 8924
rect 6356 8884 6357 8924
rect 6315 8875 6357 8884
rect 8331 8924 8373 8933
rect 8331 8884 8332 8924
rect 8372 8884 8373 8924
rect 8331 8875 8373 8884
rect 14763 8924 14805 8933
rect 14763 8884 14764 8924
rect 14804 8884 14805 8924
rect 14763 8875 14805 8884
rect 19083 8924 19125 8933
rect 19083 8884 19084 8924
rect 19124 8884 19125 8924
rect 19083 8875 19125 8884
rect 3339 8840 3381 8849
rect 3339 8800 3340 8840
rect 3380 8800 3381 8840
rect 3339 8791 3381 8800
rect 15339 8840 15381 8849
rect 15339 8800 15340 8840
rect 15380 8800 15381 8840
rect 15339 8791 15381 8800
rect 20235 8840 20277 8849
rect 20235 8800 20236 8840
rect 20276 8800 20277 8840
rect 20235 8791 20277 8800
rect 4491 8756 4533 8765
rect 4491 8716 4492 8756
rect 4532 8716 4533 8756
rect 4491 8707 4533 8716
rect 9291 8756 9333 8765
rect 9291 8716 9292 8756
rect 9332 8716 9333 8756
rect 9291 8707 9333 8716
rect 20035 8756 20093 8757
rect 20035 8716 20044 8756
rect 20084 8716 20093 8756
rect 20035 8715 20093 8716
rect 10299 8681 10341 8690
rect 19816 8687 19858 8696
rect 1891 8672 1949 8673
rect 1891 8632 1900 8672
rect 1940 8632 1949 8672
rect 1891 8631 1949 8632
rect 3139 8672 3197 8673
rect 3139 8632 3148 8672
rect 3188 8632 3197 8672
rect 3139 8631 3197 8632
rect 3907 8672 3965 8673
rect 3907 8632 3916 8672
rect 3956 8632 3965 8672
rect 3907 8631 3965 8632
rect 4107 8672 4149 8681
rect 4107 8632 4108 8672
rect 4148 8632 4149 8672
rect 4107 8623 4149 8632
rect 4195 8672 4253 8673
rect 4195 8632 4204 8672
rect 4244 8632 4253 8672
rect 4195 8631 4253 8632
rect 4395 8672 4437 8681
rect 4395 8632 4396 8672
rect 4436 8632 4437 8672
rect 4395 8623 4437 8632
rect 4683 8672 4725 8681
rect 4683 8632 4684 8672
rect 4724 8632 4725 8672
rect 4683 8623 4725 8632
rect 4867 8672 4925 8673
rect 4867 8632 4876 8672
rect 4916 8632 4925 8672
rect 4867 8631 4925 8632
rect 6115 8672 6173 8673
rect 6115 8632 6124 8672
rect 6164 8632 6173 8672
rect 6115 8631 6173 8632
rect 6883 8672 6941 8673
rect 6883 8632 6892 8672
rect 6932 8632 6941 8672
rect 6883 8631 6941 8632
rect 8131 8672 8189 8673
rect 8131 8632 8140 8672
rect 8180 8632 8189 8672
rect 8131 8631 8189 8632
rect 8715 8672 8757 8681
rect 8715 8632 8716 8672
rect 8756 8632 8757 8672
rect 8715 8623 8757 8632
rect 8811 8672 8853 8681
rect 8811 8632 8812 8672
rect 8852 8632 8853 8672
rect 8811 8623 8853 8632
rect 9195 8672 9237 8681
rect 9195 8632 9196 8672
rect 9236 8632 9237 8672
rect 9195 8623 9237 8632
rect 9763 8672 9821 8673
rect 9763 8632 9772 8672
rect 9812 8632 9821 8672
rect 10299 8641 10300 8681
rect 10340 8641 10341 8681
rect 10299 8632 10341 8641
rect 10731 8672 10773 8681
rect 10731 8632 10732 8672
rect 10772 8632 10773 8672
rect 9763 8631 9821 8632
rect 10731 8623 10773 8632
rect 10827 8672 10869 8681
rect 10827 8632 10828 8672
rect 10868 8632 10869 8672
rect 10827 8623 10869 8632
rect 11203 8672 11261 8673
rect 11203 8632 11212 8672
rect 11252 8632 11261 8672
rect 11203 8631 11261 8632
rect 12451 8672 12509 8673
rect 12451 8632 12460 8672
rect 12500 8632 12509 8672
rect 12451 8631 12509 8632
rect 13315 8672 13373 8673
rect 13315 8632 13324 8672
rect 13364 8632 13373 8672
rect 13315 8631 13373 8632
rect 14563 8672 14621 8673
rect 14563 8632 14572 8672
rect 14612 8632 14621 8672
rect 14563 8631 14621 8632
rect 15427 8672 15485 8673
rect 15427 8632 15436 8672
rect 15476 8632 15485 8672
rect 15427 8631 15485 8632
rect 16875 8672 16917 8681
rect 16875 8632 16876 8672
rect 16916 8632 16917 8672
rect 16875 8623 16917 8632
rect 16971 8672 17013 8681
rect 16971 8632 16972 8672
rect 17012 8632 17013 8672
rect 16971 8623 17013 8632
rect 17635 8672 17693 8673
rect 17635 8632 17644 8672
rect 17684 8632 17693 8672
rect 17635 8631 17693 8632
rect 18883 8672 18941 8673
rect 18883 8632 18892 8672
rect 18932 8632 18941 8672
rect 18883 8631 18941 8632
rect 19267 8672 19325 8673
rect 19267 8632 19276 8672
rect 19316 8632 19325 8672
rect 19267 8631 19325 8632
rect 19363 8672 19421 8673
rect 19363 8632 19372 8672
rect 19412 8632 19421 8672
rect 19363 8631 19421 8632
rect 19563 8672 19605 8681
rect 19563 8632 19564 8672
rect 19604 8632 19605 8672
rect 19563 8623 19605 8632
rect 19659 8672 19701 8681
rect 19659 8632 19660 8672
rect 19700 8632 19701 8672
rect 19816 8647 19817 8687
rect 19857 8647 19858 8687
rect 19816 8638 19858 8647
rect 19659 8623 19701 8632
rect 6603 8504 6645 8513
rect 6603 8464 6604 8504
rect 6644 8464 6645 8504
rect 6603 8455 6645 8464
rect 10443 8504 10485 8513
rect 10443 8464 10444 8504
rect 10484 8464 10485 8504
rect 10443 8455 10485 8464
rect 11011 8504 11069 8505
rect 11011 8464 11020 8504
rect 11060 8464 11069 8504
rect 11011 8463 11069 8464
rect 12651 8504 12693 8513
rect 12651 8464 12652 8504
rect 12692 8464 12693 8504
rect 12651 8455 12693 8464
rect 15043 8504 15101 8505
rect 15043 8464 15052 8504
rect 15092 8464 15101 8504
rect 15043 8463 15101 8464
rect 17155 8504 17213 8505
rect 17155 8464 17164 8504
rect 17204 8464 17213 8504
rect 17155 8463 17213 8464
rect 17347 8504 17405 8505
rect 17347 8464 17356 8504
rect 17396 8464 17405 8504
rect 17347 8463 17405 8464
rect 19083 8504 19125 8513
rect 19083 8464 19084 8504
rect 19124 8464 19125 8504
rect 19083 8455 19125 8464
rect 19747 8504 19805 8505
rect 19747 8464 19756 8504
rect 19796 8464 19805 8504
rect 19747 8463 19805 8464
rect 1152 8336 20452 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20452 8336
rect 1152 8272 20452 8296
rect 3619 8168 3677 8169
rect 3619 8128 3628 8168
rect 3668 8128 3677 8168
rect 3619 8127 3677 8128
rect 3915 8168 3957 8177
rect 3915 8128 3916 8168
rect 3956 8128 3957 8168
rect 3915 8119 3957 8128
rect 8619 8168 8661 8177
rect 8619 8128 8620 8168
rect 8660 8128 8661 8168
rect 8619 8119 8661 8128
rect 10347 8168 10389 8177
rect 10347 8128 10348 8168
rect 10388 8128 10389 8168
rect 10347 8119 10389 8128
rect 14859 8168 14901 8177
rect 14859 8128 14860 8168
rect 14900 8128 14901 8168
rect 14859 8119 14901 8128
rect 19747 8168 19805 8169
rect 19747 8128 19756 8168
rect 19796 8128 19805 8168
rect 19747 8127 19805 8128
rect 20139 8168 20181 8177
rect 20139 8128 20140 8168
rect 20180 8128 20181 8168
rect 20139 8119 20181 8128
rect 12747 8084 12789 8093
rect 12747 8044 12748 8084
rect 12788 8044 12789 8084
rect 12747 8035 12789 8044
rect 2955 8000 2997 8009
rect 2955 7960 2956 8000
rect 2996 7960 2997 8000
rect 2955 7951 2997 7960
rect 3051 8000 3093 8009
rect 3051 7960 3052 8000
rect 3092 7960 3093 8000
rect 3051 7951 3093 7960
rect 3147 8000 3189 8009
rect 3147 7960 3148 8000
rect 3188 7960 3189 8000
rect 3147 7951 3189 7960
rect 3243 8000 3285 8009
rect 3243 7960 3244 8000
rect 3284 7960 3285 8000
rect 3243 7951 3285 7960
rect 3427 8000 3485 8001
rect 3427 7960 3436 8000
rect 3476 7960 3485 8000
rect 3427 7959 3485 7960
rect 3531 8000 3573 8009
rect 3531 7960 3532 8000
rect 3572 7960 3573 8000
rect 3531 7951 3573 7960
rect 3723 8000 3765 8009
rect 3723 7960 3724 8000
rect 3764 7960 3765 8000
rect 3723 7951 3765 7960
rect 3907 8000 3965 8001
rect 3907 7960 3916 8000
rect 3956 7960 3965 8000
rect 3907 7959 3965 7960
rect 4107 8000 4149 8009
rect 4107 7960 4108 8000
rect 4148 7960 4149 8000
rect 4107 7951 4149 7960
rect 4195 8000 4253 8001
rect 4195 7960 4204 8000
rect 4244 7960 4253 8000
rect 4195 7959 4253 7960
rect 4683 8000 4725 8009
rect 4683 7960 4684 8000
rect 4724 7960 4725 8000
rect 4683 7951 4725 7960
rect 4779 8000 4821 8009
rect 4779 7960 4780 8000
rect 4820 7960 4821 8000
rect 4779 7951 4821 7960
rect 4971 8000 5013 8009
rect 4971 7960 4972 8000
rect 5012 7960 5013 8000
rect 4971 7951 5013 7960
rect 7171 8000 7229 8001
rect 7171 7960 7180 8000
rect 7220 7960 7229 8000
rect 7171 7959 7229 7960
rect 8419 8000 8477 8001
rect 8419 7960 8428 8000
rect 8468 7960 8477 8000
rect 8419 7959 8477 7960
rect 8899 8000 8957 8001
rect 8899 7960 8908 8000
rect 8948 7960 8957 8000
rect 8899 7959 8957 7960
rect 10147 8000 10205 8001
rect 10147 7960 10156 8000
rect 10196 7960 10205 8000
rect 10147 7959 10205 7960
rect 11019 8000 11061 8009
rect 11019 7960 11020 8000
rect 11060 7960 11061 8000
rect 11019 7951 11061 7960
rect 11115 8000 11157 8009
rect 11115 7960 11116 8000
rect 11156 7960 11157 8000
rect 11115 7951 11157 7960
rect 12067 8000 12125 8001
rect 12067 7960 12076 8000
rect 12116 7960 12125 8000
rect 13411 8000 13469 8001
rect 12067 7959 12125 7960
rect 12603 7990 12645 7999
rect 12603 7950 12604 7990
rect 12644 7950 12645 7990
rect 13411 7960 13420 8000
rect 13460 7960 13469 8000
rect 13411 7959 13469 7960
rect 14659 8000 14717 8001
rect 14659 7960 14668 8000
rect 14708 7960 14717 8000
rect 14659 7959 14717 7960
rect 17635 8000 17693 8001
rect 17635 7960 17644 8000
rect 17684 7960 17693 8000
rect 17635 7959 17693 7960
rect 18883 8000 18941 8001
rect 18883 7960 18892 8000
rect 18932 7960 18941 8000
rect 18883 7959 18941 7960
rect 19467 8000 19509 8009
rect 19467 7960 19468 8000
rect 19508 7960 19509 8000
rect 19467 7951 19509 7960
rect 19563 8000 19605 8009
rect 19563 7960 19564 8000
rect 19604 7960 19605 8000
rect 19563 7951 19605 7960
rect 19947 8000 19989 8009
rect 19947 7960 19948 8000
rect 19988 7960 19989 8000
rect 19947 7951 19989 7960
rect 20043 8000 20085 8009
rect 20043 7960 20044 8000
rect 20084 7960 20085 8000
rect 20043 7951 20085 7960
rect 20235 8000 20277 8009
rect 20235 7960 20236 8000
rect 20276 7960 20277 8000
rect 20235 7951 20277 7960
rect 12603 7941 12645 7950
rect 11499 7916 11541 7925
rect 11499 7876 11500 7916
rect 11540 7876 11541 7916
rect 11499 7867 11541 7876
rect 11595 7916 11637 7925
rect 11595 7876 11596 7916
rect 11636 7876 11637 7916
rect 11595 7867 11637 7876
rect 4675 7832 4733 7833
rect 4675 7792 4684 7832
rect 4724 7792 4733 7832
rect 4675 7791 4733 7792
rect 6315 7832 6357 7841
rect 6315 7792 6316 7832
rect 6356 7792 6357 7832
rect 6315 7783 6357 7792
rect 6603 7832 6645 7841
rect 6603 7792 6604 7832
rect 6644 7792 6645 7832
rect 6603 7783 6645 7792
rect 15051 7832 15093 7841
rect 15051 7792 15052 7832
rect 15092 7792 15093 7832
rect 15051 7783 15093 7792
rect 17355 7832 17397 7841
rect 17355 7792 17356 7832
rect 17396 7792 17397 7832
rect 17355 7783 17397 7792
rect 19083 7748 19125 7757
rect 19083 7708 19084 7748
rect 19124 7708 19125 7748
rect 19083 7699 19125 7708
rect 1152 7580 20352 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 20352 7580
rect 1152 7516 20352 7540
rect 4491 7412 4533 7421
rect 4491 7372 4492 7412
rect 4532 7372 4533 7412
rect 4491 7363 4533 7372
rect 20235 7412 20277 7421
rect 20235 7372 20236 7412
rect 20276 7372 20277 7412
rect 20235 7363 20277 7372
rect 12363 7328 12405 7337
rect 12363 7288 12364 7328
rect 12404 7288 12405 7328
rect 12363 7279 12405 7288
rect 15051 7328 15093 7337
rect 15051 7288 15052 7328
rect 15092 7288 15093 7328
rect 15051 7279 15093 7288
rect 18795 7328 18837 7337
rect 18795 7288 18796 7328
rect 18836 7288 18837 7328
rect 18795 7279 18837 7288
rect 19267 7328 19325 7329
rect 19267 7288 19276 7328
rect 19316 7288 19325 7328
rect 19267 7287 19325 7288
rect 8811 7244 8853 7253
rect 8811 7204 8812 7244
rect 8852 7204 8853 7244
rect 8811 7195 8853 7204
rect 13131 7244 13173 7253
rect 13131 7204 13132 7244
rect 13172 7204 13173 7244
rect 13131 7195 13173 7204
rect 13227 7244 13269 7253
rect 13227 7204 13228 7244
rect 13268 7204 13269 7244
rect 13227 7195 13269 7204
rect 16011 7244 16053 7253
rect 16011 7204 16012 7244
rect 16052 7204 16053 7244
rect 16011 7195 16053 7204
rect 20035 7244 20093 7245
rect 20035 7204 20044 7244
rect 20084 7204 20093 7244
rect 20035 7203 20093 7204
rect 9819 7169 9861 7178
rect 4203 7160 4245 7169
rect 4203 7120 4204 7160
rect 4244 7120 4245 7160
rect 4203 7111 4245 7120
rect 4491 7160 4533 7169
rect 4491 7120 4492 7160
rect 4532 7120 4533 7160
rect 4491 7111 4533 7120
rect 6499 7160 6557 7161
rect 6499 7120 6508 7160
rect 6548 7120 6557 7160
rect 6499 7119 6557 7120
rect 7747 7160 7805 7161
rect 7747 7120 7756 7160
rect 7796 7120 7805 7160
rect 7747 7119 7805 7120
rect 8235 7160 8277 7169
rect 8235 7120 8236 7160
rect 8276 7120 8277 7160
rect 8235 7111 8277 7120
rect 8331 7160 8373 7169
rect 8331 7120 8332 7160
rect 8372 7120 8373 7160
rect 8331 7111 8373 7120
rect 8715 7160 8757 7169
rect 8715 7120 8716 7160
rect 8756 7120 8757 7160
rect 8715 7111 8757 7120
rect 9283 7160 9341 7161
rect 9283 7120 9292 7160
rect 9332 7120 9341 7160
rect 9819 7129 9820 7169
rect 9860 7129 9861 7169
rect 9819 7120 9861 7129
rect 10915 7160 10973 7161
rect 10915 7120 10924 7160
rect 10964 7120 10973 7160
rect 9283 7119 9341 7120
rect 10915 7119 10973 7120
rect 12163 7160 12221 7161
rect 12163 7120 12172 7160
rect 12212 7120 12221 7160
rect 12163 7119 12221 7120
rect 12651 7160 12693 7169
rect 12651 7120 12652 7160
rect 12692 7120 12693 7160
rect 12651 7111 12693 7120
rect 12747 7160 12789 7169
rect 14187 7165 14229 7174
rect 12747 7120 12748 7160
rect 12788 7120 12789 7160
rect 12747 7111 12789 7120
rect 13699 7160 13757 7161
rect 13699 7120 13708 7160
rect 13748 7120 13757 7160
rect 13699 7119 13757 7120
rect 14187 7125 14188 7165
rect 14228 7125 14229 7165
rect 14187 7116 14229 7125
rect 15435 7160 15477 7169
rect 15435 7120 15436 7160
rect 15476 7120 15477 7160
rect 15435 7111 15477 7120
rect 15531 7160 15573 7169
rect 15531 7120 15532 7160
rect 15572 7120 15573 7160
rect 15531 7111 15573 7120
rect 15915 7160 15957 7169
rect 16971 7165 17013 7174
rect 15915 7120 15916 7160
rect 15956 7120 15957 7160
rect 15915 7111 15957 7120
rect 16483 7160 16541 7161
rect 16483 7120 16492 7160
rect 16532 7120 16541 7160
rect 16483 7119 16541 7120
rect 16971 7125 16972 7165
rect 17012 7125 17013 7165
rect 16971 7116 17013 7125
rect 17347 7160 17405 7161
rect 17347 7120 17356 7160
rect 17396 7120 17405 7160
rect 17347 7119 17405 7120
rect 18595 7160 18653 7161
rect 18595 7120 18604 7160
rect 18644 7120 18653 7160
rect 18595 7119 18653 7120
rect 18987 7160 19029 7169
rect 18987 7120 18988 7160
rect 19028 7120 19029 7160
rect 18987 7111 19029 7120
rect 19179 7160 19221 7169
rect 19179 7120 19180 7160
rect 19220 7120 19221 7160
rect 19179 7111 19221 7120
rect 19275 7160 19317 7169
rect 19275 7120 19276 7160
rect 19316 7120 19317 7160
rect 19275 7111 19317 7120
rect 19755 7160 19797 7169
rect 19755 7120 19756 7160
rect 19796 7120 19797 7160
rect 19755 7111 19797 7120
rect 19851 7160 19893 7169
rect 19851 7120 19852 7160
rect 19892 7120 19893 7160
rect 19851 7111 19893 7120
rect 7947 7076 7989 7085
rect 7947 7036 7948 7076
rect 7988 7036 7989 7076
rect 7947 7027 7989 7036
rect 17163 7076 17205 7085
rect 17163 7036 17164 7076
rect 17204 7036 17205 7076
rect 17163 7027 17205 7036
rect 9963 6992 10005 7001
rect 9963 6952 9964 6992
rect 10004 6952 10005 6992
rect 9963 6943 10005 6952
rect 14379 6992 14421 7001
rect 14379 6952 14380 6992
rect 14420 6952 14421 6992
rect 14379 6943 14421 6952
rect 19555 6992 19613 6993
rect 19555 6952 19564 6992
rect 19604 6952 19613 6992
rect 19555 6951 19613 6952
rect 1152 6824 20452 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20452 6824
rect 1152 6760 20452 6784
rect 6603 6656 6645 6665
rect 6603 6616 6604 6656
rect 6644 6616 6645 6656
rect 6603 6607 6645 6616
rect 9867 6656 9909 6665
rect 9867 6616 9868 6656
rect 9908 6616 9909 6656
rect 9867 6607 9909 6616
rect 14187 6656 14229 6665
rect 14187 6616 14188 6656
rect 14228 6616 14229 6656
rect 14187 6607 14229 6616
rect 16491 6656 16533 6665
rect 16491 6616 16492 6656
rect 16532 6616 16533 6656
rect 16491 6607 16533 6616
rect 20139 6656 20181 6665
rect 20139 6616 20140 6656
rect 20180 6616 20181 6656
rect 20139 6607 20181 6616
rect 8419 6488 8477 6489
rect 8419 6448 8428 6488
rect 8468 6448 8477 6488
rect 8419 6447 8477 6448
rect 9667 6488 9725 6489
rect 9667 6448 9676 6488
rect 9716 6448 9725 6488
rect 9667 6447 9725 6448
rect 12739 6488 12797 6489
rect 12739 6448 12748 6488
rect 12788 6448 12797 6488
rect 12739 6447 12797 6448
rect 13987 6488 14045 6489
rect 13987 6448 13996 6488
rect 14036 6448 14045 6488
rect 13987 6447 14045 6448
rect 15043 6488 15101 6489
rect 15043 6448 15052 6488
rect 15092 6448 15101 6488
rect 15043 6447 15101 6448
rect 16291 6488 16349 6489
rect 16291 6448 16300 6488
rect 16340 6448 16349 6488
rect 16291 6447 16349 6448
rect 18691 6488 18749 6489
rect 18691 6448 18700 6488
rect 18740 6448 18749 6488
rect 18691 6447 18749 6448
rect 19939 6488 19997 6489
rect 19939 6448 19948 6488
rect 19988 6448 19997 6488
rect 19939 6447 19997 6448
rect 10147 6404 10205 6405
rect 10147 6364 10156 6404
rect 10196 6364 10205 6404
rect 10147 6363 10205 6364
rect 11683 6404 11741 6405
rect 11683 6364 11692 6404
rect 11732 6364 11741 6404
rect 11683 6363 11741 6364
rect 11499 6320 11541 6329
rect 11499 6280 11500 6320
rect 11540 6280 11541 6320
rect 11499 6271 11541 6280
rect 17355 6320 17397 6329
rect 17355 6280 17356 6320
rect 17396 6280 17397 6320
rect 17355 6271 17397 6280
rect 10347 6236 10389 6245
rect 10347 6196 10348 6236
rect 10388 6196 10389 6236
rect 10347 6187 10389 6196
rect 1152 6068 20352 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 20352 6068
rect 1152 6004 20352 6028
rect 14859 5900 14901 5909
rect 14859 5860 14860 5900
rect 14900 5860 14901 5900
rect 14859 5851 14901 5860
rect 6603 5816 6645 5825
rect 6603 5776 6604 5816
rect 6644 5776 6645 5816
rect 6603 5767 6645 5776
rect 15051 5816 15093 5825
rect 15051 5776 15052 5816
rect 15092 5776 15093 5816
rect 15051 5767 15093 5776
rect 13411 5648 13469 5649
rect 13411 5608 13420 5648
rect 13460 5608 13469 5648
rect 13411 5607 13469 5608
rect 14659 5648 14717 5649
rect 14659 5608 14668 5648
rect 14708 5608 14717 5648
rect 14659 5607 14717 5608
rect 19659 5648 19701 5657
rect 19659 5608 19660 5648
rect 19700 5608 19701 5648
rect 19659 5599 19701 5608
rect 19755 5648 19797 5657
rect 19755 5608 19756 5648
rect 19796 5608 19797 5648
rect 19755 5599 19797 5608
rect 17347 5480 17405 5481
rect 17347 5440 17356 5480
rect 17396 5440 17405 5480
rect 17347 5439 17405 5440
rect 19459 5480 19517 5481
rect 19459 5440 19468 5480
rect 19508 5440 19517 5480
rect 19459 5439 19517 5440
rect 1152 5312 20452 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20452 5312
rect 1152 5248 20452 5272
rect 6603 5144 6645 5153
rect 6603 5104 6604 5144
rect 6644 5104 6645 5144
rect 6603 5095 6645 5104
rect 15043 5144 15101 5145
rect 15043 5104 15052 5144
rect 15092 5104 15101 5144
rect 15043 5103 15101 5104
rect 17355 4808 17397 4817
rect 17355 4768 17356 4808
rect 17396 4768 17397 4808
rect 17355 4759 17397 4768
rect 1152 4556 20352 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 20352 4556
rect 1152 4492 20352 4516
rect 6603 4304 6645 4313
rect 6603 4264 6604 4304
rect 6644 4264 6645 4304
rect 6603 4255 6645 4264
rect 15051 4304 15093 4313
rect 15051 4264 15052 4304
rect 15092 4264 15093 4304
rect 15051 4255 15093 4264
rect 17347 3968 17405 3969
rect 17347 3928 17356 3968
rect 17396 3928 17405 3968
rect 17347 3927 17405 3928
rect 1152 3800 20452 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20452 3800
rect 1152 3736 20452 3760
rect 6603 3632 6645 3641
rect 6603 3592 6604 3632
rect 6644 3592 6645 3632
rect 6603 3583 6645 3592
rect 15043 3632 15101 3633
rect 15043 3592 15052 3632
rect 15092 3592 15101 3632
rect 15043 3591 15101 3592
rect 17347 3632 17405 3633
rect 17347 3592 17356 3632
rect 17396 3592 17405 3632
rect 17347 3591 17405 3592
rect 1152 3044 20352 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 20352 3044
rect 1152 2980 20352 3004
rect 6891 2876 6933 2885
rect 6891 2836 6892 2876
rect 6932 2836 6933 2876
rect 6891 2827 6933 2836
rect 15051 2792 15093 2801
rect 15051 2752 15052 2792
rect 15092 2752 15093 2792
rect 15051 2743 15093 2752
rect 7075 2708 7133 2709
rect 7075 2668 7084 2708
rect 7124 2668 7133 2708
rect 7075 2667 7133 2668
rect 11395 2708 11453 2709
rect 11395 2668 11404 2708
rect 11444 2668 11453 2708
rect 11395 2667 11453 2668
rect 13795 2708 13853 2709
rect 13795 2668 13804 2708
rect 13844 2668 13853 2708
rect 13795 2667 13853 2668
rect 14371 2708 14429 2709
rect 14371 2668 14380 2708
rect 14420 2668 14429 2708
rect 14371 2667 14429 2668
rect 11595 2456 11637 2465
rect 11595 2416 11596 2456
rect 11636 2416 11637 2456
rect 11595 2407 11637 2416
rect 13995 2456 14037 2465
rect 13995 2416 13996 2456
rect 14036 2416 14037 2456
rect 13995 2407 14037 2416
rect 14571 2456 14613 2465
rect 14571 2416 14572 2456
rect 14612 2416 14613 2456
rect 14571 2407 14613 2416
rect 1152 2288 20452 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20452 2288
rect 1152 2224 20452 2248
rect 5739 2120 5781 2129
rect 5739 2080 5740 2120
rect 5780 2080 5781 2120
rect 5739 2071 5781 2080
rect 6123 2120 6165 2129
rect 6123 2080 6124 2120
rect 6164 2080 6165 2120
rect 6123 2071 6165 2080
rect 6507 2120 6549 2129
rect 6507 2080 6508 2120
rect 6548 2080 6549 2120
rect 6507 2071 6549 2080
rect 6891 2120 6933 2129
rect 6891 2080 6892 2120
rect 6932 2080 6933 2120
rect 6891 2071 6933 2080
rect 7275 2120 7317 2129
rect 7275 2080 7276 2120
rect 7316 2080 7317 2120
rect 7275 2071 7317 2080
rect 7659 2120 7701 2129
rect 7659 2080 7660 2120
rect 7700 2080 7701 2120
rect 7659 2071 7701 2080
rect 13891 2120 13949 2121
rect 13891 2080 13900 2120
rect 13940 2080 13949 2120
rect 13891 2079 13949 2080
rect 15243 2120 15285 2129
rect 15243 2080 15244 2120
rect 15284 2080 15285 2120
rect 15243 2071 15285 2080
rect 17259 2120 17301 2129
rect 17259 2080 17260 2120
rect 17300 2080 17301 2120
rect 17259 2071 17301 2080
rect 17643 2120 17685 2129
rect 17643 2080 17644 2120
rect 17684 2080 17685 2120
rect 17643 2071 17685 2080
rect 18027 2120 18069 2129
rect 18027 2080 18028 2120
rect 18068 2080 18069 2120
rect 18027 2071 18069 2080
rect 18411 2120 18453 2129
rect 18411 2080 18412 2120
rect 18452 2080 18453 2120
rect 18411 2071 18453 2080
rect 18795 2120 18837 2129
rect 18795 2080 18796 2120
rect 18836 2080 18837 2120
rect 18795 2071 18837 2080
rect 19179 2120 19221 2129
rect 19179 2080 19180 2120
rect 19220 2080 19221 2120
rect 19179 2071 19221 2080
rect 19563 2120 19605 2129
rect 19563 2080 19564 2120
rect 19604 2080 19605 2120
rect 19563 2071 19605 2080
rect 19947 2120 19989 2129
rect 19947 2080 19948 2120
rect 19988 2080 19989 2120
rect 19947 2071 19989 2080
rect 10147 1881 10205 1882
rect 5923 1868 5981 1869
rect 5923 1828 5932 1868
rect 5972 1828 5981 1868
rect 5923 1827 5981 1828
rect 6307 1868 6365 1869
rect 6307 1828 6316 1868
rect 6356 1828 6365 1868
rect 6307 1827 6365 1828
rect 6691 1868 6749 1869
rect 6691 1828 6700 1868
rect 6740 1828 6749 1868
rect 6691 1827 6749 1828
rect 7075 1868 7133 1869
rect 7075 1828 7084 1868
rect 7124 1828 7133 1868
rect 7075 1827 7133 1828
rect 7459 1868 7517 1869
rect 7459 1828 7468 1868
rect 7508 1828 7517 1868
rect 7459 1827 7517 1828
rect 7843 1868 7901 1869
rect 7843 1828 7852 1868
rect 7892 1828 7901 1868
rect 7843 1827 7901 1828
rect 8131 1868 8189 1869
rect 8131 1828 8140 1868
rect 8180 1828 8189 1868
rect 8131 1827 8189 1828
rect 8611 1868 8669 1869
rect 8611 1828 8620 1868
rect 8660 1828 8669 1868
rect 8611 1827 8669 1828
rect 8995 1868 9053 1869
rect 8995 1828 9004 1868
rect 9044 1828 9053 1868
rect 8995 1827 9053 1828
rect 9571 1868 9629 1869
rect 9571 1828 9580 1868
rect 9620 1828 9629 1868
rect 9571 1827 9629 1828
rect 9763 1868 9821 1869
rect 9763 1828 9772 1868
rect 9812 1828 9821 1868
rect 10147 1841 10156 1881
rect 10196 1841 10205 1881
rect 10147 1840 10205 1841
rect 10531 1868 10589 1869
rect 9763 1827 9821 1828
rect 10531 1828 10540 1868
rect 10580 1828 10589 1868
rect 10531 1827 10589 1828
rect 10915 1868 10973 1869
rect 10915 1828 10924 1868
rect 10964 1828 10973 1868
rect 10915 1827 10973 1828
rect 11491 1868 11549 1869
rect 11491 1828 11500 1868
rect 11540 1828 11549 1868
rect 11491 1827 11549 1828
rect 11683 1868 11741 1869
rect 11683 1828 11692 1868
rect 11732 1828 11741 1868
rect 11683 1827 11741 1828
rect 12067 1868 12125 1869
rect 12067 1828 12076 1868
rect 12116 1828 12125 1868
rect 12067 1827 12125 1828
rect 12739 1868 12797 1869
rect 12739 1828 12748 1868
rect 12788 1828 12797 1868
rect 12739 1827 12797 1828
rect 13315 1868 13373 1869
rect 13315 1828 13324 1868
rect 13364 1828 13373 1868
rect 13315 1827 13373 1828
rect 14275 1868 14333 1869
rect 14275 1828 14284 1868
rect 14324 1828 14333 1868
rect 14275 1827 14333 1828
rect 14659 1868 14717 1869
rect 14659 1828 14668 1868
rect 14708 1828 14717 1868
rect 14659 1827 14717 1828
rect 15619 1868 15677 1869
rect 15619 1828 15628 1868
rect 15668 1828 15677 1868
rect 15619 1827 15677 1828
rect 16003 1868 16061 1869
rect 16003 1828 16012 1868
rect 16052 1828 16061 1868
rect 16003 1827 16061 1828
rect 16387 1868 16445 1869
rect 16387 1828 16396 1868
rect 16436 1828 16445 1868
rect 16387 1827 16445 1828
rect 16771 1868 16829 1869
rect 16771 1828 16780 1868
rect 16820 1828 16829 1868
rect 16771 1827 16829 1828
rect 17443 1868 17501 1869
rect 17443 1828 17452 1868
rect 17492 1828 17501 1868
rect 17443 1827 17501 1828
rect 17827 1868 17885 1869
rect 17827 1828 17836 1868
rect 17876 1828 17885 1868
rect 17827 1827 17885 1828
rect 18211 1868 18269 1869
rect 18211 1828 18220 1868
rect 18260 1828 18269 1868
rect 18211 1827 18269 1828
rect 18595 1868 18653 1869
rect 18595 1828 18604 1868
rect 18644 1828 18653 1868
rect 18595 1827 18653 1828
rect 18979 1868 19037 1869
rect 18979 1828 18988 1868
rect 19028 1828 19037 1868
rect 18979 1827 19037 1828
rect 19363 1868 19421 1869
rect 19363 1828 19372 1868
rect 19412 1828 19421 1868
rect 19363 1827 19421 1828
rect 19747 1868 19805 1869
rect 19747 1828 19756 1868
rect 19796 1828 19805 1868
rect 19747 1827 19805 1828
rect 20120 1865 20162 1874
rect 20120 1825 20121 1865
rect 20161 1825 20162 1865
rect 20120 1816 20162 1825
rect 9195 1784 9237 1793
rect 9195 1744 9196 1784
rect 9236 1744 9237 1784
rect 9195 1735 9237 1744
rect 15435 1784 15477 1793
rect 15435 1744 15436 1784
rect 15476 1744 15477 1784
rect 15435 1735 15477 1744
rect 8331 1700 8373 1709
rect 8331 1660 8332 1700
rect 8372 1660 8373 1700
rect 8331 1651 8373 1660
rect 8811 1700 8853 1709
rect 8811 1660 8812 1700
rect 8852 1660 8853 1700
rect 8811 1651 8853 1660
rect 9387 1700 9429 1709
rect 9387 1660 9388 1700
rect 9428 1660 9429 1700
rect 9387 1651 9429 1660
rect 9963 1700 10005 1709
rect 9963 1660 9964 1700
rect 10004 1660 10005 1700
rect 9963 1651 10005 1660
rect 10347 1700 10389 1709
rect 10347 1660 10348 1700
rect 10388 1660 10389 1700
rect 10347 1651 10389 1660
rect 10731 1700 10773 1709
rect 10731 1660 10732 1700
rect 10772 1660 10773 1700
rect 10731 1651 10773 1660
rect 11115 1700 11157 1709
rect 11115 1660 11116 1700
rect 11156 1660 11157 1700
rect 11115 1651 11157 1660
rect 11307 1700 11349 1709
rect 11307 1660 11308 1700
rect 11348 1660 11349 1700
rect 11307 1651 11349 1660
rect 11883 1700 11925 1709
rect 11883 1660 11884 1700
rect 11924 1660 11925 1700
rect 11883 1651 11925 1660
rect 12267 1700 12309 1709
rect 12267 1660 12268 1700
rect 12308 1660 12309 1700
rect 12267 1651 12309 1660
rect 12939 1700 12981 1709
rect 12939 1660 12940 1700
rect 12980 1660 12981 1700
rect 12939 1651 12981 1660
rect 13131 1700 13173 1709
rect 13131 1660 13132 1700
rect 13172 1660 13173 1700
rect 13131 1651 13173 1660
rect 14091 1700 14133 1709
rect 14091 1660 14092 1700
rect 14132 1660 14133 1700
rect 14091 1651 14133 1660
rect 14475 1700 14517 1709
rect 14475 1660 14476 1700
rect 14516 1660 14517 1700
rect 14475 1651 14517 1660
rect 15819 1700 15861 1709
rect 15819 1660 15820 1700
rect 15860 1660 15861 1700
rect 15819 1651 15861 1660
rect 16203 1700 16245 1709
rect 16203 1660 16204 1700
rect 16244 1660 16245 1700
rect 16203 1651 16245 1660
rect 16587 1700 16629 1709
rect 16587 1660 16588 1700
rect 16628 1660 16629 1700
rect 16587 1651 16629 1660
rect 1152 1532 20352 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 20352 1532
rect 1152 1468 20352 1492
rect 6507 1280 6549 1289
rect 6507 1240 6508 1280
rect 6548 1240 6549 1280
rect 6507 1231 6549 1240
rect 14187 1280 14229 1289
rect 14187 1240 14188 1280
rect 14228 1240 14229 1280
rect 14187 1231 14229 1240
rect 18027 1280 18069 1289
rect 18027 1240 18028 1280
rect 18068 1240 18069 1280
rect 18027 1231 18069 1240
rect 18411 1280 18453 1289
rect 18411 1240 18412 1280
rect 18452 1240 18453 1280
rect 18411 1231 18453 1240
rect 18795 1280 18837 1289
rect 18795 1240 18796 1280
rect 18836 1240 18837 1280
rect 18795 1231 18837 1240
rect 6691 1196 6749 1197
rect 6691 1156 6700 1196
rect 6740 1156 6749 1196
rect 6691 1155 6749 1156
rect 6883 1196 6941 1197
rect 6883 1156 6892 1196
rect 6932 1156 6941 1196
rect 6883 1155 6941 1156
rect 9379 1196 9437 1197
rect 9379 1156 9388 1196
rect 9428 1156 9437 1196
rect 9379 1155 9437 1156
rect 10339 1196 10397 1197
rect 10339 1156 10348 1196
rect 10388 1156 10397 1196
rect 10339 1155 10397 1156
rect 11107 1196 11165 1197
rect 11107 1156 11116 1196
rect 11156 1156 11165 1196
rect 11107 1155 11165 1156
rect 11587 1196 11645 1197
rect 11587 1156 11596 1196
rect 11636 1156 11645 1196
rect 11587 1155 11645 1156
rect 13027 1196 13085 1197
rect 13027 1156 13036 1196
rect 13076 1156 13085 1196
rect 13027 1155 13085 1156
rect 13411 1196 13469 1197
rect 13411 1156 13420 1196
rect 13460 1156 13469 1196
rect 13411 1155 13469 1156
rect 13803 1196 13845 1205
rect 13803 1156 13804 1196
rect 13844 1156 13845 1196
rect 13803 1147 13845 1156
rect 14563 1196 14621 1197
rect 14563 1156 14572 1196
rect 14612 1156 14621 1196
rect 14563 1155 14621 1156
rect 14947 1196 15005 1197
rect 14947 1156 14956 1196
rect 14996 1156 15005 1196
rect 14947 1155 15005 1156
rect 15331 1196 15389 1197
rect 15331 1156 15340 1196
rect 15380 1156 15389 1196
rect 15331 1155 15389 1156
rect 15715 1196 15773 1197
rect 15715 1156 15724 1196
rect 15764 1156 15773 1196
rect 15715 1155 15773 1156
rect 16099 1196 16157 1197
rect 16099 1156 16108 1196
rect 16148 1156 16157 1196
rect 16099 1155 16157 1156
rect 18211 1196 18269 1197
rect 18211 1156 18220 1196
rect 18260 1156 18269 1196
rect 18211 1155 18269 1156
rect 18595 1196 18653 1197
rect 18595 1156 18604 1196
rect 18644 1156 18653 1196
rect 18595 1155 18653 1156
rect 18979 1196 19037 1197
rect 18979 1156 18988 1196
rect 19028 1156 19037 1196
rect 18979 1155 19037 1156
rect 19363 1196 19421 1197
rect 19363 1156 19372 1196
rect 19412 1156 19421 1196
rect 19363 1155 19421 1156
rect 7083 944 7125 953
rect 7083 904 7084 944
rect 7124 904 7125 944
rect 7083 895 7125 904
rect 9195 944 9237 953
rect 9195 904 9196 944
rect 9236 904 9237 944
rect 9195 895 9237 904
rect 10539 944 10581 953
rect 10539 904 10540 944
rect 10580 904 10581 944
rect 10539 895 10581 904
rect 11307 944 11349 953
rect 11307 904 11308 944
rect 11348 904 11349 944
rect 11307 895 11349 904
rect 11787 944 11829 953
rect 11787 904 11788 944
rect 11828 904 11829 944
rect 11787 895 11829 904
rect 13227 944 13269 953
rect 13227 904 13228 944
rect 13268 904 13269 944
rect 13227 895 13269 904
rect 13611 944 13653 953
rect 13611 904 13612 944
rect 13652 904 13653 944
rect 13611 895 13653 904
rect 14379 944 14421 953
rect 14379 904 14380 944
rect 14420 904 14421 944
rect 14379 895 14421 904
rect 14763 944 14805 953
rect 14763 904 14764 944
rect 14804 904 14805 944
rect 14763 895 14805 904
rect 15147 944 15189 953
rect 15147 904 15148 944
rect 15188 904 15189 944
rect 15147 895 15189 904
rect 15531 944 15573 953
rect 15531 904 15532 944
rect 15572 904 15573 944
rect 15531 895 15573 904
rect 15915 944 15957 953
rect 15915 904 15916 944
rect 15956 904 15957 944
rect 15915 895 15957 904
rect 19179 944 19221 953
rect 19179 904 19180 944
rect 19220 904 19221 944
rect 19179 895 19221 904
rect 1152 776 20452 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20452 776
rect 1152 712 20452 736
<< via1 >>
rect 3688 84652 3728 84692
rect 3770 84652 3810 84692
rect 3852 84652 3892 84692
rect 3934 84652 3974 84692
rect 4016 84652 4056 84692
rect 18808 84652 18848 84692
rect 18890 84652 18930 84692
rect 18972 84652 19012 84692
rect 19054 84652 19094 84692
rect 19136 84652 19176 84692
rect 4300 84400 4340 84440
rect 4492 84316 4532 84356
rect 4928 83896 4968 83936
rect 5010 83896 5050 83936
rect 5092 83896 5132 83936
rect 5174 83896 5214 83936
rect 5256 83896 5296 83936
rect 20048 83896 20088 83936
rect 20130 83896 20170 83936
rect 20212 83896 20252 83936
rect 20294 83896 20334 83936
rect 20376 83896 20416 83936
rect 1708 83728 1748 83768
rect 1900 83728 1940 83768
rect 2284 83728 2324 83768
rect 2668 83728 2708 83768
rect 3052 83728 3092 83768
rect 3436 83728 3476 83768
rect 3820 83728 3860 83768
rect 4204 83728 4244 83768
rect 4588 83728 4628 83768
rect 4972 83728 5012 83768
rect 5356 83728 5396 83768
rect 5932 83728 5972 83768
rect 6700 83728 6740 83768
rect 7180 83728 7220 83768
rect 7564 83728 7604 83768
rect 7756 83728 7796 83768
rect 8332 83728 8372 83768
rect 8524 83728 8564 83768
rect 13324 83728 13364 83768
rect 14956 83728 14996 83768
rect 15532 83728 15572 83768
rect 15724 83728 15764 83768
rect 18124 83728 18164 83768
rect 19180 83728 19220 83768
rect 19564 83728 19604 83768
rect 1516 83476 1556 83516
rect 2092 83476 2132 83516
rect 2476 83476 2516 83516
rect 2860 83476 2900 83516
rect 3244 83476 3284 83516
rect 3628 83476 3668 83516
rect 4012 83476 4052 83516
rect 4396 83476 4436 83516
rect 4780 83476 4820 83516
rect 5164 83476 5204 83516
rect 5548 83476 5588 83516
rect 6124 83476 6164 83516
rect 6508 83476 6548 83516
rect 6988 83476 7028 83516
rect 7372 83476 7412 83516
rect 7948 83476 7988 83516
rect 8140 83476 8180 83516
rect 8716 83476 8756 83516
rect 13516 83476 13556 83516
rect 15148 83476 15188 83516
rect 15340 83476 15380 83516
rect 15916 83476 15956 83516
rect 18316 83476 18356 83516
rect 18988 83476 19028 83516
rect 19372 83476 19412 83516
rect 3688 83140 3728 83180
rect 3770 83140 3810 83180
rect 3852 83140 3892 83180
rect 3934 83140 3974 83180
rect 4016 83140 4056 83180
rect 18808 83140 18848 83180
rect 18890 83140 18930 83180
rect 18972 83140 19012 83180
rect 19054 83140 19094 83180
rect 19136 83140 19176 83180
rect 2668 82972 2708 83012
rect 3052 82972 3092 83012
rect 3436 82972 3476 83012
rect 3916 82972 3956 83012
rect 4588 82972 4628 83012
rect 19180 82972 19220 83012
rect 19564 82972 19604 83012
rect 2860 82804 2900 82844
rect 3244 82804 3284 82844
rect 3628 82804 3668 82844
rect 4108 82804 4148 82844
rect 4780 82804 4820 82844
rect 18988 82804 19028 82844
rect 19372 82804 19412 82844
rect 4928 82384 4968 82424
rect 5010 82384 5050 82424
rect 5092 82384 5132 82424
rect 5174 82384 5214 82424
rect 5256 82384 5296 82424
rect 20048 82384 20088 82424
rect 20130 82384 20170 82424
rect 20212 82384 20252 82424
rect 20294 82384 20334 82424
rect 20376 82384 20416 82424
rect 14284 82216 14324 82256
rect 15724 82216 15764 82256
rect 14092 81964 14132 82004
rect 15532 81964 15572 82004
rect 3688 81628 3728 81668
rect 3770 81628 3810 81668
rect 3852 81628 3892 81668
rect 3934 81628 3974 81668
rect 4016 81628 4056 81668
rect 18808 81628 18848 81668
rect 18890 81628 18930 81668
rect 18972 81628 19012 81668
rect 19054 81628 19094 81668
rect 19136 81628 19176 81668
rect 19564 81460 19604 81500
rect 19180 81376 19220 81416
rect 18988 81292 19028 81332
rect 19372 81292 19412 81332
rect 4928 80872 4968 80912
rect 5010 80872 5050 80912
rect 5092 80872 5132 80912
rect 5174 80872 5214 80912
rect 5256 80872 5296 80912
rect 20048 80872 20088 80912
rect 20130 80872 20170 80912
rect 20212 80872 20252 80912
rect 20294 80872 20334 80912
rect 20376 80872 20416 80912
rect 13228 80536 13268 80576
rect 14476 80536 14516 80576
rect 18700 80452 18740 80492
rect 19372 80452 19412 80492
rect 19756 80452 19796 80492
rect 18892 80368 18932 80408
rect 19948 80368 19988 80408
rect 14668 80284 14708 80324
rect 19564 80284 19604 80324
rect 3688 80116 3728 80156
rect 3770 80116 3810 80156
rect 3852 80116 3892 80156
rect 3934 80116 3974 80156
rect 4016 80116 4056 80156
rect 18808 80116 18848 80156
rect 18890 80116 18930 80156
rect 18972 80116 19012 80156
rect 19054 80116 19094 80156
rect 19136 80116 19176 80156
rect 15724 79948 15764 79988
rect 15916 79948 15956 79988
rect 16684 79948 16724 79988
rect 19180 79948 19220 79988
rect 15532 79780 15572 79820
rect 16108 79780 16148 79820
rect 16492 79780 16532 79820
rect 18988 79780 19028 79820
rect 19372 79780 19412 79820
rect 19756 79780 19796 79820
rect 11020 79696 11060 79736
rect 12268 79696 12308 79736
rect 13420 79696 13460 79736
rect 14668 79696 14708 79736
rect 10732 79528 10772 79568
rect 12460 79528 12500 79568
rect 14860 79528 14900 79568
rect 19564 79528 19604 79568
rect 19948 79528 19988 79568
rect 4928 79360 4968 79400
rect 5010 79360 5050 79400
rect 5092 79360 5132 79400
rect 5174 79360 5214 79400
rect 5256 79360 5296 79400
rect 20048 79360 20088 79400
rect 20130 79360 20170 79400
rect 20212 79360 20252 79400
rect 20294 79360 20334 79400
rect 20376 79360 20416 79400
rect 19180 79192 19220 79232
rect 10540 79108 10580 79148
rect 12556 79108 12596 79148
rect 14860 79108 14900 79148
rect 9100 79024 9140 79064
rect 10348 79024 10388 79064
rect 10828 79024 10868 79064
rect 10924 79024 10964 79064
rect 11404 79024 11444 79064
rect 11884 79024 11924 79064
rect 12412 79014 12452 79054
rect 13132 79024 13172 79064
rect 13228 79024 13268 79064
rect 13708 79024 13748 79064
rect 14188 79024 14228 79064
rect 14716 79014 14756 79054
rect 15340 79024 15380 79064
rect 16588 79024 16628 79064
rect 11308 78940 11348 78980
rect 13612 78940 13652 78980
rect 18988 78940 19028 78980
rect 19372 78940 19412 78980
rect 19756 78940 19796 78980
rect 16780 78772 16820 78812
rect 19564 78772 19604 78812
rect 19948 78772 19988 78812
rect 3688 78604 3728 78644
rect 3770 78604 3810 78644
rect 3852 78604 3892 78644
rect 3934 78604 3974 78644
rect 4016 78604 4056 78644
rect 18808 78604 18848 78644
rect 18890 78604 18930 78644
rect 18972 78604 19012 78644
rect 19054 78604 19094 78644
rect 19136 78604 19176 78644
rect 13132 78436 13172 78476
rect 18796 78436 18836 78476
rect 19180 78436 19220 78476
rect 8428 78352 8468 78392
rect 19564 78352 19604 78392
rect 18604 78268 18644 78308
rect 18988 78268 19028 78308
rect 19372 78268 19412 78308
rect 19756 78268 19796 78308
rect 11692 78184 11732 78224
rect 12940 78184 12980 78224
rect 14956 78184 14996 78224
rect 15052 78184 15092 78224
rect 15436 78184 15476 78224
rect 16540 78226 16580 78266
rect 15532 78184 15572 78224
rect 16012 78184 16052 78224
rect 10732 78100 10772 78140
rect 16684 78016 16724 78056
rect 19948 78016 19988 78056
rect 4928 77848 4968 77888
rect 5010 77848 5050 77888
rect 5092 77848 5132 77888
rect 5174 77848 5214 77888
rect 5256 77848 5296 77888
rect 20048 77848 20088 77888
rect 20130 77848 20170 77888
rect 20212 77848 20252 77888
rect 20294 77848 20334 77888
rect 20376 77848 20416 77888
rect 8428 77680 8468 77720
rect 16684 77680 16724 77720
rect 17068 77680 17108 77720
rect 8812 77512 8852 77552
rect 10060 77512 10100 77552
rect 10636 77512 10676 77552
rect 11884 77512 11924 77552
rect 13036 77512 13076 77552
rect 14284 77512 14324 77552
rect 15052 77512 15092 77552
rect 16300 77512 16340 77552
rect 17740 77512 17780 77552
rect 18988 77512 19028 77552
rect 16876 77428 16916 77468
rect 17260 77428 17300 77468
rect 19354 77441 19394 77481
rect 19756 77428 19796 77468
rect 10252 77260 10292 77300
rect 12076 77260 12116 77300
rect 14476 77260 14516 77300
rect 16492 77260 16532 77300
rect 19180 77260 19220 77300
rect 19564 77260 19604 77300
rect 19948 77260 19988 77300
rect 3688 77092 3728 77132
rect 3770 77092 3810 77132
rect 3852 77092 3892 77132
rect 3934 77092 3974 77132
rect 4016 77092 4056 77132
rect 18808 77092 18848 77132
rect 18890 77092 18930 77132
rect 18972 77092 19012 77132
rect 19054 77092 19094 77132
rect 19136 77092 19176 77132
rect 8908 76756 8948 76796
rect 10924 76756 10964 76796
rect 6700 76672 6740 76712
rect 7948 76672 7988 76712
rect 8428 76672 8468 76712
rect 8524 76672 8564 76712
rect 9004 76672 9044 76712
rect 9484 76672 9524 76712
rect 9964 76677 10004 76717
rect 10444 76672 10484 76712
rect 10540 76672 10580 76712
rect 12028 76714 12068 76754
rect 15628 76756 15668 76796
rect 18604 76756 18644 76796
rect 18988 76756 19028 76796
rect 19564 76756 19604 76796
rect 19948 76756 19988 76796
rect 11020 76672 11060 76712
rect 11500 76672 11540 76712
rect 13036 76672 13076 76712
rect 13132 76672 13172 76712
rect 13516 76672 13556 76712
rect 13612 76672 13652 76712
rect 14092 76672 14132 76712
rect 14572 76686 14612 76726
rect 15052 76672 15092 76712
rect 15148 76672 15188 76712
rect 15532 76672 15572 76712
rect 16108 76672 16148 76712
rect 16588 76686 16628 76726
rect 17164 76672 17204 76712
rect 18412 76672 18452 76712
rect 8140 76588 8180 76628
rect 10156 76504 10196 76544
rect 12172 76504 12212 76544
rect 14764 76504 14804 76544
rect 16780 76504 16820 76544
rect 16972 76504 17012 76544
rect 18796 76504 18836 76544
rect 19180 76504 19220 76544
rect 19756 76504 19796 76544
rect 20140 76504 20180 76544
rect 4928 76336 4968 76376
rect 5010 76336 5050 76376
rect 5092 76336 5132 76376
rect 5174 76336 5214 76376
rect 5256 76336 5296 76376
rect 20048 76336 20088 76376
rect 20130 76336 20170 76376
rect 20212 76336 20252 76376
rect 20294 76336 20334 76376
rect 20376 76336 20416 76376
rect 8428 76168 8468 76208
rect 10156 76168 10196 76208
rect 14764 76168 14804 76208
rect 15436 76168 15476 76208
rect 19372 76084 19412 76124
rect 6700 76000 6740 76040
rect 7948 76000 7988 76040
rect 8716 76000 8756 76040
rect 9964 76000 10004 76040
rect 11500 76000 11540 76040
rect 12748 76000 12788 76040
rect 13324 76000 13364 76040
rect 14572 76000 14612 76040
rect 15628 76000 15668 76040
rect 16876 76000 16916 76040
rect 17644 76000 17684 76040
rect 17740 76000 17780 76040
rect 18220 76000 18260 76040
rect 18700 76000 18740 76040
rect 19228 75990 19268 76030
rect 15244 75916 15284 75956
rect 18124 75916 18164 75956
rect 19564 75916 19604 75956
rect 19948 75916 19988 75956
rect 10348 75832 10388 75872
rect 12940 75832 12980 75872
rect 17260 75832 17300 75872
rect 8140 75748 8180 75788
rect 17068 75748 17108 75788
rect 19756 75748 19796 75788
rect 20140 75748 20180 75788
rect 3688 75580 3728 75620
rect 3770 75580 3810 75620
rect 3852 75580 3892 75620
rect 3934 75580 3974 75620
rect 4016 75580 4056 75620
rect 18808 75580 18848 75620
rect 18890 75580 18930 75620
rect 18972 75580 19012 75620
rect 19054 75580 19094 75620
rect 19136 75580 19176 75620
rect 8428 75328 8468 75368
rect 18220 75202 18260 75242
rect 6700 75160 6740 75200
rect 7948 75160 7988 75200
rect 9196 75160 9236 75200
rect 10444 75160 10484 75200
rect 10828 75160 10868 75200
rect 12076 75160 12116 75200
rect 13036 75160 13076 75200
rect 14284 75160 14324 75200
rect 15340 75160 15380 75200
rect 16588 75160 16628 75200
rect 16972 75160 17012 75200
rect 18796 75160 18836 75200
rect 20044 75160 20084 75200
rect 8140 74992 8180 75032
rect 8332 74992 8372 75032
rect 10636 74992 10676 75032
rect 12268 74992 12308 75032
rect 14476 74992 14516 75032
rect 16780 74992 16820 75032
rect 18412 74992 18452 75032
rect 18604 74992 18644 75032
rect 4928 74824 4968 74864
rect 5010 74824 5050 74864
rect 5092 74824 5132 74864
rect 5174 74824 5214 74864
rect 5256 74824 5296 74864
rect 20048 74824 20088 74864
rect 20130 74824 20170 74864
rect 20212 74824 20252 74864
rect 20294 74824 20334 74864
rect 20376 74824 20416 74864
rect 10252 74656 10292 74696
rect 14380 74572 14420 74612
rect 16972 74572 17012 74612
rect 19276 74572 19316 74612
rect 5164 74488 5204 74528
rect 6412 74488 6452 74528
rect 6796 74488 6836 74528
rect 8044 74488 8084 74528
rect 8524 74488 8564 74528
rect 8620 74488 8660 74528
rect 9004 74488 9044 74528
rect 9580 74488 9620 74528
rect 10060 74483 10100 74523
rect 10924 74488 10964 74528
rect 12172 74488 12212 74528
rect 12652 74488 12692 74528
rect 12748 74488 12788 74528
rect 13708 74488 13748 74528
rect 14236 74478 14276 74518
rect 15244 74488 15284 74528
rect 15340 74488 15380 74528
rect 15724 74488 15764 74528
rect 16300 74488 16340 74528
rect 16780 74483 16820 74523
rect 17548 74488 17588 74528
rect 17644 74488 17684 74528
rect 18028 74488 18068 74528
rect 18604 74488 18644 74528
rect 19084 74483 19124 74523
rect 9100 74404 9140 74444
rect 13132 74404 13172 74444
rect 13228 74404 13268 74444
rect 15820 74404 15860 74444
rect 18124 74404 18164 74444
rect 19450 74417 19490 74457
rect 19852 74404 19892 74444
rect 6604 74236 6644 74276
rect 8236 74236 8276 74276
rect 12364 74236 12404 74276
rect 19660 74236 19700 74276
rect 20044 74236 20084 74276
rect 3688 74068 3728 74108
rect 3770 74068 3810 74108
rect 3852 74068 3892 74108
rect 3934 74068 3974 74108
rect 4016 74068 4056 74108
rect 18808 74068 18848 74108
rect 18890 74068 18930 74108
rect 18972 74068 19012 74108
rect 19054 74068 19094 74108
rect 19136 74068 19176 74108
rect 14860 73900 14900 73940
rect 19948 73900 19988 73940
rect 5932 73732 5972 73772
rect 9004 73732 9044 73772
rect 11884 73732 11924 73772
rect 11980 73732 12020 73772
rect 18988 73732 19028 73772
rect 19372 73732 19412 73772
rect 19756 73732 19796 73772
rect 3724 73648 3764 73688
rect 4972 73648 5012 73688
rect 5452 73648 5492 73688
rect 5548 73648 5588 73688
rect 6028 73648 6068 73688
rect 6508 73648 6548 73688
rect 6988 73662 7028 73702
rect 8524 73648 8564 73688
rect 8620 73648 8660 73688
rect 9100 73648 9140 73688
rect 9580 73648 9620 73688
rect 10060 73653 10100 73693
rect 11404 73648 11444 73688
rect 11500 73648 11540 73688
rect 12460 73648 12500 73688
rect 12940 73662 12980 73702
rect 13420 73648 13460 73688
rect 14668 73648 14708 73688
rect 15052 73648 15092 73688
rect 16300 73669 16340 73709
rect 17164 73648 17204 73688
rect 18412 73648 18452 73688
rect 5164 73564 5204 73604
rect 13132 73564 13172 73604
rect 7180 73480 7220 73520
rect 10252 73480 10292 73520
rect 16492 73480 16532 73520
rect 18604 73480 18644 73520
rect 19180 73480 19220 73520
rect 19564 73480 19604 73520
rect 4928 73312 4968 73352
rect 5010 73312 5050 73352
rect 5092 73312 5132 73352
rect 5174 73312 5214 73352
rect 5256 73312 5296 73352
rect 20048 73312 20088 73352
rect 20130 73312 20170 73352
rect 20212 73312 20252 73352
rect 20294 73312 20334 73352
rect 20376 73312 20416 73352
rect 18412 73144 18452 73184
rect 8524 73060 8564 73100
rect 13804 73060 13844 73100
rect 3916 72976 3956 73016
rect 5164 72976 5204 73016
rect 7084 72976 7124 73016
rect 8716 72976 8756 73016
rect 9964 72976 10004 73016
rect 10348 72976 10388 73016
rect 11596 72976 11636 73016
rect 12076 72976 12116 73016
rect 8332 72934 8372 72974
rect 12172 72976 12212 73016
rect 13132 72976 13172 73016
rect 13612 72962 13652 73002
rect 14956 72976 14996 73016
rect 16204 72976 16244 73016
rect 16684 72976 16724 73016
rect 16780 72976 16820 73016
rect 17164 72976 17204 73016
rect 17740 72976 17780 73016
rect 18268 72966 18308 73006
rect 12556 72892 12596 72932
rect 12652 72892 12692 72932
rect 17260 72892 17300 72932
rect 18604 72892 18644 72932
rect 18988 72892 19028 72932
rect 19372 72892 19412 72932
rect 19756 72892 19796 72932
rect 10156 72808 10196 72848
rect 18796 72808 18836 72848
rect 19180 72808 19220 72848
rect 5356 72724 5396 72764
rect 11788 72724 11828 72764
rect 16396 72724 16436 72764
rect 19564 72724 19604 72764
rect 19948 72724 19988 72764
rect 3688 72556 3728 72596
rect 3770 72556 3810 72596
rect 3852 72556 3892 72596
rect 3934 72556 3974 72596
rect 4016 72556 4056 72596
rect 18808 72556 18848 72596
rect 18890 72556 18930 72596
rect 18972 72556 19012 72596
rect 19054 72556 19094 72596
rect 19136 72556 19176 72596
rect 19180 72388 19220 72428
rect 1228 72136 1268 72176
rect 2476 72136 2516 72176
rect 4300 72136 4340 72176
rect 5548 72136 5588 72176
rect 5932 72136 5972 72176
rect 7180 72136 7220 72176
rect 7564 72136 7604 72176
rect 8812 72136 8852 72176
rect 10348 72136 10388 72176
rect 11596 72136 11636 72176
rect 11980 72136 12020 72176
rect 13228 72136 13268 72176
rect 13900 72136 13940 72176
rect 15148 72136 15188 72176
rect 16780 72136 16820 72176
rect 17260 72178 17300 72218
rect 18988 72220 19028 72260
rect 19372 72220 19412 72260
rect 19756 72220 19796 72260
rect 17356 72178 17396 72218
rect 16876 72116 16916 72156
rect 17836 72136 17876 72176
rect 18364 72145 18404 72185
rect 2668 71968 2708 72008
rect 5740 71968 5780 72008
rect 7372 71968 7412 72008
rect 9004 71968 9044 72008
rect 11788 71968 11828 72008
rect 13420 71968 13460 72008
rect 15340 71968 15380 72008
rect 18508 71968 18548 72008
rect 19564 71968 19604 72008
rect 19948 71968 19988 72008
rect 4928 71800 4968 71840
rect 5010 71800 5050 71840
rect 5092 71800 5132 71840
rect 5174 71800 5214 71840
rect 5256 71800 5296 71840
rect 20048 71800 20088 71840
rect 20130 71800 20170 71840
rect 20212 71800 20252 71840
rect 20294 71800 20334 71840
rect 20376 71800 20416 71840
rect 8332 71632 8372 71672
rect 15724 71632 15764 71672
rect 6316 71548 6356 71588
rect 10732 71548 10772 71588
rect 13708 71548 13748 71588
rect 1516 71464 1556 71504
rect 2764 71464 2804 71504
rect 4588 71464 4628 71504
rect 4684 71464 4724 71504
rect 5068 71464 5108 71504
rect 5644 71464 5684 71504
rect 6124 71450 6164 71490
rect 6604 71464 6644 71504
rect 6700 71464 6740 71504
rect 7660 71464 7700 71504
rect 8140 71459 8180 71499
rect 9004 71464 9044 71504
rect 9100 71464 9140 71504
rect 10060 71464 10100 71504
rect 10540 71450 10580 71490
rect 11980 71464 12020 71504
rect 12076 71464 12116 71504
rect 13036 71464 13076 71504
rect 13516 71450 13556 71490
rect 13996 71464 14036 71504
rect 14092 71464 14132 71504
rect 14476 71464 14516 71504
rect 15052 71464 15092 71504
rect 15532 71459 15572 71499
rect 15916 71464 15956 71504
rect 17164 71464 17204 71504
rect 17740 71464 17780 71504
rect 18988 71464 19028 71504
rect 5164 71380 5204 71420
rect 7084 71380 7124 71420
rect 7180 71380 7220 71420
rect 8524 71380 8564 71420
rect 9484 71380 9524 71420
rect 9580 71380 9620 71420
rect 12460 71380 12500 71420
rect 12556 71380 12596 71420
rect 14572 71380 14612 71420
rect 19372 71380 19412 71420
rect 19948 71380 19988 71420
rect 2956 71212 2996 71252
rect 8716 71212 8756 71252
rect 17356 71212 17396 71252
rect 19180 71212 19220 71252
rect 19564 71212 19604 71252
rect 20140 71212 20180 71252
rect 3688 71044 3728 71084
rect 3770 71044 3810 71084
rect 3852 71044 3892 71084
rect 3934 71044 3974 71084
rect 4016 71044 4056 71084
rect 18808 71044 18848 71084
rect 18890 71044 18930 71084
rect 18972 71044 19012 71084
rect 19054 71044 19094 71084
rect 19136 71044 19176 71084
rect 5452 70876 5492 70916
rect 8716 70876 8756 70916
rect 13420 70876 13460 70916
rect 19948 70792 19988 70832
rect 9004 70708 9044 70748
rect 19372 70708 19412 70748
rect 19756 70708 19796 70748
rect 2380 70624 2420 70664
rect 3628 70624 3668 70664
rect 4012 70624 4052 70664
rect 5260 70624 5300 70664
rect 5644 70624 5684 70664
rect 6892 70624 6932 70664
rect 7276 70624 7316 70664
rect 8524 70624 8564 70664
rect 10348 70624 10388 70664
rect 11596 70624 11636 70664
rect 11980 70624 12020 70664
rect 13228 70624 13268 70664
rect 13900 70624 13940 70664
rect 15148 70624 15188 70664
rect 16108 70624 16148 70664
rect 17356 70624 17396 70664
rect 17932 70624 17972 70664
rect 19180 70624 19220 70664
rect 17740 70540 17780 70580
rect 3820 70456 3860 70496
rect 7084 70456 7124 70496
rect 11788 70456 11828 70496
rect 15340 70456 15380 70496
rect 17548 70456 17588 70496
rect 19564 70456 19604 70496
rect 4928 70288 4968 70328
rect 5010 70288 5050 70328
rect 5092 70288 5132 70328
rect 5174 70288 5214 70328
rect 5256 70288 5296 70328
rect 20048 70288 20088 70328
rect 20130 70288 20170 70328
rect 20212 70288 20252 70328
rect 20294 70288 20334 70328
rect 20376 70288 20416 70328
rect 11884 70120 11924 70160
rect 17356 70120 17396 70160
rect 9868 70036 9908 70076
rect 4588 69994 4628 70034
rect 19372 70036 19412 70076
rect 1228 69952 1268 69992
rect 2476 69952 2516 69992
rect 2956 69952 2996 69992
rect 4204 69952 4244 69992
rect 5836 69952 5876 69992
rect 6220 69952 6260 69992
rect 7468 69952 7508 69992
rect 8428 69952 8468 69992
rect 9676 69952 9716 69992
rect 10156 69952 10196 69992
rect 10252 69952 10292 69992
rect 11212 69952 11252 69992
rect 11740 69942 11780 69982
rect 13516 69952 13556 69992
rect 14764 69952 14804 69992
rect 15628 69952 15668 69992
rect 15724 69952 15764 69992
rect 16684 69952 16724 69992
rect 17164 69947 17204 69987
rect 17644 69952 17684 69992
rect 17740 69952 17780 69992
rect 18124 69952 18164 69992
rect 18700 69952 18740 69992
rect 19228 69942 19268 69982
rect 10636 69868 10676 69908
rect 10732 69868 10772 69908
rect 16108 69868 16148 69908
rect 16204 69868 16244 69908
rect 18220 69868 18260 69908
rect 19564 69868 19604 69908
rect 19948 69868 19988 69908
rect 2668 69700 2708 69740
rect 4396 69700 4436 69740
rect 6028 69700 6068 69740
rect 7660 69700 7700 69740
rect 14956 69700 14996 69740
rect 19756 69700 19796 69740
rect 20140 69700 20180 69740
rect 3688 69532 3728 69572
rect 3770 69532 3810 69572
rect 3852 69532 3892 69572
rect 3934 69532 3974 69572
rect 4016 69532 4056 69572
rect 18808 69532 18848 69572
rect 18890 69532 18930 69572
rect 18972 69532 19012 69572
rect 19054 69532 19094 69572
rect 19136 69532 19176 69572
rect 11212 69280 11252 69320
rect 17932 69280 17972 69320
rect 17740 69196 17780 69236
rect 19756 69196 19796 69236
rect 2860 69112 2900 69152
rect 2956 69112 2996 69152
rect 3340 69112 3380 69152
rect 3436 69112 3476 69152
rect 3916 69112 3956 69152
rect 4396 69126 4436 69166
rect 4780 69112 4820 69152
rect 6028 69133 6068 69173
rect 6796 69112 6836 69152
rect 6892 69112 6932 69152
rect 7276 69112 7316 69152
rect 7372 69112 7412 69152
rect 7852 69112 7892 69152
rect 8332 69126 8372 69166
rect 8908 69112 8948 69152
rect 10156 69112 10196 69152
rect 10732 69112 10772 69152
rect 11884 69112 11924 69152
rect 13132 69112 13172 69152
rect 13612 69112 13652 69152
rect 13708 69112 13748 69152
rect 14092 69112 14132 69152
rect 14188 69112 14228 69152
rect 14668 69112 14708 69152
rect 15148 69126 15188 69166
rect 16108 69154 16148 69194
rect 17356 69112 17396 69152
rect 18124 69112 18164 69152
rect 19372 69112 19412 69152
rect 8524 69028 8564 69068
rect 13324 69028 13364 69068
rect 15340 69028 15380 69068
rect 4588 68944 4628 68984
rect 6220 68944 6260 68984
rect 10348 68944 10388 68984
rect 17548 68944 17588 68984
rect 19564 68944 19604 68984
rect 19948 68944 19988 68984
rect 4928 68776 4968 68816
rect 5010 68776 5050 68816
rect 5092 68776 5132 68816
rect 5174 68776 5214 68816
rect 5256 68776 5296 68816
rect 20048 68776 20088 68816
rect 20130 68776 20170 68816
rect 20212 68776 20252 68816
rect 20294 68776 20334 68816
rect 20376 68776 20416 68816
rect 12364 68608 12404 68648
rect 19372 68608 19412 68648
rect 5164 68524 5204 68564
rect 8044 68524 8084 68564
rect 1516 68440 1556 68480
rect 2764 68440 2804 68480
rect 3436 68440 3476 68480
rect 3532 68440 3572 68480
rect 4012 68440 4052 68480
rect 4492 68440 4532 68480
rect 4972 68435 5012 68475
rect 6316 68440 6356 68480
rect 6412 68440 6452 68480
rect 7372 68440 7412 68480
rect 7852 68435 7892 68475
rect 8236 68440 8276 68480
rect 9484 68440 9524 68480
rect 10636 68440 10676 68480
rect 10732 68440 10772 68480
rect 11212 68440 11252 68480
rect 11692 68440 11732 68480
rect 12172 68426 12212 68466
rect 14092 68440 14132 68480
rect 15340 68440 15380 68480
rect 15724 68440 15764 68480
rect 16972 68440 17012 68480
rect 17644 68440 17684 68480
rect 17740 68440 17780 68480
rect 18220 68440 18260 68480
rect 18700 68440 18740 68480
rect 19228 68430 19268 68470
rect 3916 68356 3956 68396
rect 6796 68356 6836 68396
rect 6892 68356 6932 68396
rect 11116 68356 11156 68396
rect 18124 68356 18164 68396
rect 19564 68356 19604 68396
rect 19948 68356 19988 68396
rect 2956 68188 2996 68228
rect 9676 68188 9716 68228
rect 15532 68188 15572 68228
rect 17164 68188 17204 68228
rect 19756 68188 19796 68228
rect 20140 68188 20180 68228
rect 3688 68020 3728 68060
rect 3770 68020 3810 68060
rect 3852 68020 3892 68060
rect 3934 68020 3974 68060
rect 4016 68020 4056 68060
rect 18808 68020 18848 68060
rect 18890 68020 18930 68060
rect 18972 68020 19012 68060
rect 19054 68020 19094 68060
rect 19136 68020 19176 68060
rect 11596 67852 11636 67892
rect 15916 67852 15956 67892
rect 10252 67684 10292 67724
rect 15724 67684 15764 67724
rect 19756 67684 19796 67724
rect 1324 67600 1364 67640
rect 2572 67600 2612 67640
rect 2956 67600 2996 67640
rect 4204 67600 4244 67640
rect 4588 67600 4628 67640
rect 5836 67600 5876 67640
rect 6220 67600 6260 67640
rect 7468 67600 7508 67640
rect 7852 67600 7892 67640
rect 9100 67600 9140 67640
rect 9676 67600 9716 67640
rect 9772 67600 9812 67640
rect 11260 67642 11300 67682
rect 10156 67600 10196 67640
rect 10732 67600 10772 67640
rect 11788 67600 11828 67640
rect 13036 67600 13076 67640
rect 13420 67600 13460 67640
rect 14668 67600 14708 67640
rect 16204 67600 16244 67640
rect 16300 67580 16340 67620
rect 16684 67600 16724 67640
rect 16780 67600 16820 67640
rect 17260 67600 17300 67640
rect 17740 67614 17780 67654
rect 18124 67600 18164 67640
rect 19372 67600 19412 67640
rect 11404 67516 11444 67556
rect 17932 67516 17972 67556
rect 2764 67432 2804 67472
rect 4396 67432 4436 67472
rect 6028 67432 6068 67472
rect 7660 67432 7700 67472
rect 9292 67432 9332 67472
rect 14860 67432 14900 67472
rect 19564 67432 19604 67472
rect 19948 67432 19988 67472
rect 4928 67264 4968 67304
rect 5010 67264 5050 67304
rect 5092 67264 5132 67304
rect 5174 67264 5214 67304
rect 5256 67264 5296 67304
rect 20048 67264 20088 67304
rect 20130 67264 20170 67304
rect 20212 67264 20252 67304
rect 20294 67264 20334 67304
rect 20376 67264 20416 67304
rect 9676 67096 9716 67136
rect 11500 67096 11540 67136
rect 15244 67096 15284 67136
rect 19852 67096 19892 67136
rect 20236 67096 20276 67136
rect 13228 67012 13268 67052
rect 1228 66928 1268 66968
rect 2476 66928 2516 66968
rect 3340 66928 3380 66968
rect 4588 66928 4628 66968
rect 4972 66928 5012 66968
rect 6220 66928 6260 66968
rect 7948 66928 7988 66968
rect 8044 66928 8084 66968
rect 8524 66928 8564 66968
rect 9004 66928 9044 66968
rect 9484 66923 9524 66963
rect 10060 66928 10100 66968
rect 11308 66928 11348 66968
rect 11788 66928 11828 66968
rect 13036 66928 13076 66968
rect 13516 66948 13556 66988
rect 13612 66928 13652 66968
rect 13996 66928 14036 66968
rect 14572 66928 14612 66968
rect 15052 66923 15092 66963
rect 16876 66928 16916 66968
rect 17260 66928 17300 66968
rect 18508 66928 18548 66968
rect 8428 66844 8468 66884
rect 15628 66886 15668 66926
rect 14092 66844 14132 66884
rect 19660 66844 19700 66884
rect 20044 66844 20084 66884
rect 4780 66760 4820 66800
rect 6412 66760 6452 66800
rect 2668 66676 2708 66716
rect 17068 66676 17108 66716
rect 18700 66676 18740 66716
rect 3688 66508 3728 66548
rect 3770 66508 3810 66548
rect 3852 66508 3892 66548
rect 3934 66508 3974 66548
rect 4016 66508 4056 66548
rect 18808 66508 18848 66548
rect 18890 66508 18930 66548
rect 18972 66508 19012 66548
rect 19054 66508 19094 66548
rect 19136 66508 19176 66548
rect 17164 66256 17204 66296
rect 19948 66256 19988 66296
rect 4204 66172 4244 66212
rect 6316 66172 6356 66212
rect 6412 66172 6452 66212
rect 18028 66172 18068 66212
rect 19372 66172 19412 66212
rect 19756 66172 19796 66212
rect 1420 66088 1460 66128
rect 2668 66088 2708 66128
rect 3628 66088 3668 66128
rect 3724 66088 3764 66128
rect 4108 66088 4148 66128
rect 4684 66088 4724 66128
rect 5164 66102 5204 66142
rect 5836 66088 5876 66128
rect 5932 66088 5972 66128
rect 6892 66088 6932 66128
rect 7372 66102 7412 66142
rect 9100 66088 9140 66128
rect 10348 66088 10388 66128
rect 10732 66088 10772 66128
rect 11980 66088 12020 66128
rect 12364 66088 12404 66128
rect 13612 66088 13652 66128
rect 13996 66088 14036 66128
rect 15244 66088 15284 66128
rect 17452 66088 17492 66128
rect 17548 66088 17588 66128
rect 17932 66088 17972 66128
rect 18508 66088 18548 66128
rect 19036 66097 19076 66137
rect 7564 66004 7604 66044
rect 2860 65920 2900 65960
rect 5356 65920 5396 65960
rect 10540 65920 10580 65960
rect 12172 65920 12212 65960
rect 13804 65920 13844 65960
rect 15436 65920 15476 65960
rect 19180 65920 19220 65960
rect 19564 65920 19604 65960
rect 4928 65752 4968 65792
rect 5010 65752 5050 65792
rect 5092 65752 5132 65792
rect 5174 65752 5214 65792
rect 5256 65752 5296 65792
rect 20048 65752 20088 65792
rect 20130 65752 20170 65792
rect 20212 65752 20252 65792
rect 20294 65752 20334 65792
rect 20376 65752 20416 65792
rect 16300 65584 16340 65624
rect 4492 65500 4532 65540
rect 12556 65500 12596 65540
rect 15436 65500 15476 65540
rect 18316 65500 18356 65540
rect 2764 65416 2804 65456
rect 2860 65416 2900 65456
rect 3244 65416 3284 65456
rect 3820 65416 3860 65456
rect 3340 65374 3380 65414
rect 4300 65411 4340 65451
rect 5836 65416 5876 65456
rect 7084 65416 7124 65456
rect 7468 65416 7508 65456
rect 8716 65416 8756 65456
rect 9100 65416 9140 65456
rect 10348 65416 10388 65456
rect 10828 65416 10868 65456
rect 10924 65416 10964 65456
rect 11308 65416 11348 65456
rect 11404 65416 11444 65456
rect 11884 65416 11924 65456
rect 12364 65411 12404 65451
rect 13708 65416 13748 65456
rect 13804 65416 13844 65456
rect 14188 65416 14228 65456
rect 14284 65416 14324 65456
rect 14764 65416 14804 65456
rect 15292 65406 15332 65446
rect 16588 65416 16628 65456
rect 16684 65416 16724 65456
rect 17068 65416 17108 65456
rect 17164 65416 17204 65456
rect 17644 65416 17684 65456
rect 18124 65411 18164 65451
rect 18988 65332 19028 65372
rect 19372 65332 19412 65372
rect 19756 65332 19796 65372
rect 19564 65248 19604 65288
rect 19948 65248 19988 65288
rect 7276 65164 7316 65204
rect 8908 65164 8948 65204
rect 10540 65164 10580 65204
rect 19180 65164 19220 65204
rect 3688 64996 3728 65036
rect 3770 64996 3810 65036
rect 3852 64996 3892 65036
rect 3934 64996 3974 65036
rect 4016 64996 4056 65036
rect 18808 64996 18848 65036
rect 18890 64996 18930 65036
rect 18972 64996 19012 65036
rect 19054 64996 19094 65036
rect 19136 64996 19176 65036
rect 19948 64828 19988 64868
rect 8140 64660 8180 64700
rect 10252 64660 10292 64700
rect 10348 64660 10388 64700
rect 19372 64660 19412 64700
rect 19756 64660 19796 64700
rect 2572 64576 2612 64616
rect 3820 64576 3860 64616
rect 4204 64576 4244 64616
rect 5452 64576 5492 64616
rect 5836 64576 5876 64616
rect 7084 64576 7124 64616
rect 7564 64576 7604 64616
rect 7660 64576 7700 64616
rect 8044 64576 8084 64616
rect 8620 64576 8660 64616
rect 9100 64590 9140 64630
rect 9772 64576 9812 64616
rect 9868 64576 9908 64616
rect 10828 64576 10868 64616
rect 11308 64590 11348 64630
rect 12364 64576 12404 64616
rect 13612 64576 13652 64616
rect 13996 64576 14036 64616
rect 15244 64576 15284 64616
rect 15724 64576 15764 64616
rect 16972 64576 17012 64616
rect 17740 64576 17780 64616
rect 18988 64576 19028 64616
rect 5644 64492 5684 64532
rect 11500 64492 11540 64532
rect 4012 64408 4052 64448
rect 7276 64408 7316 64448
rect 9292 64408 9332 64448
rect 13804 64408 13844 64448
rect 15436 64408 15476 64448
rect 17164 64408 17204 64448
rect 19180 64408 19220 64448
rect 19564 64408 19604 64448
rect 4928 64240 4968 64280
rect 5010 64240 5050 64280
rect 5092 64240 5132 64280
rect 5174 64240 5214 64280
rect 5256 64240 5296 64280
rect 20048 64240 20088 64280
rect 20130 64240 20170 64280
rect 20212 64240 20252 64280
rect 20294 64240 20334 64280
rect 20376 64240 20416 64280
rect 19180 64072 19220 64112
rect 19948 64072 19988 64112
rect 5164 63988 5204 64028
rect 8140 63988 8180 64028
rect 12556 63988 12596 64028
rect 15628 63988 15668 64028
rect 1708 63904 1748 63944
rect 2956 63904 2996 63944
rect 3436 63904 3476 63944
rect 3532 63904 3572 63944
rect 4012 63904 4052 63944
rect 4492 63904 4532 63944
rect 4972 63899 5012 63939
rect 6412 63904 6452 63944
rect 6508 63904 6548 63944
rect 7468 63904 7508 63944
rect 7948 63899 7988 63939
rect 9100 63904 9140 63944
rect 10348 63904 10388 63944
rect 10828 63904 10868 63944
rect 10924 63904 10964 63944
rect 11404 63904 11444 63944
rect 11884 63904 11924 63944
rect 12364 63899 12404 63939
rect 13900 63904 13940 63944
rect 13996 63904 14036 63944
rect 14956 63904 14996 63944
rect 15436 63899 15476 63939
rect 17452 63904 17492 63944
rect 17548 63904 17588 63944
rect 18508 63904 18548 63944
rect 19036 63894 19076 63934
rect 3916 63820 3956 63860
rect 6892 63820 6932 63860
rect 6988 63820 7028 63860
rect 11308 63820 11348 63860
rect 14380 63820 14420 63860
rect 14476 63820 14516 63860
rect 17932 63820 17972 63860
rect 18028 63820 18068 63860
rect 19372 63820 19412 63860
rect 19756 63820 19796 63860
rect 10540 63736 10580 63776
rect 19564 63736 19604 63776
rect 3148 63652 3188 63692
rect 3688 63484 3728 63524
rect 3770 63484 3810 63524
rect 3852 63484 3892 63524
rect 3934 63484 3974 63524
rect 4016 63484 4056 63524
rect 18808 63484 18848 63524
rect 18890 63484 18930 63524
rect 18972 63484 19012 63524
rect 19054 63484 19094 63524
rect 19136 63484 19176 63524
rect 10444 63316 10484 63356
rect 8812 63232 8852 63272
rect 17164 63232 17204 63272
rect 19660 63232 19700 63272
rect 3436 63148 3476 63188
rect 19468 63148 19508 63188
rect 2860 63064 2900 63104
rect 2956 63064 2996 63104
rect 3340 63064 3380 63104
rect 3916 63064 3956 63104
rect 4396 63078 4436 63118
rect 5644 63064 5684 63104
rect 6892 63064 6932 63104
rect 7372 63064 7412 63104
rect 8620 63064 8660 63104
rect 9004 63064 9044 63104
rect 10252 63064 10292 63104
rect 10636 63064 10676 63104
rect 11884 63064 11924 63104
rect 13804 63064 13844 63104
rect 15052 63064 15092 63104
rect 15532 63064 15572 63104
rect 16780 63064 16820 63104
rect 17548 63064 17588 63104
rect 17644 63064 17684 63104
rect 18028 63064 18068 63104
rect 18124 63064 18164 63104
rect 18604 63064 18644 63104
rect 19132 63073 19172 63113
rect 4588 62980 4628 63020
rect 7084 62980 7124 63020
rect 16972 62980 17012 63020
rect 19276 62980 19316 63020
rect 12076 62896 12116 62936
rect 15244 62896 15284 62936
rect 17164 62896 17204 62936
rect 4928 62728 4968 62768
rect 5010 62728 5050 62768
rect 5092 62728 5132 62768
rect 5174 62728 5214 62768
rect 5256 62728 5296 62768
rect 20048 62728 20088 62768
rect 20130 62728 20170 62768
rect 20212 62728 20252 62768
rect 20294 62728 20334 62768
rect 20376 62728 20416 62768
rect 9292 62560 9332 62600
rect 16780 62560 16820 62600
rect 19468 62560 19508 62600
rect 19852 62560 19892 62600
rect 20236 62560 20276 62600
rect 15628 62476 15668 62516
rect 1228 62392 1268 62432
rect 2476 62392 2516 62432
rect 2956 62392 2996 62432
rect 4204 62392 4244 62432
rect 4588 62392 4628 62432
rect 5836 62392 5876 62432
rect 7564 62392 7604 62432
rect 7660 62392 7700 62432
rect 8620 62392 8660 62432
rect 9100 62387 9140 62427
rect 10924 62392 10964 62432
rect 12172 62392 12212 62432
rect 13900 62392 13940 62432
rect 13996 62392 14036 62432
rect 14956 62392 14996 62432
rect 15436 62387 15476 62427
rect 18028 62392 18068 62432
rect 19276 62392 19316 62432
rect 8044 62308 8084 62348
rect 8140 62308 8180 62348
rect 14380 62308 14420 62348
rect 14476 62308 14516 62348
rect 16588 62308 16628 62348
rect 19660 62308 19700 62348
rect 20044 62308 20084 62348
rect 2668 62140 2708 62180
rect 4396 62140 4436 62180
rect 6028 62140 6068 62180
rect 12364 62140 12404 62180
rect 3688 61972 3728 62012
rect 3770 61972 3810 62012
rect 3852 61972 3892 62012
rect 3934 61972 3974 62012
rect 4016 61972 4056 62012
rect 18808 61972 18848 62012
rect 18890 61972 18930 62012
rect 18972 61972 19012 62012
rect 19054 61972 19094 62012
rect 19136 61972 19176 62012
rect 13900 61804 13940 61844
rect 10252 61720 10292 61760
rect 18796 61720 18836 61760
rect 19948 61720 19988 61760
rect 3436 61636 3476 61676
rect 11116 61636 11156 61676
rect 18604 61636 18644 61676
rect 18988 61636 19028 61676
rect 19372 61636 19412 61676
rect 19756 61636 19796 61676
rect 2860 61552 2900 61592
rect 2956 61552 2996 61592
rect 3340 61552 3380 61592
rect 3916 61552 3956 61592
rect 4396 61557 4436 61597
rect 5356 61552 5396 61592
rect 6604 61552 6644 61592
rect 7180 61552 7220 61592
rect 8428 61552 8468 61592
rect 8812 61552 8852 61592
rect 10060 61552 10100 61592
rect 10540 61571 10580 61611
rect 10636 61552 10676 61592
rect 11020 61552 11060 61592
rect 11596 61552 11636 61592
rect 12076 61566 12116 61606
rect 12460 61552 12500 61592
rect 13708 61552 13748 61592
rect 14572 61552 14612 61592
rect 15820 61552 15860 61592
rect 16204 61552 16244 61592
rect 17452 61552 17492 61592
rect 12268 61468 12308 61508
rect 4588 61384 4628 61424
rect 6796 61384 6836 61424
rect 8620 61384 8660 61424
rect 16012 61384 16052 61424
rect 17644 61384 17684 61424
rect 19180 61384 19220 61424
rect 19564 61384 19604 61424
rect 4928 61216 4968 61256
rect 5010 61216 5050 61256
rect 5092 61216 5132 61256
rect 5174 61216 5214 61256
rect 5256 61216 5296 61256
rect 20048 61216 20088 61256
rect 20130 61216 20170 61256
rect 20212 61216 20252 61256
rect 20294 61216 20334 61256
rect 20376 61216 20416 61256
rect 2860 61048 2900 61088
rect 8908 61048 8948 61088
rect 12460 61048 12500 61088
rect 17836 61048 17876 61088
rect 19852 61048 19892 61088
rect 4876 60964 4916 61004
rect 1420 60880 1460 60920
rect 2668 60880 2708 60920
rect 3148 60880 3188 60920
rect 3244 60880 3284 60920
rect 3724 60880 3764 60920
rect 4204 60880 4244 60920
rect 4684 60875 4724 60915
rect 5452 60880 5492 60920
rect 6700 60880 6740 60920
rect 7180 60880 7220 60920
rect 7276 60880 7316 60920
rect 8236 60880 8276 60920
rect 8716 60875 8756 60915
rect 9100 60880 9140 60920
rect 10060 60880 10100 60920
rect 10732 60880 10772 60920
rect 10828 60880 10868 60920
rect 11788 60880 11828 60920
rect 12316 60870 12356 60910
rect 13324 60880 13364 60920
rect 14572 60880 14612 60920
rect 16108 60880 16148 60920
rect 16204 60880 16244 60920
rect 17164 60880 17204 60920
rect 17644 60875 17684 60915
rect 18124 60880 18164 60920
rect 18220 60880 18260 60920
rect 19180 60880 19220 60920
rect 19660 60866 19700 60906
rect 3628 60796 3668 60836
rect 7660 60796 7700 60836
rect 7756 60796 7796 60836
rect 11212 60796 11252 60836
rect 11308 60796 11348 60836
rect 16588 60796 16628 60836
rect 16684 60796 16724 60836
rect 18604 60796 18644 60836
rect 18700 60796 18740 60836
rect 20044 60796 20084 60836
rect 6892 60628 6932 60668
rect 14764 60628 14804 60668
rect 20236 60628 20276 60668
rect 3688 60460 3728 60500
rect 3770 60460 3810 60500
rect 3852 60460 3892 60500
rect 3934 60460 3974 60500
rect 4016 60460 4056 60500
rect 18808 60460 18848 60500
rect 18890 60460 18930 60500
rect 18972 60460 19012 60500
rect 19054 60460 19094 60500
rect 19136 60460 19176 60500
rect 2668 60292 2708 60332
rect 10636 60292 10676 60332
rect 17452 60292 17492 60332
rect 19564 60292 19604 60332
rect 6700 60124 6740 60164
rect 13804 60124 13844 60164
rect 19756 60124 19796 60164
rect 1228 60040 1268 60080
rect 2476 60040 2516 60080
rect 3052 60040 3092 60080
rect 4300 60040 4340 60080
rect 6124 60040 6164 60080
rect 6220 60040 6260 60080
rect 6604 60040 6644 60080
rect 7180 60040 7220 60080
rect 7660 60054 7700 60094
rect 9196 60040 9236 60080
rect 10444 60040 10484 60080
rect 11500 60040 11540 60080
rect 12748 60040 12788 60080
rect 13228 60040 13268 60080
rect 13324 60040 13364 60080
rect 13708 60040 13748 60080
rect 14284 60040 14324 60080
rect 14764 60054 14804 60094
rect 15148 60040 15188 60080
rect 15244 60040 15284 60080
rect 15436 60040 15476 60080
rect 16012 60040 16052 60080
rect 17260 60040 17300 60080
rect 18124 60040 18164 60080
rect 19372 60040 19412 60080
rect 12940 59956 12980 59996
rect 14956 59956 14996 59996
rect 4492 59872 4532 59912
rect 7852 59872 7892 59912
rect 15340 59872 15380 59912
rect 19948 59872 19988 59912
rect 4928 59704 4968 59744
rect 5010 59704 5050 59744
rect 5092 59704 5132 59744
rect 5174 59704 5214 59744
rect 5256 59704 5296 59744
rect 20048 59704 20088 59744
rect 20130 59704 20170 59744
rect 20212 59704 20252 59744
rect 20294 59704 20334 59744
rect 20376 59704 20416 59744
rect 11308 59536 11348 59576
rect 15436 59536 15476 59576
rect 16876 59536 16916 59576
rect 19180 59536 19220 59576
rect 19948 59536 19988 59576
rect 4876 59452 4916 59492
rect 9292 59452 9332 59492
rect 3148 59368 3188 59408
rect 3244 59368 3284 59408
rect 3724 59368 3764 59408
rect 4204 59368 4244 59408
rect 4684 59363 4724 59403
rect 6028 59368 6068 59408
rect 7276 59368 7316 59408
rect 7852 59368 7892 59408
rect 9100 59368 9140 59408
rect 9580 59368 9620 59408
rect 9676 59368 9716 59408
rect 10636 59368 10676 59408
rect 11116 59354 11156 59394
rect 13996 59368 14036 59408
rect 15244 59368 15284 59408
rect 15628 59368 15668 59408
rect 15724 59353 15764 59393
rect 15916 59368 15956 59408
rect 16012 59368 16052 59408
rect 16113 59368 16153 59408
rect 17452 59368 17492 59408
rect 17548 59368 17588 59408
rect 17932 59368 17972 59408
rect 18028 59368 18068 59408
rect 18508 59368 18548 59408
rect 19036 59358 19076 59398
rect 3628 59284 3668 59324
rect 10060 59284 10100 59324
rect 10156 59284 10196 59324
rect 16684 59284 16724 59324
rect 19372 59284 19412 59324
rect 19756 59284 19796 59324
rect 2764 59200 2804 59240
rect 7468 59200 7508 59240
rect 17068 59200 17108 59240
rect 19564 59200 19604 59240
rect 15628 59116 15668 59156
rect 3688 58948 3728 58988
rect 3770 58948 3810 58988
rect 3852 58948 3892 58988
rect 3934 58948 3974 58988
rect 4016 58948 4056 58988
rect 18808 58948 18848 58988
rect 18890 58948 18930 58988
rect 18972 58948 19012 58988
rect 19054 58948 19094 58988
rect 19136 58948 19176 58988
rect 15340 58780 15380 58820
rect 19084 58780 19124 58820
rect 19564 58780 19604 58820
rect 19948 58780 19988 58820
rect 3148 58696 3188 58736
rect 5740 58612 5780 58652
rect 5836 58612 5876 58652
rect 12172 58612 12212 58652
rect 12268 58612 12308 58652
rect 19372 58612 19412 58652
rect 19756 58612 19796 58652
rect 1420 58528 1460 58568
rect 2668 58528 2708 58568
rect 3532 58528 3572 58568
rect 4780 58528 4820 58568
rect 5260 58528 5300 58568
rect 5356 58528 5396 58568
rect 6316 58528 6356 58568
rect 6796 58533 6836 58573
rect 7564 58528 7604 58568
rect 7660 58528 7700 58568
rect 8044 58528 8084 58568
rect 8140 58528 8180 58568
rect 8620 58528 8660 58568
rect 9100 58533 9140 58573
rect 9964 58528 10004 58568
rect 11212 58528 11252 58568
rect 11692 58528 11732 58568
rect 11788 58528 11828 58568
rect 12748 58528 12788 58568
rect 13276 58537 13316 58577
rect 13708 58528 13748 58568
rect 14956 58528 14996 58568
rect 15532 58528 15572 58568
rect 16780 58528 16820 58568
rect 16972 58528 17012 58568
rect 17068 58528 17108 58568
rect 17644 58528 17684 58568
rect 18892 58528 18932 58568
rect 4972 58444 5012 58484
rect 6988 58444 7028 58484
rect 9292 58444 9332 58484
rect 11404 58444 11444 58484
rect 13420 58444 13460 58484
rect 2860 58360 2900 58400
rect 15148 58360 15188 58400
rect 17260 58360 17300 58400
rect 4928 58192 4968 58232
rect 5010 58192 5050 58232
rect 5092 58192 5132 58232
rect 5174 58192 5214 58232
rect 5256 58192 5296 58232
rect 20048 58192 20088 58232
rect 20130 58192 20170 58232
rect 20212 58192 20252 58232
rect 20294 58192 20334 58232
rect 20376 58192 20416 58232
rect 4108 58024 4148 58064
rect 6796 58024 6836 58064
rect 9004 58024 9044 58064
rect 13324 58024 13364 58064
rect 11212 57940 11252 57980
rect 15628 57940 15668 57980
rect 17356 57940 17396 57980
rect 1324 57856 1364 57896
rect 2572 57856 2612 57896
rect 3148 57856 3188 57896
rect 3340 57856 3380 57896
rect 3436 57856 3476 57896
rect 3628 57856 3668 57896
rect 3724 57856 3764 57896
rect 3916 57856 3956 57896
rect 4012 57856 4052 57896
rect 4113 57856 4153 57896
rect 5356 57856 5396 57896
rect 6604 57856 6644 57896
rect 7564 57856 7604 57896
rect 8812 57856 8852 57896
rect 11020 57856 11060 57896
rect 11884 57856 11924 57896
rect 13132 57856 13172 57896
rect 13996 57856 14036 57896
rect 15244 57856 15284 57896
rect 15724 57856 15764 57896
rect 15916 57856 15956 57896
rect 17164 57856 17204 57896
rect 17548 57856 17588 57896
rect 9772 57814 9812 57854
rect 17644 57856 17684 57896
rect 17740 57856 17780 57896
rect 17836 57856 17876 57896
rect 18124 57856 18164 57896
rect 18412 57856 18452 57896
rect 18508 57898 18548 57938
rect 18988 57856 19028 57896
rect 19084 57856 19124 57896
rect 19180 57856 19220 57896
rect 19276 57856 19316 57896
rect 19468 57856 19508 57896
rect 19660 57856 19700 57896
rect 19852 57772 19892 57812
rect 3436 57688 3476 57728
rect 20044 57688 20084 57728
rect 2764 57604 2804 57644
rect 15436 57604 15476 57644
rect 19660 57604 19700 57644
rect 18796 57562 18836 57602
rect 3688 57436 3728 57476
rect 3770 57436 3810 57476
rect 3852 57436 3892 57476
rect 3934 57436 3974 57476
rect 4016 57436 4056 57476
rect 18808 57436 18848 57476
rect 18890 57436 18930 57476
rect 18972 57436 19012 57476
rect 19054 57436 19094 57476
rect 19136 57436 19176 57476
rect 2764 57268 2804 57308
rect 7180 57268 7220 57308
rect 17740 57268 17780 57308
rect 19948 57184 19988 57224
rect 3628 57100 3668 57140
rect 10060 57100 10100 57140
rect 10156 57100 10196 57140
rect 18028 57100 18068 57140
rect 1324 57016 1364 57056
rect 2572 57016 2612 57056
rect 3052 57016 3092 57056
rect 3148 57016 3188 57056
rect 3532 57016 3572 57056
rect 4108 57016 4148 57056
rect 4636 57025 4676 57065
rect 4972 57016 5012 57056
rect 5068 57016 5108 57056
rect 6988 57016 7028 57056
rect 7180 57016 7220 57056
rect 7372 57016 7412 57056
rect 7468 57016 7508 57056
rect 7564 57016 7604 57056
rect 7852 57016 7892 57056
rect 9100 57016 9140 57056
rect 9580 57016 9620 57056
rect 9676 57016 9716 57056
rect 10636 57016 10676 57056
rect 11116 57021 11156 57061
rect 11980 57016 12020 57056
rect 13228 57016 13268 57056
rect 13708 57016 13748 57056
rect 13804 57016 13844 57056
rect 14188 57016 14228 57056
rect 14284 57016 14324 57056
rect 14764 57016 14804 57056
rect 15244 57030 15284 57070
rect 16300 57016 16340 57056
rect 17548 57016 17588 57056
rect 17932 57016 17972 57056
rect 18124 57016 18164 57056
rect 18316 57016 18356 57056
rect 19564 57016 19604 57056
rect 19948 57016 19988 57056
rect 20140 57030 20180 57070
rect 20236 57016 20276 57056
rect 4780 56932 4820 56972
rect 9292 56932 9332 56972
rect 11308 56932 11348 56972
rect 13420 56932 13460 56972
rect 19756 56932 19796 56972
rect 5260 56848 5300 56888
rect 7660 56848 7700 56888
rect 15436 56848 15476 56888
rect 17740 56848 17780 56888
rect 4928 56680 4968 56720
rect 5010 56680 5050 56720
rect 5092 56680 5132 56720
rect 5174 56680 5214 56720
rect 5256 56680 5296 56720
rect 20048 56680 20088 56720
rect 20130 56680 20170 56720
rect 20212 56680 20252 56720
rect 20294 56680 20334 56720
rect 20376 56680 20416 56720
rect 3052 56512 3092 56552
rect 4876 56512 4916 56552
rect 5068 56512 5108 56552
rect 11116 56512 11156 56552
rect 16684 56512 16724 56552
rect 17164 56512 17204 56552
rect 17644 56512 17684 56552
rect 19660 56512 19700 56552
rect 7948 56428 7988 56468
rect 13420 56428 13460 56468
rect 15532 56428 15572 56468
rect 1612 56344 1652 56384
rect 2860 56344 2900 56384
rect 3436 56344 3476 56384
rect 4684 56344 4724 56384
rect 5164 56344 5204 56384
rect 5836 56344 5876 56384
rect 7084 56344 7124 56384
rect 7564 56344 7604 56384
rect 7852 56344 7892 56384
rect 8428 56344 8468 56384
rect 8620 56344 8660 56384
rect 8716 56344 8756 56384
rect 8908 56344 8948 56384
rect 9100 56344 9140 56384
rect 9676 56344 9716 56384
rect 10924 56344 10964 56384
rect 11980 56344 12020 56384
rect 13228 56344 13268 56384
rect 13804 56344 13844 56384
rect 13900 56344 13940 56384
rect 14284 56344 14324 56384
rect 14380 56344 14420 56384
rect 14860 56344 14900 56384
rect 15340 56339 15380 56379
rect 16876 56344 16916 56384
rect 16972 56344 17012 56384
rect 17356 56344 17396 56384
rect 17452 56344 17492 56384
rect 17932 56344 17972 56384
rect 18028 56344 18068 56384
rect 18508 56344 18548 56384
rect 18988 56344 19028 56384
rect 19468 56330 19508 56370
rect 19852 56344 19892 56384
rect 20044 56344 20084 56384
rect 20140 56344 20180 56384
rect 16492 56260 16532 56300
rect 18412 56260 18452 56300
rect 7276 56176 7316 56216
rect 8236 56176 8276 56216
rect 8428 56176 8468 56216
rect 8908 56176 8948 56216
rect 19852 56092 19892 56132
rect 3688 55924 3728 55964
rect 3770 55924 3810 55964
rect 3852 55924 3892 55964
rect 3934 55924 3974 55964
rect 4016 55924 4056 55964
rect 18808 55924 18848 55964
rect 18890 55924 18930 55964
rect 18972 55924 19012 55964
rect 19054 55924 19094 55964
rect 19136 55924 19176 55964
rect 5932 55756 5972 55796
rect 17164 55756 17204 55796
rect 19852 55756 19892 55796
rect 2764 55672 2804 55712
rect 10060 55672 10100 55712
rect 10924 55588 10964 55628
rect 1324 55504 1364 55544
rect 2572 55504 2612 55544
rect 3148 55504 3188 55544
rect 3244 55504 3284 55544
rect 3436 55504 3476 55544
rect 3532 55504 3572 55544
rect 3633 55504 3673 55544
rect 3916 55504 3956 55544
rect 4012 55504 4052 55544
rect 4492 55504 4532 55544
rect 5740 55504 5780 55544
rect 6220 55504 6260 55544
rect 6316 55504 6356 55544
rect 6700 55504 6740 55544
rect 6796 55504 6836 55544
rect 7276 55504 7316 55544
rect 7756 55509 7796 55549
rect 8140 55504 8180 55544
rect 8236 55504 8276 55544
rect 8332 55504 8372 55544
rect 8428 55504 8468 55544
rect 8620 55504 8660 55544
rect 9868 55504 9908 55544
rect 10348 55504 10388 55544
rect 10444 55504 10484 55544
rect 10828 55504 10868 55544
rect 11404 55504 11444 55544
rect 11932 55513 11972 55553
rect 13228 55504 13268 55544
rect 14476 55504 14516 55544
rect 15724 55504 15764 55544
rect 16972 55504 17012 55544
rect 17644 55504 17684 55544
rect 17740 55504 17780 55544
rect 18412 55504 18452 55544
rect 19660 55504 19700 55544
rect 7948 55420 7988 55460
rect 12076 55420 12116 55460
rect 3532 55336 3572 55376
rect 4204 55336 4244 55376
rect 14668 55336 14708 55376
rect 17932 55336 17972 55376
rect 4928 55168 4968 55208
rect 5010 55168 5050 55208
rect 5092 55168 5132 55208
rect 5174 55168 5214 55208
rect 5256 55168 5296 55208
rect 20048 55168 20088 55208
rect 20130 55168 20170 55208
rect 20212 55168 20252 55208
rect 20294 55168 20334 55208
rect 20376 55168 20416 55208
rect 2860 55000 2900 55040
rect 3052 55000 3092 55040
rect 6988 55000 7028 55040
rect 7660 55000 7700 55040
rect 11980 55000 12020 55040
rect 16300 55000 16340 55040
rect 17836 55000 17876 55040
rect 18124 55000 18164 55040
rect 18508 55000 18548 55040
rect 1420 54832 1460 54872
rect 2668 54832 2708 54872
rect 3148 54832 3188 54872
rect 3340 54832 3380 54872
rect 4588 54832 4628 54872
rect 5548 54832 5588 54872
rect 6796 54832 6836 54872
rect 7372 54832 7412 54872
rect 7468 54832 7508 54872
rect 8236 54832 8276 54872
rect 9484 54832 9524 54872
rect 10060 54832 10100 54872
rect 10156 54832 10196 54872
rect 10252 54832 10292 54872
rect 10348 54832 10388 54872
rect 10540 54832 10580 54872
rect 11788 54832 11828 54872
rect 12940 54832 12980 54872
rect 14188 54832 14228 54872
rect 14860 54832 14900 54872
rect 16108 54832 16148 54872
rect 16684 54832 16724 54872
rect 16876 54832 16916 54872
rect 16972 54832 17012 54872
rect 17356 54832 17396 54872
rect 17452 54832 17492 54872
rect 17548 54832 17588 54872
rect 17644 54832 17684 54872
rect 17932 54832 17972 54872
rect 18700 54832 18740 54872
rect 19948 54832 19988 54872
rect 4780 54580 4820 54620
rect 9676 54580 9716 54620
rect 14380 54580 14420 54620
rect 16684 54580 16724 54620
rect 18508 54580 18548 54620
rect 3688 54412 3728 54452
rect 3770 54412 3810 54452
rect 3852 54412 3892 54452
rect 3934 54412 3974 54452
rect 4016 54412 4056 54452
rect 18808 54412 18848 54452
rect 18890 54412 18930 54452
rect 18972 54412 19012 54452
rect 19054 54412 19094 54452
rect 19136 54412 19176 54452
rect 15340 54160 15380 54200
rect 3724 54076 3764 54116
rect 17260 54076 17300 54116
rect 19372 54076 19412 54116
rect 1420 53992 1460 54032
rect 2668 53992 2708 54032
rect 3148 53992 3188 54032
rect 3244 53992 3284 54032
rect 3628 53992 3668 54032
rect 4204 53992 4244 54032
rect 4684 54006 4724 54046
rect 5068 53992 5108 54032
rect 5164 53992 5204 54032
rect 5260 53992 5300 54032
rect 5740 53992 5780 54032
rect 6988 53992 7028 54032
rect 7276 53992 7316 54032
rect 8524 53992 8564 54032
rect 9004 53992 9044 54032
rect 9100 53992 9140 54032
rect 9484 53992 9524 54032
rect 9580 53992 9620 54032
rect 10060 53992 10100 54032
rect 10540 53997 10580 54037
rect 10924 53992 10964 54032
rect 11212 53992 11252 54032
rect 12460 53992 12500 54032
rect 12940 54011 12980 54051
rect 13036 53992 13076 54032
rect 13420 53992 13460 54032
rect 13516 53992 13556 54032
rect 13996 53992 14036 54032
rect 14476 54006 14516 54046
rect 15148 53992 15188 54032
rect 15340 53992 15380 54032
rect 15532 53992 15572 54032
rect 15628 53992 15668 54032
rect 15724 53992 15764 54032
rect 16204 53997 16244 54037
rect 16684 53992 16724 54032
rect 17164 53992 17204 54032
rect 17644 53992 17684 54032
rect 17740 53992 17780 54032
rect 18412 54006 18452 54046
rect 18892 53992 18932 54032
rect 19468 53992 19508 54032
rect 19852 53992 19892 54032
rect 19948 53992 19988 54032
rect 2860 53908 2900 53948
rect 8716 53908 8756 53948
rect 14668 53908 14708 53948
rect 16012 53908 16052 53948
rect 4876 53824 4916 53864
rect 5356 53824 5396 53864
rect 5548 53824 5588 53864
rect 10732 53824 10772 53864
rect 11020 53824 11060 53864
rect 12652 53824 12692 53864
rect 15820 53824 15860 53864
rect 18220 53824 18260 53864
rect 4928 53656 4968 53696
rect 5010 53656 5050 53696
rect 5092 53656 5132 53696
rect 5174 53656 5214 53696
rect 5256 53656 5296 53696
rect 20048 53656 20088 53696
rect 20130 53656 20170 53696
rect 20212 53656 20252 53696
rect 20294 53656 20334 53696
rect 20376 53656 20416 53696
rect 3052 53488 3092 53528
rect 5836 53488 5876 53528
rect 8044 53488 8084 53528
rect 8812 53488 8852 53528
rect 12748 53488 12788 53528
rect 15244 53488 15284 53528
rect 20140 53488 20180 53528
rect 6028 53404 6068 53444
rect 14860 53404 14900 53444
rect 1228 53320 1268 53360
rect 2476 53320 2516 53360
rect 2956 53320 2996 53360
rect 3148 53320 3188 53360
rect 3244 53320 3284 53360
rect 4396 53320 4436 53360
rect 5644 53320 5684 53360
rect 6220 53315 6260 53355
rect 6700 53320 6740 53360
rect 7180 53320 7220 53360
rect 7660 53320 7700 53360
rect 7756 53320 7796 53360
rect 8236 53320 8276 53360
rect 8332 53320 8372 53360
rect 8524 53320 8564 53360
rect 8620 53320 8660 53360
rect 9004 53320 9044 53360
rect 10252 53320 10292 53360
rect 10828 53320 10868 53360
rect 10924 53320 10964 53360
rect 11116 53320 11156 53360
rect 11308 53320 11348 53360
rect 12556 53320 12596 53360
rect 13132 53320 13172 53360
rect 13228 53320 13268 53360
rect 13612 53320 13652 53360
rect 13708 53320 13748 53360
rect 14188 53320 14228 53360
rect 14716 53310 14756 53350
rect 15436 53320 15476 53360
rect 16876 53320 16916 53360
rect 16684 53278 16724 53318
rect 16972 53320 17012 53360
rect 17068 53320 17108 53360
rect 17164 53320 17204 53360
rect 17548 53320 17588 53360
rect 17644 53320 17684 53360
rect 17740 53320 17780 53360
rect 17836 53320 17876 53360
rect 18028 53320 18068 53360
rect 19276 53320 19316 53360
rect 19660 53320 19700 53360
rect 19852 53320 19892 53360
rect 19948 53320 19988 53360
rect 20236 53320 20276 53360
rect 7276 53236 7316 53276
rect 19468 53152 19508 53192
rect 2668 53068 2708 53108
rect 10444 53068 10484 53108
rect 11116 53068 11156 53108
rect 19660 53068 19700 53108
rect 3688 52900 3728 52940
rect 3770 52900 3810 52940
rect 3852 52900 3892 52940
rect 3934 52900 3974 52940
rect 4016 52900 4056 52940
rect 18808 52900 18848 52940
rect 18890 52900 18930 52940
rect 18972 52900 19012 52940
rect 19054 52900 19094 52940
rect 19136 52900 19176 52940
rect 11404 52732 11444 52772
rect 16108 52732 16148 52772
rect 18220 52732 18260 52772
rect 3724 52648 3764 52688
rect 12940 52648 12980 52688
rect 17164 52648 17204 52688
rect 11692 52564 11732 52604
rect 1420 52480 1460 52520
rect 2668 52480 2708 52520
rect 3052 52480 3092 52520
rect 3340 52480 3380 52520
rect 3532 52480 3572 52520
rect 3724 52480 3764 52520
rect 3820 52480 3860 52520
rect 4204 52480 4244 52520
rect 5452 52480 5492 52520
rect 5836 52480 5876 52520
rect 6028 52493 6068 52533
rect 6220 52480 6260 52520
rect 6412 52480 6452 52520
rect 6508 52480 6548 52520
rect 6892 52480 6932 52520
rect 8140 52480 8180 52520
rect 8332 52480 8372 52520
rect 9580 52480 9620 52520
rect 10156 52480 10196 52520
rect 10348 52522 10388 52562
rect 16588 52564 16628 52604
rect 10252 52480 10292 52520
rect 10732 52480 10772 52520
rect 10828 52480 10868 52520
rect 10924 52480 10964 52520
rect 11212 52480 11252 52520
rect 11596 52480 11636 52520
rect 11788 52480 11828 52520
rect 12460 52480 12500 52520
rect 12556 52480 12596 52520
rect 12748 52480 12788 52520
rect 12940 52480 12980 52520
rect 13036 52480 13076 52520
rect 13228 52480 13268 52520
rect 13324 52480 13364 52520
rect 13516 52480 13556 52520
rect 13612 52480 13652 52520
rect 13713 52480 13753 52520
rect 14188 52480 14228 52520
rect 14284 52480 14324 52520
rect 14668 52480 14708 52520
rect 15916 52480 15956 52520
rect 16492 52480 16532 52520
rect 16684 52480 16724 52520
rect 16876 52480 16916 52520
rect 17164 52480 17204 52520
rect 17356 52480 17396 52520
rect 17548 52480 17588 52520
rect 17644 52480 17684 52520
rect 17836 52480 17876 52520
rect 18028 52480 18068 52520
rect 18412 52480 18452 52520
rect 19660 52480 19700 52520
rect 19852 52480 19892 52520
rect 19948 52480 19988 52520
rect 20044 52480 20084 52520
rect 20140 52525 20180 52565
rect 5644 52396 5684 52436
rect 6316 52396 6356 52436
rect 17452 52396 17492 52436
rect 2860 52312 2900 52352
rect 3244 52312 3284 52352
rect 5932 52312 5972 52352
rect 6700 52312 6740 52352
rect 9772 52312 9812 52352
rect 10444 52312 10484 52352
rect 10636 52312 10676 52352
rect 11116 52312 11156 52352
rect 12268 52312 12308 52352
rect 13708 52312 13748 52352
rect 17932 52312 17972 52352
rect 4928 52144 4968 52184
rect 5010 52144 5050 52184
rect 5092 52144 5132 52184
rect 5174 52144 5214 52184
rect 5256 52144 5296 52184
rect 20048 52144 20088 52184
rect 20130 52144 20170 52184
rect 20212 52144 20252 52184
rect 20294 52144 20334 52184
rect 20376 52144 20416 52184
rect 3052 51976 3092 52016
rect 5452 51976 5492 52016
rect 6604 51976 6644 52016
rect 12940 51976 12980 52016
rect 15820 51976 15860 52016
rect 17932 51976 17972 52016
rect 1420 51808 1460 51848
rect 2668 51808 2708 51848
rect 3244 51803 3284 51843
rect 3724 51808 3764 51848
rect 4204 51808 4244 51848
rect 4300 51808 4340 51848
rect 4684 51808 4724 51848
rect 4780 51808 4820 51848
rect 5356 51808 5396 51848
rect 5644 51808 5684 51848
rect 5740 51808 5780 51848
rect 5932 51808 5972 51848
rect 6124 51808 6164 51848
rect 6220 51808 6260 51848
rect 6412 51808 6452 51848
rect 6748 51798 6788 51838
rect 7276 51808 7316 51848
rect 7756 51808 7796 51848
rect 8236 51808 8276 51848
rect 8332 51808 8372 51848
rect 9868 51808 9908 51848
rect 11116 51808 11156 51848
rect 11500 51808 11540 51848
rect 12748 51808 12788 51848
rect 13516 51808 13556 51848
rect 14764 51808 14804 51848
rect 15916 51808 15956 51848
rect 16204 51808 16244 51848
rect 16300 51808 16340 51848
rect 16684 51808 16724 51848
rect 17260 51808 17300 51848
rect 17740 51794 17780 51834
rect 18124 51808 18164 51848
rect 18413 51823 18453 51863
rect 18700 51808 18740 51848
rect 19948 51808 19988 51848
rect 7852 51724 7892 51764
rect 16780 51724 16820 51764
rect 2860 51640 2900 51680
rect 5932 51640 5972 51680
rect 6412 51556 6452 51596
rect 11308 51556 11348 51596
rect 13324 51556 13364 51596
rect 18124 51556 18164 51596
rect 20140 51556 20180 51596
rect 3688 51388 3728 51428
rect 3770 51388 3810 51428
rect 3852 51388 3892 51428
rect 3934 51388 3974 51428
rect 4016 51388 4056 51428
rect 18808 51388 18848 51428
rect 18890 51388 18930 51428
rect 18972 51388 19012 51428
rect 19054 51388 19094 51428
rect 19136 51388 19176 51428
rect 6124 51220 6164 51260
rect 12748 51220 12788 51260
rect 3052 51136 3092 51176
rect 18028 51136 18068 51176
rect 3532 51052 3572 51092
rect 8620 51052 8660 51092
rect 14188 51052 14228 51092
rect 19564 51052 19604 51092
rect 1228 50968 1268 51008
rect 2476 50968 2516 51008
rect 3052 50968 3092 51008
rect 3340 50968 3380 51008
rect 3628 50968 3668 51008
rect 3820 50968 3860 51008
rect 3916 50968 3956 51008
rect 4012 50968 4052 51008
rect 4108 50968 4148 51008
rect 4684 50968 4724 51008
rect 5932 50968 5972 51008
rect 6316 50968 6356 51008
rect 7564 50968 7604 51008
rect 8044 50968 8084 51008
rect 8140 50968 8180 51008
rect 8524 50968 8564 51008
rect 9100 50968 9140 51008
rect 9628 50977 9668 51017
rect 11308 50968 11348 51008
rect 12556 50968 12596 51008
rect 13228 50982 13268 51022
rect 13708 50968 13748 51008
rect 14284 50968 14324 51008
rect 14668 50968 14708 51008
rect 14764 50968 14804 51008
rect 15532 50968 15572 51008
rect 16780 50968 16820 51008
rect 17356 50968 17396 51008
rect 17548 50968 17588 51008
rect 17644 50968 17684 51008
rect 18028 50968 18068 51008
rect 18604 50982 18644 51022
rect 19084 50968 19124 51008
rect 19660 50968 19700 51008
rect 20044 50968 20084 51008
rect 20140 50948 20180 50988
rect 7756 50884 7796 50924
rect 13036 50884 13076 50924
rect 18412 50884 18452 50924
rect 2668 50800 2708 50840
rect 2860 50800 2900 50840
rect 9772 50800 9812 50840
rect 16972 50800 17012 50840
rect 17452 50800 17492 50840
rect 17836 50800 17876 50840
rect 4928 50632 4968 50672
rect 5010 50632 5050 50672
rect 5092 50632 5132 50672
rect 5174 50632 5214 50672
rect 5256 50632 5296 50672
rect 20048 50632 20088 50672
rect 20130 50632 20170 50672
rect 20212 50632 20252 50672
rect 20294 50632 20334 50672
rect 20376 50632 20416 50672
rect 16972 50464 17012 50504
rect 7948 50380 7988 50420
rect 12652 50380 12692 50420
rect 18988 50380 19028 50420
rect 19276 50380 19316 50420
rect 2572 50296 2612 50336
rect 3820 50296 3860 50336
rect 4108 50296 4148 50336
rect 4588 50296 4628 50336
rect 5836 50296 5876 50336
rect 6412 50296 6452 50336
rect 7372 50296 7412 50336
rect 7660 50251 7700 50291
rect 7756 50296 7796 50336
rect 7852 50296 7892 50336
rect 8236 50296 8276 50336
rect 9484 50296 9524 50336
rect 11212 50296 11252 50336
rect 12460 50296 12500 50336
rect 13036 50296 13076 50336
rect 14284 50296 14324 50336
rect 15532 50296 15572 50336
rect 16780 50296 16820 50336
rect 17164 50283 17204 50323
rect 17356 50296 17396 50336
rect 17548 50296 17588 50336
rect 18796 50296 18836 50336
rect 19180 50296 19220 50336
rect 19372 50296 19412 50336
rect 19468 50296 19508 50336
rect 19660 50251 19700 50291
rect 19756 50296 19796 50336
rect 19948 50296 19988 50336
rect 19852 50254 19892 50294
rect 20140 50296 20180 50336
rect 20236 50296 20276 50336
rect 2380 50044 2420 50084
rect 4012 50044 4052 50084
rect 6028 50044 6068 50084
rect 9676 50044 9716 50084
rect 12844 50044 12884 50084
rect 17164 50044 17204 50084
rect 3688 49876 3728 49916
rect 3770 49876 3810 49916
rect 3852 49876 3892 49916
rect 3934 49876 3974 49916
rect 4016 49876 4056 49916
rect 18808 49876 18848 49916
rect 18890 49876 18930 49916
rect 18972 49876 19012 49916
rect 19054 49876 19094 49916
rect 19136 49876 19176 49916
rect 7084 49708 7124 49748
rect 7276 49708 7316 49748
rect 8236 49708 8276 49748
rect 15244 49708 15284 49748
rect 16684 49708 16724 49748
rect 18412 49708 18452 49748
rect 3820 49540 3860 49580
rect 3916 49540 3956 49580
rect 10156 49540 10196 49580
rect 13900 49540 13940 49580
rect 2860 49470 2900 49510
rect 3340 49456 3380 49496
rect 4300 49456 4340 49496
rect 4396 49456 4436 49496
rect 4780 49456 4820 49496
rect 4876 49456 4916 49496
rect 4972 49456 5012 49496
rect 5644 49456 5684 49496
rect 6892 49456 6932 49496
rect 7564 49456 7604 49496
rect 7660 49456 7700 49496
rect 7948 49456 7988 49496
rect 8236 49456 8276 49496
rect 8428 49456 8468 49496
rect 9580 49456 9620 49496
rect 9676 49456 9716 49496
rect 10060 49456 10100 49496
rect 10636 49456 10676 49496
rect 11116 49461 11156 49501
rect 12940 49461 12980 49501
rect 13420 49456 13460 49496
rect 13996 49456 14036 49496
rect 14380 49456 14420 49496
rect 14476 49456 14516 49496
rect 15052 49456 15092 49496
rect 15244 49456 15284 49496
rect 15436 49456 15476 49496
rect 15532 49456 15572 49496
rect 15628 49456 15668 49496
rect 15724 49456 15764 49496
rect 16012 49456 16052 49496
rect 16300 49456 16340 49496
rect 16396 49456 16436 49496
rect 16972 49456 17012 49496
rect 18220 49456 18260 49496
rect 18604 49456 18644 49496
rect 19852 49456 19892 49496
rect 2668 49372 2708 49412
rect 11308 49372 11348 49412
rect 4684 49288 4724 49328
rect 12748 49288 12788 49328
rect 18412 49288 18452 49328
rect 20044 49288 20084 49328
rect 4928 49120 4968 49160
rect 5010 49120 5050 49160
rect 5092 49120 5132 49160
rect 5174 49120 5214 49160
rect 5256 49120 5296 49160
rect 20048 49120 20088 49160
rect 20130 49120 20170 49160
rect 20212 49120 20252 49160
rect 20294 49120 20334 49160
rect 20376 49120 20416 49160
rect 3628 48952 3668 48992
rect 9484 48952 9524 48992
rect 13132 48952 13172 48992
rect 17164 48952 17204 48992
rect 17356 48952 17396 48992
rect 17836 48952 17876 48992
rect 7468 48868 7508 48908
rect 11500 48868 11540 48908
rect 15148 48868 15188 48908
rect 1324 48784 1364 48824
rect 2572 48784 2612 48824
rect 3148 48784 3188 48824
rect 3244 48784 3284 48824
rect 3436 48784 3476 48824
rect 3772 48774 3812 48814
rect 4300 48784 4340 48824
rect 4780 48784 4820 48824
rect 4876 48784 4916 48824
rect 5260 48784 5300 48824
rect 5356 48784 5396 48824
rect 5740 48784 5780 48824
rect 5836 48784 5876 48824
rect 6220 48784 6260 48824
rect 6316 48784 6356 48824
rect 6796 48784 6836 48824
rect 7276 48779 7316 48819
rect 7660 48784 7700 48824
rect 7852 48784 7892 48824
rect 8044 48784 8084 48824
rect 9292 48784 9332 48824
rect 9772 48784 9812 48824
rect 9868 48784 9908 48824
rect 10252 48784 10292 48824
rect 10348 48784 10388 48824
rect 10828 48784 10868 48824
rect 11356 48774 11396 48814
rect 11692 48784 11732 48824
rect 12940 48784 12980 48824
rect 13708 48784 13748 48824
rect 14956 48784 14996 48824
rect 15436 48784 15476 48824
rect 15532 48784 15572 48824
rect 16492 48784 16532 48824
rect 16972 48779 17012 48819
rect 17452 48784 17492 48824
rect 17548 48784 17588 48824
rect 17644 48784 17684 48824
rect 18028 48779 18068 48819
rect 18508 48784 18548 48824
rect 18988 48784 19028 48824
rect 19084 48784 19124 48824
rect 19468 48784 19508 48824
rect 19564 48784 19604 48824
rect 19852 48784 19892 48824
rect 20044 48784 20084 48824
rect 20140 48784 20180 48824
rect 15916 48700 15956 48740
rect 16012 48700 16052 48740
rect 3436 48616 3476 48656
rect 7660 48616 7700 48656
rect 2764 48532 2804 48572
rect 19852 48532 19892 48572
rect 3688 48364 3728 48404
rect 3770 48364 3810 48404
rect 3852 48364 3892 48404
rect 3934 48364 3974 48404
rect 4016 48364 4056 48404
rect 18808 48364 18848 48404
rect 18890 48364 18930 48404
rect 18972 48364 19012 48404
rect 19054 48364 19094 48404
rect 19136 48364 19176 48404
rect 3244 48196 3284 48236
rect 11692 48196 11732 48236
rect 16204 48196 16244 48236
rect 18412 48196 18452 48236
rect 20044 48196 20084 48236
rect 6796 48112 6836 48152
rect 13036 48028 13076 48068
rect 13132 48028 13172 48068
rect 1228 47944 1268 47984
rect 2476 47944 2516 47984
rect 2860 47944 2900 47984
rect 3052 47944 3092 47984
rect 3436 47944 3476 47984
rect 4684 47944 4724 47984
rect 5356 47944 5396 47984
rect 6604 47944 6644 47984
rect 6988 47944 7028 47984
rect 7084 47944 7124 47984
rect 7468 47944 7508 47984
rect 7564 47944 7604 47984
rect 7660 47944 7700 47984
rect 7756 47944 7796 47984
rect 8620 47944 8660 47984
rect 9868 47944 9908 47984
rect 10252 47944 10292 47984
rect 11500 47944 11540 47984
rect 12556 47944 12596 47984
rect 12652 47944 12692 47984
rect 13612 47944 13652 47984
rect 14092 47949 14132 47989
rect 14764 47944 14804 47984
rect 16012 47944 16052 47984
rect 16396 47944 16436 47984
rect 16492 47944 16532 47984
rect 16972 47944 17012 47984
rect 18220 47944 18260 47984
rect 18604 47944 18644 47984
rect 19852 47944 19892 47984
rect 14284 47860 14324 47900
rect 2668 47776 2708 47816
rect 2956 47776 2996 47816
rect 7276 47776 7316 47816
rect 10060 47776 10100 47816
rect 16684 47776 16724 47816
rect 4928 47608 4968 47648
rect 5010 47608 5050 47648
rect 5092 47608 5132 47648
rect 5174 47608 5214 47648
rect 5256 47608 5296 47648
rect 20048 47608 20088 47648
rect 20130 47608 20170 47648
rect 20212 47608 20252 47648
rect 20294 47608 20334 47648
rect 20376 47608 20416 47648
rect 6412 47440 6452 47480
rect 12364 47440 12404 47480
rect 13996 47440 14036 47480
rect 16396 47440 16436 47480
rect 2572 47356 2612 47396
rect 10348 47356 10388 47396
rect 2476 47272 2516 47312
rect 2668 47272 2708 47312
rect 2764 47272 2804 47312
rect 2956 47272 2996 47312
rect 4204 47272 4244 47312
rect 4588 47272 4628 47312
rect 4876 47272 4916 47312
rect 6604 47272 6644 47312
rect 6700 47272 6740 47312
rect 6892 47272 6932 47312
rect 8140 47272 8180 47312
rect 8620 47272 8660 47312
rect 8716 47272 8756 47312
rect 9676 47272 9716 47312
rect 10156 47267 10196 47307
rect 10924 47272 10964 47312
rect 12172 47272 12212 47312
rect 12556 47272 12596 47312
rect 13804 47272 13844 47312
rect 14956 47272 14996 47312
rect 16204 47272 16244 47312
rect 16780 47272 16820 47312
rect 18028 47272 18068 47312
rect 18604 47272 18644 47312
rect 19852 47272 19892 47312
rect 9100 47188 9140 47228
rect 9196 47188 9236 47228
rect 8332 47104 8372 47144
rect 4396 47020 4436 47060
rect 4588 47020 4628 47060
rect 18220 47020 18260 47060
rect 20044 47020 20084 47060
rect 3688 46852 3728 46892
rect 3770 46852 3810 46892
rect 3852 46852 3892 46892
rect 3934 46852 3974 46892
rect 4016 46852 4056 46892
rect 18808 46852 18848 46892
rect 18890 46852 18930 46892
rect 18972 46852 19012 46892
rect 19054 46852 19094 46892
rect 19136 46852 19176 46892
rect 3436 46516 3476 46556
rect 10732 46516 10772 46556
rect 1228 46432 1268 46472
rect 2476 46432 2516 46472
rect 2956 46432 2996 46472
rect 3052 46432 3092 46472
rect 3532 46432 3572 46472
rect 4012 46432 4052 46472
rect 4492 46446 4532 46486
rect 4972 46432 5012 46472
rect 5068 46432 5108 46472
rect 5164 46432 5204 46472
rect 6124 46474 6164 46514
rect 6220 46474 6260 46514
rect 6316 46432 6356 46472
rect 6412 46432 6452 46472
rect 6700 46432 6740 46472
rect 7084 46432 7124 46472
rect 7276 46474 7316 46514
rect 13420 46516 13460 46556
rect 19084 46516 19124 46556
rect 7180 46432 7220 46472
rect 7756 46432 7796 46472
rect 7852 46432 7892 46472
rect 8044 46432 8084 46472
rect 8236 46432 8276 46472
rect 8428 46432 8468 46472
rect 9676 46432 9716 46472
rect 10156 46432 10196 46472
rect 10252 46432 10292 46472
rect 10636 46432 10676 46472
rect 11212 46432 11252 46472
rect 11692 46437 11732 46477
rect 12844 46432 12884 46472
rect 12940 46432 12980 46472
rect 13324 46432 13364 46472
rect 13900 46432 13940 46472
rect 14380 46437 14420 46477
rect 15340 46432 15380 46472
rect 16588 46432 16628 46472
rect 16972 46432 17012 46472
rect 17068 46432 17108 46472
rect 17164 46432 17204 46472
rect 18508 46432 18548 46472
rect 18604 46432 18644 46472
rect 18988 46432 19028 46472
rect 19564 46432 19604 46472
rect 20044 46437 20084 46477
rect 2668 46348 2708 46388
rect 9868 46348 9908 46388
rect 14572 46348 14612 46388
rect 20236 46348 20276 46388
rect 4684 46264 4724 46304
rect 4876 46264 4916 46304
rect 6892 46264 6932 46304
rect 7372 46264 7412 46304
rect 7564 46264 7604 46304
rect 8140 46264 8180 46304
rect 11884 46264 11924 46304
rect 16780 46264 16820 46304
rect 17260 46264 17300 46304
rect 6604 46198 6644 46238
rect 4928 46096 4968 46136
rect 5010 46096 5050 46136
rect 5092 46096 5132 46136
rect 5174 46096 5214 46136
rect 5256 46096 5296 46136
rect 20048 46096 20088 46136
rect 20130 46096 20170 46136
rect 20212 46096 20252 46136
rect 20294 46096 20334 46136
rect 20376 46096 20416 46136
rect 2860 45928 2900 45968
rect 12652 45928 12692 45968
rect 14284 45928 14324 45968
rect 14476 45928 14516 45968
rect 3340 45844 3380 45884
rect 7564 45844 7604 45884
rect 17260 45844 17300 45884
rect 1420 45760 1460 45800
rect 2668 45760 2708 45800
rect 3532 45746 3572 45786
rect 4012 45760 4052 45800
rect 4972 45760 5012 45800
rect 5068 45760 5108 45800
rect 5836 45760 5876 45800
rect 5932 45760 5972 45800
rect 6316 45760 6356 45800
rect 6412 45760 6452 45800
rect 6892 45760 6932 45800
rect 7372 45746 7412 45786
rect 7948 45760 7988 45800
rect 9196 45760 9236 45800
rect 9580 45760 9620 45800
rect 10828 45760 10868 45800
rect 11212 45760 11252 45800
rect 12460 45760 12500 45800
rect 12844 45760 12884 45800
rect 14092 45760 14132 45800
rect 14668 45760 14708 45800
rect 14764 45760 14804 45800
rect 15532 45760 15572 45800
rect 15628 45760 15668 45800
rect 16012 45760 16052 45800
rect 16108 45760 16148 45800
rect 16588 45760 16628 45800
rect 17068 45755 17108 45795
rect 17452 45760 17492 45800
rect 17740 45760 17780 45800
rect 17932 45760 17972 45800
rect 18028 45760 18068 45800
rect 18220 45760 18260 45800
rect 18412 45760 18452 45800
rect 19660 45760 19700 45800
rect 4492 45676 4532 45716
rect 4588 45676 4628 45716
rect 11020 45592 11060 45632
rect 17932 45592 17972 45632
rect 9388 45508 9428 45548
rect 17740 45508 17780 45548
rect 19852 45508 19892 45548
rect 3688 45340 3728 45380
rect 3770 45340 3810 45380
rect 3852 45340 3892 45380
rect 3934 45340 3974 45380
rect 4016 45340 4056 45380
rect 18808 45340 18848 45380
rect 18890 45340 18930 45380
rect 18972 45340 19012 45380
rect 19054 45340 19094 45380
rect 19136 45340 19176 45380
rect 3436 45172 3476 45212
rect 6988 45172 7028 45212
rect 4012 45088 4052 45128
rect 4396 45088 4436 45128
rect 1996 44920 2036 44960
rect 3244 44920 3284 44960
rect 3724 44920 3764 44960
rect 3916 44920 3956 44960
rect 4012 44920 4052 44960
rect 4396 44912 4436 44952
rect 4684 44920 4724 44960
rect 4972 44920 5012 44960
rect 5548 44920 5588 44960
rect 6796 44920 6836 44960
rect 7180 44920 7220 44960
rect 7276 44920 7316 44960
rect 7372 44920 7412 44960
rect 7468 44920 7508 44960
rect 7660 44920 7700 44960
rect 7756 44920 7796 44960
rect 7948 44920 7988 44960
rect 8140 44920 8180 44960
rect 8236 44920 8276 44960
rect 8764 44962 8804 45002
rect 9772 45004 9812 45044
rect 9868 45004 9908 45044
rect 13804 45004 13844 45044
rect 13900 45004 13940 45044
rect 18892 45004 18932 45044
rect 18988 45004 19028 45044
rect 9292 44920 9332 44960
rect 10252 44920 10292 44960
rect 10348 44920 10388 44960
rect 11404 44920 11444 44960
rect 12652 44920 12692 44960
rect 13324 44920 13364 44960
rect 13420 44920 13460 44960
rect 14380 44920 14420 44960
rect 14860 44925 14900 44965
rect 15244 44920 15284 44960
rect 15436 44920 15476 44960
rect 16684 44920 16724 44960
rect 17932 44920 17972 44960
rect 18412 44920 18452 44960
rect 18508 44920 18548 44960
rect 19468 44920 19508 44960
rect 19948 44934 19988 44974
rect 8620 44836 8660 44876
rect 4204 44752 4244 44792
rect 4876 44752 4916 44792
rect 7852 44752 7892 44792
rect 12844 44752 12884 44792
rect 15052 44710 15092 44750
rect 15340 44752 15380 44792
rect 16300 44752 16340 44792
rect 18124 44752 18164 44792
rect 20140 44752 20180 44792
rect 4928 44584 4968 44624
rect 5010 44584 5050 44624
rect 5092 44584 5132 44624
rect 5174 44584 5214 44624
rect 5256 44584 5296 44624
rect 20048 44584 20088 44624
rect 20130 44584 20170 44624
rect 20212 44584 20252 44624
rect 20294 44584 20334 44624
rect 20376 44584 20416 44624
rect 4588 44416 4628 44456
rect 6316 44416 6356 44456
rect 8332 44416 8372 44456
rect 13612 44416 13652 44456
rect 16108 44416 16148 44456
rect 10348 44332 10388 44372
rect 19948 44332 19988 44372
rect 3148 44248 3188 44288
rect 4396 44248 4436 44288
rect 4876 44248 4916 44288
rect 6124 44248 6164 44288
rect 6892 44248 6932 44288
rect 8140 44248 8180 44288
rect 8620 44248 8660 44288
rect 8716 44248 8756 44288
rect 9100 44248 9140 44288
rect 9196 44248 9236 44288
rect 9676 44248 9716 44288
rect 10156 44234 10196 44274
rect 11788 44248 11828 44288
rect 11980 44248 12020 44288
rect 13228 44248 13268 44288
rect 13804 44248 13844 44288
rect 13900 44248 13940 44288
rect 14092 44248 14132 44288
rect 14188 44248 14228 44288
rect 14284 44248 14324 44288
rect 14380 44248 14420 44288
rect 14668 44248 14708 44288
rect 15916 44248 15956 44288
rect 16780 44248 16820 44288
rect 17164 44248 17204 44288
rect 17260 44248 17300 44288
rect 17452 44248 17492 44288
rect 18220 44248 18260 44288
rect 18316 44248 18356 44288
rect 18700 44248 18740 44288
rect 18796 44248 18836 44288
rect 19276 44248 19316 44288
rect 19804 44238 19844 44278
rect 13420 44080 13460 44120
rect 16300 44080 16340 44120
rect 16780 44080 16820 44120
rect 11692 43996 11732 44036
rect 16588 43996 16628 44036
rect 3688 43828 3728 43868
rect 3770 43828 3810 43868
rect 3852 43828 3892 43868
rect 3934 43828 3974 43868
rect 4016 43828 4056 43868
rect 18808 43828 18848 43868
rect 18890 43828 18930 43868
rect 18972 43828 19012 43868
rect 19054 43828 19094 43868
rect 19136 43828 19176 43868
rect 6700 43660 6740 43700
rect 8332 43660 8372 43700
rect 10156 43660 10196 43700
rect 16108 43660 16148 43700
rect 18604 43660 18644 43700
rect 5068 43576 5108 43616
rect 3628 43408 3668 43448
rect 4876 43408 4916 43448
rect 5260 43408 5300 43448
rect 6508 43408 6548 43448
rect 6892 43408 6932 43448
rect 8140 43408 8180 43448
rect 8716 43408 8756 43448
rect 9964 43408 10004 43448
rect 11308 43408 11348 43448
rect 12556 43408 12596 43448
rect 13132 43408 13172 43448
rect 13228 43387 13268 43427
rect 13324 43408 13364 43448
rect 13420 43408 13460 43448
rect 13708 43408 13748 43448
rect 14092 43408 14132 43448
rect 14188 43408 14228 43448
rect 14284 43408 14324 43448
rect 14668 43408 14708 43448
rect 15916 43408 15956 43448
rect 16588 43408 16628 43448
rect 16780 43408 16820 43448
rect 16876 43408 16916 43448
rect 17164 43408 17204 43448
rect 18412 43408 18452 43448
rect 12748 43240 12788 43280
rect 13612 43240 13652 43280
rect 13900 43240 13940 43280
rect 14380 43240 14420 43280
rect 16300 43240 16340 43280
rect 16684 43240 16724 43280
rect 18988 43240 19028 43280
rect 4928 43072 4968 43112
rect 5010 43072 5050 43112
rect 5092 43072 5132 43112
rect 5174 43072 5214 43112
rect 5256 43072 5296 43112
rect 20048 43072 20088 43112
rect 20130 43072 20170 43112
rect 20212 43072 20252 43112
rect 20294 43072 20334 43112
rect 20376 43072 20416 43112
rect 16300 42904 16340 42944
rect 4876 42820 4916 42860
rect 9580 42820 9620 42860
rect 1420 42736 1460 42776
rect 2668 42736 2708 42776
rect 3148 42736 3188 42776
rect 3244 42736 3284 42776
rect 4204 42736 4244 42776
rect 4684 42722 4724 42762
rect 5356 42736 5396 42776
rect 6604 42736 6644 42776
rect 6796 42736 6836 42776
rect 8044 42736 8084 42776
rect 10732 42736 10772 42776
rect 11980 42736 12020 42776
rect 12748 42736 12788 42776
rect 13996 42736 14036 42776
rect 14668 42736 14708 42776
rect 15916 42736 15956 42776
rect 3628 42652 3668 42692
rect 3724 42652 3764 42692
rect 9100 42652 9140 42692
rect 20044 42652 20084 42692
rect 16396 42568 16436 42608
rect 17260 42568 17300 42608
rect 18988 42568 19028 42608
rect 19756 42568 19796 42608
rect 20236 42568 20276 42608
rect 2860 42484 2900 42524
rect 5164 42484 5204 42524
rect 8236 42484 8276 42524
rect 12172 42484 12212 42524
rect 14188 42484 14228 42524
rect 16108 42484 16148 42524
rect 3688 42316 3728 42356
rect 3770 42316 3810 42356
rect 3852 42316 3892 42356
rect 3934 42316 3974 42356
rect 4016 42316 4056 42356
rect 18808 42316 18848 42356
rect 18890 42316 18930 42356
rect 18972 42316 19012 42356
rect 19054 42316 19094 42356
rect 19136 42316 19176 42356
rect 3916 42148 3956 42188
rect 18124 42148 18164 42188
rect 9100 42064 9140 42104
rect 19852 42064 19892 42104
rect 4780 41980 4820 42020
rect 10252 41980 10292 42020
rect 12844 41980 12884 42020
rect 14956 41980 14996 42020
rect 17932 41980 17972 42020
rect 19276 41980 19316 42020
rect 19660 41980 19700 42020
rect 2476 41896 2516 41936
rect 3724 41896 3764 41936
rect 4204 41896 4244 41936
rect 4300 41896 4340 41936
rect 4684 41896 4724 41936
rect 5260 41896 5300 41936
rect 5740 41910 5780 41950
rect 7372 41896 7412 41936
rect 8620 41896 8660 41936
rect 9676 41896 9716 41936
rect 9772 41896 9812 41936
rect 10156 41896 10196 41936
rect 10732 41896 10772 41936
rect 11212 41901 11252 41941
rect 12268 41896 12308 41936
rect 12364 41896 12404 41936
rect 12748 41896 12788 41936
rect 13324 41896 13364 41936
rect 13804 41901 13844 41941
rect 14380 41896 14420 41936
rect 14476 41896 14516 41936
rect 15964 41938 16004 41978
rect 14860 41896 14900 41936
rect 15436 41896 15476 41936
rect 16492 41896 16532 41936
rect 17740 41896 17780 41936
rect 18988 41896 19028 41936
rect 8812 41812 8852 41852
rect 5932 41728 5972 41768
rect 11404 41728 11444 41768
rect 13996 41728 14036 41768
rect 16108 41728 16148 41768
rect 16300 41728 16340 41768
rect 19468 41728 19508 41768
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 3244 41392 3284 41432
rect 11788 41392 11828 41432
rect 13420 41392 13460 41432
rect 16396 41392 16436 41432
rect 18988 41392 19028 41432
rect 19852 41392 19892 41432
rect 5452 41308 5492 41348
rect 8236 41308 8276 41348
rect 10252 41308 10292 41348
rect 16108 41308 16148 41348
rect 1804 41224 1844 41264
rect 3052 41224 3092 41264
rect 3724 41224 3764 41264
rect 3820 41224 3860 41264
rect 4300 41224 4340 41264
rect 4780 41224 4820 41264
rect 5308 41214 5348 41254
rect 6796 41224 6836 41264
rect 8044 41224 8084 41264
rect 8524 41224 8564 41264
rect 8620 41224 8660 41264
rect 9580 41224 9620 41264
rect 10060 41219 10100 41259
rect 11980 41224 12020 41264
rect 13228 41224 13268 41264
rect 14380 41224 14420 41264
rect 14476 41224 14516 41264
rect 14956 41224 14996 41264
rect 15436 41224 15476 41264
rect 15964 41214 16004 41254
rect 4204 41140 4244 41180
rect 9004 41140 9044 41180
rect 9100 41140 9140 41180
rect 14860 41140 14900 41180
rect 19276 41140 19316 41180
rect 19660 41140 19700 41180
rect 17260 41056 17300 41096
rect 19468 41056 19508 41096
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 8236 40636 8276 40676
rect 14092 40636 14132 40676
rect 19564 40636 19604 40676
rect 3340 40552 3380 40592
rect 16396 40552 16436 40592
rect 18028 40552 18068 40592
rect 14956 40468 14996 40508
rect 17836 40468 17876 40508
rect 18988 40468 19028 40508
rect 19372 40468 19412 40508
rect 1900 40384 1940 40424
rect 3148 40384 3188 40424
rect 3532 40384 3572 40424
rect 4780 40384 4820 40424
rect 5164 40384 5204 40424
rect 6412 40384 6452 40424
rect 6796 40384 6836 40424
rect 8044 40384 8084 40424
rect 10732 40384 10772 40424
rect 11980 40384 12020 40424
rect 12652 40384 12692 40424
rect 13900 40384 13940 40424
rect 14380 40384 14420 40424
rect 14476 40384 14516 40424
rect 14860 40384 14900 40424
rect 15436 40384 15476 40424
rect 15916 40389 15956 40429
rect 4972 40300 5012 40340
rect 6604 40300 6644 40340
rect 8428 40216 8468 40256
rect 9100 40216 9140 40256
rect 12172 40216 12212 40256
rect 16108 40216 16148 40256
rect 17260 40216 17300 40256
rect 19180 40216 19220 40256
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 2668 39880 2708 39920
rect 9100 39880 9140 39920
rect 14668 39880 14708 39920
rect 16396 39880 16436 39920
rect 17260 39880 17300 39920
rect 18988 39880 19028 39920
rect 5548 39796 5588 39836
rect 8140 39796 8180 39836
rect 11116 39796 11156 39836
rect 14188 39796 14228 39836
rect 1228 39712 1268 39752
rect 2476 39712 2516 39752
rect 3820 39712 3860 39752
rect 3916 39712 3956 39752
rect 4396 39712 4436 39752
rect 4876 39712 4916 39752
rect 5356 39707 5396 39747
rect 6412 39712 6452 39752
rect 6508 39712 6548 39752
rect 6892 39712 6932 39752
rect 7468 39712 7508 39752
rect 7948 39698 7988 39738
rect 9388 39712 9428 39752
rect 9484 39712 9524 39752
rect 9964 39712 10004 39752
rect 10444 39712 10484 39752
rect 10924 39698 10964 39738
rect 12460 39712 12500 39752
rect 12556 39712 12596 39752
rect 13036 39712 13076 39752
rect 13516 39712 13556 39752
rect 13996 39698 14036 39738
rect 14860 39712 14900 39752
rect 16108 39712 16148 39752
rect 4300 39628 4340 39668
rect 6988 39628 7028 39668
rect 9868 39628 9908 39668
rect 12940 39628 12980 39668
rect 19276 39628 19316 39668
rect 19660 39628 19700 39668
rect 9004 39544 9044 39584
rect 16300 39544 16340 39584
rect 17356 39544 17396 39584
rect 19852 39544 19892 39584
rect 19468 39460 19508 39500
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 7180 39040 7220 39080
rect 8812 39040 8852 39080
rect 12460 39040 12500 39080
rect 16300 39040 16340 39080
rect 17260 39040 17300 39080
rect 19852 39040 19892 39080
rect 3052 38956 3092 38996
rect 14956 38956 14996 38996
rect 19276 38956 19316 38996
rect 19660 38956 19700 38996
rect 20044 38956 20084 38996
rect 2476 38872 2516 38912
rect 2572 38872 2612 38912
rect 2956 38872 2996 38912
rect 3532 38872 3572 38912
rect 4012 38877 4052 38917
rect 5740 38872 5780 38912
rect 6988 38872 7028 38912
rect 7372 38872 7412 38912
rect 8620 38872 8660 38912
rect 9004 38872 9044 38912
rect 10252 38872 10292 38912
rect 11020 38872 11060 38912
rect 12268 38872 12308 38912
rect 12652 38872 12692 38912
rect 13900 38872 13940 38912
rect 14380 38872 14420 38912
rect 14476 38872 14516 38912
rect 14860 38872 14900 38912
rect 15436 38872 15476 38912
rect 15964 38881 16004 38921
rect 17452 38872 17492 38912
rect 18700 38872 18740 38912
rect 4204 38788 4244 38828
rect 14092 38788 14132 38828
rect 16108 38788 16148 38828
rect 10444 38704 10484 38744
rect 18988 38704 19028 38744
rect 19468 38704 19508 38744
rect 20236 38704 20276 38744
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 2668 38368 2708 38408
rect 4684 38368 4724 38408
rect 9004 38368 9044 38408
rect 16108 38368 16148 38408
rect 16396 38368 16436 38408
rect 17260 38368 17300 38408
rect 18988 38368 19028 38408
rect 19468 38368 19508 38408
rect 7948 38284 7988 38324
rect 11884 38284 11924 38324
rect 13996 38284 14036 38324
rect 1228 38200 1268 38240
rect 2476 38200 2516 38240
rect 2956 38200 2996 38240
rect 3052 38200 3092 38240
rect 3436 38200 3476 38240
rect 3532 38200 3572 38240
rect 4012 38200 4052 38240
rect 4492 38186 4532 38226
rect 6220 38200 6260 38240
rect 6316 38200 6356 38240
rect 6700 38200 6740 38240
rect 6796 38200 6836 38240
rect 7276 38200 7316 38240
rect 7756 38186 7796 38226
rect 8140 38200 8180 38240
rect 8332 38200 8372 38240
rect 9676 38200 9716 38240
rect 9868 38200 9908 38240
rect 10156 38200 10196 38240
rect 10252 38200 10292 38240
rect 11212 38200 11252 38240
rect 11692 38195 11732 38235
rect 12268 38200 12308 38240
rect 12364 38200 12404 38240
rect 13324 38200 13364 38240
rect 13804 38186 13844 38226
rect 14668 38200 14708 38240
rect 15916 38200 15956 38240
rect 10636 38116 10676 38156
rect 10732 38116 10772 38156
rect 12748 38116 12788 38156
rect 12844 38116 12884 38156
rect 18604 38116 18644 38156
rect 19276 38116 19316 38156
rect 19660 38116 19700 38156
rect 20044 38116 20084 38156
rect 19084 38032 19124 38072
rect 20236 38032 20276 38072
rect 8140 37948 8180 37988
rect 9772 37948 9812 37988
rect 18796 37948 18836 37988
rect 19852 37948 19892 37988
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 3916 37612 3956 37652
rect 5548 37612 5588 37652
rect 7180 37612 7220 37652
rect 8812 37612 8852 37652
rect 12076 37612 12116 37652
rect 13708 37612 13748 37652
rect 10156 37528 10196 37568
rect 19084 37528 19124 37568
rect 15820 37444 15860 37484
rect 15916 37444 15956 37484
rect 19276 37444 19316 37484
rect 19660 37444 19700 37484
rect 20044 37444 20084 37484
rect 2476 37360 2516 37400
rect 3724 37360 3764 37400
rect 4108 37360 4148 37400
rect 5356 37360 5396 37400
rect 5740 37360 5780 37400
rect 6988 37360 7028 37400
rect 7372 37360 7412 37400
rect 8620 37360 8660 37400
rect 9388 37360 9428 37400
rect 9580 37360 9620 37400
rect 9676 37360 9716 37400
rect 10636 37360 10676 37400
rect 11884 37360 11924 37400
rect 12268 37360 12308 37400
rect 13516 37360 13556 37400
rect 15340 37360 15380 37400
rect 15436 37360 15476 37400
rect 16396 37360 16436 37400
rect 16924 37369 16964 37409
rect 17068 37276 17108 37316
rect 9004 37192 9044 37232
rect 9388 37192 9428 37232
rect 10060 37192 10100 37232
rect 17260 37192 17300 37232
rect 19468 37192 19508 37232
rect 19852 37192 19892 37232
rect 20236 37192 20276 37232
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 2668 36856 2708 36896
rect 9580 36856 9620 36896
rect 19084 36856 19124 36896
rect 12940 36772 12980 36812
rect 14956 36772 14996 36812
rect 16972 36772 17012 36812
rect 1228 36688 1268 36728
rect 2476 36688 2516 36728
rect 3340 36688 3380 36728
rect 4588 36688 4628 36728
rect 5548 36688 5588 36728
rect 6796 36688 6836 36728
rect 7372 36688 7412 36728
rect 8620 36688 8660 36728
rect 9772 36688 9812 36728
rect 9868 36688 9908 36728
rect 10636 36688 10676 36728
rect 10924 36688 10964 36728
rect 11020 36688 11060 36728
rect 11500 36688 11540 36728
rect 12748 36688 12788 36728
rect 13228 36688 13268 36728
rect 13324 36688 13364 36728
rect 14284 36688 14324 36728
rect 14764 36674 14804 36714
rect 15244 36688 15284 36728
rect 15340 36688 15380 36728
rect 15724 36688 15764 36728
rect 15820 36688 15860 36728
rect 16300 36688 16340 36728
rect 16780 36674 16820 36714
rect 13708 36604 13748 36644
rect 13804 36604 13844 36644
rect 6988 36520 7028 36560
rect 8812 36520 8852 36560
rect 9004 36520 9044 36560
rect 10060 36520 10100 36560
rect 17260 36520 17300 36560
rect 4780 36436 4820 36476
rect 11308 36436 11348 36476
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 2668 36100 2708 36140
rect 7180 36100 7220 36140
rect 14284 36100 14324 36140
rect 15148 36100 15188 36140
rect 19756 36100 19796 36140
rect 20140 36100 20180 36140
rect 8812 36016 8852 36056
rect 10060 36016 10100 36056
rect 1228 35848 1268 35888
rect 2476 35848 2516 35888
rect 2956 35848 2996 35888
rect 3052 35848 3092 35888
rect 3436 35848 3476 35888
rect 4540 35890 4580 35930
rect 18124 35932 18164 35972
rect 19564 35932 19604 35972
rect 19948 35932 19988 35972
rect 3532 35848 3572 35888
rect 4012 35848 4052 35888
rect 5260 35848 5300 35888
rect 6508 35848 6548 35888
rect 6892 35848 6932 35888
rect 6988 35848 7028 35888
rect 7180 35848 7220 35888
rect 7372 35848 7412 35888
rect 8620 35848 8660 35888
rect 9388 35848 9428 35888
rect 9676 35848 9716 35888
rect 10540 35848 10580 35888
rect 11788 35848 11828 35888
rect 11980 35848 12020 35888
rect 12172 35848 12212 35888
rect 12460 35848 12500 35888
rect 12652 35837 12692 35877
rect 12844 35848 12884 35888
rect 14092 35848 14132 35888
rect 15340 35848 15380 35888
rect 16588 35848 16628 35888
rect 17644 35848 17684 35888
rect 17740 35848 17780 35888
rect 18220 35848 18260 35888
rect 18700 35848 18740 35888
rect 19180 35853 19220 35893
rect 9772 35764 9812 35804
rect 4684 35680 4724 35720
rect 6700 35680 6740 35720
rect 9004 35680 9044 35720
rect 10348 35680 10388 35720
rect 12076 35680 12116 35720
rect 12556 35680 12596 35720
rect 17260 35680 17300 35720
rect 19372 35680 19412 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 4300 35260 4340 35300
rect 7564 35260 7604 35300
rect 8236 35260 8276 35300
rect 9772 35260 9812 35300
rect 14572 35260 14612 35300
rect 16396 35260 16436 35300
rect 17548 35260 17588 35300
rect 2572 35176 2612 35216
rect 2668 35176 2708 35216
rect 3628 35176 3668 35216
rect 4108 35162 4148 35202
rect 4780 35176 4820 35216
rect 5068 35176 5108 35216
rect 5260 35176 5300 35216
rect 5452 35176 5492 35216
rect 5548 35176 5588 35216
rect 5836 35176 5876 35216
rect 5932 35176 5972 35216
rect 6892 35176 6932 35216
rect 2092 35092 2132 35132
rect 3052 35092 3092 35132
rect 3148 35092 3188 35132
rect 6316 35134 6356 35174
rect 7372 35171 7412 35211
rect 7852 35176 7892 35216
rect 8140 35176 8180 35216
rect 9388 35176 9428 35216
rect 9676 35176 9716 35216
rect 10252 35176 10292 35216
rect 10348 35176 10388 35216
rect 10540 35176 10580 35216
rect 11788 35176 11828 35216
rect 12172 35176 12212 35216
rect 12364 35176 12404 35216
rect 12460 35176 12500 35216
rect 13132 35176 13172 35216
rect 14380 35176 14420 35216
rect 14956 35176 14996 35216
rect 16204 35176 16244 35216
rect 17740 35176 17780 35216
rect 18988 35176 19028 35216
rect 6412 35092 6452 35132
rect 19468 35092 19508 35132
rect 19852 35092 19892 35132
rect 5260 35008 5300 35048
rect 9004 35008 9044 35048
rect 12844 35008 12884 35048
rect 17260 35008 17300 35048
rect 19660 35008 19700 35048
rect 20044 35008 20084 35048
rect 1900 34924 1940 34964
rect 5068 34924 5108 34964
rect 8524 34924 8564 34964
rect 10060 34924 10100 34964
rect 11980 34924 12020 34964
rect 12172 34924 12212 34964
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 2668 34588 2708 34628
rect 5932 34588 5972 34628
rect 16876 34588 16916 34628
rect 19660 34588 19700 34628
rect 9964 34504 10004 34544
rect 8332 34420 8372 34460
rect 15052 34420 15092 34460
rect 16684 34420 16724 34460
rect 19468 34420 19508 34460
rect 19852 34420 19892 34460
rect 1228 34336 1268 34376
rect 2476 34336 2516 34376
rect 3052 34336 3092 34376
rect 4300 34336 4340 34376
rect 4492 34336 4532 34376
rect 5740 34336 5780 34376
rect 6124 34336 6164 34376
rect 7372 34336 7412 34376
rect 7756 34336 7796 34376
rect 8044 34336 8084 34376
rect 8524 34336 8564 34376
rect 9772 34336 9812 34376
rect 10252 34336 10292 34376
rect 10348 34336 10388 34376
rect 10732 34336 10772 34376
rect 10828 34336 10868 34376
rect 11308 34336 11348 34376
rect 11788 34341 11828 34381
rect 12172 34336 12212 34376
rect 12268 34336 12308 34376
rect 12460 34336 12500 34376
rect 12748 34336 12788 34376
rect 13996 34336 14036 34376
rect 14476 34336 14516 34376
rect 14572 34336 14612 34376
rect 14956 34336 14996 34376
rect 15532 34336 15572 34376
rect 16012 34341 16052 34381
rect 17548 34336 17588 34376
rect 17644 34336 17684 34376
rect 18028 34336 18068 34376
rect 18124 34336 18164 34376
rect 18604 34336 18644 34376
rect 19132 34345 19172 34385
rect 11980 34252 12020 34292
rect 14188 34252 14228 34292
rect 2860 34168 2900 34208
rect 5932 34168 5972 34208
rect 7564 34168 7604 34208
rect 7948 34168 7988 34208
rect 12364 34168 12404 34208
rect 16204 34168 16244 34208
rect 19276 34168 19316 34208
rect 20044 34168 20084 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 2860 33832 2900 33872
rect 3244 33832 3284 33872
rect 5260 33832 5300 33872
rect 9772 33832 9812 33872
rect 15916 33832 15956 33872
rect 18604 33832 18644 33872
rect 19564 33832 19604 33872
rect 19948 33832 19988 33872
rect 7564 33748 7604 33788
rect 1228 33664 1268 33704
rect 2476 33664 2516 33704
rect 2956 33664 2996 33704
rect 3436 33659 3476 33699
rect 3916 33664 3956 33704
rect 4876 33664 4916 33704
rect 4972 33664 5012 33704
rect 5356 33664 5396 33704
rect 5452 33664 5492 33704
rect 5548 33664 5588 33704
rect 5836 33664 5876 33704
rect 5932 33664 5972 33704
rect 6892 33664 6932 33704
rect 7420 33654 7460 33694
rect 7756 33664 7796 33704
rect 9004 33664 9044 33704
rect 9484 33664 9524 33704
rect 9580 33664 9620 33704
rect 10828 33664 10868 33704
rect 12076 33664 12116 33704
rect 14092 33664 14132 33704
rect 14476 33664 14516 33704
rect 15724 33664 15764 33704
rect 17164 33664 17204 33704
rect 18412 33664 18452 33704
rect 4396 33580 4436 33620
rect 4492 33580 4532 33620
rect 6316 33580 6356 33620
rect 12844 33622 12884 33662
rect 6412 33580 6452 33620
rect 12460 33580 12500 33620
rect 19383 33593 19423 33633
rect 19756 33580 19796 33620
rect 2668 33412 2708 33452
rect 9196 33412 9236 33452
rect 12268 33412 12308 33452
rect 12652 33412 12692 33452
rect 14284 33412 14324 33452
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 2668 33076 2708 33116
rect 3916 33076 3956 33116
rect 5548 33076 5588 33116
rect 18796 33076 18836 33116
rect 19180 33076 19220 33116
rect 19564 33076 19604 33116
rect 19756 32992 19796 33032
rect 8044 32908 8084 32948
rect 2476 32824 2516 32864
rect 3052 32824 3092 32864
rect 1228 32782 1268 32822
rect 3148 32824 3188 32864
rect 3374 32831 3414 32871
rect 3532 32824 3572 32864
rect 3628 32824 3668 32864
rect 3820 32824 3860 32864
rect 3916 32824 3956 32864
rect 4108 32824 4148 32864
rect 5356 32824 5396 32864
rect 5740 32824 5780 32864
rect 6988 32824 7028 32864
rect 7468 32824 7508 32864
rect 7564 32824 7604 32864
rect 9052 32866 9092 32906
rect 10540 32908 10580 32948
rect 10636 32908 10676 32948
rect 17164 32908 17204 32948
rect 7948 32824 7988 32864
rect 8524 32824 8564 32864
rect 10060 32824 10100 32864
rect 10156 32824 10196 32864
rect 11116 32824 11156 32864
rect 11596 32829 11636 32869
rect 13612 32866 13652 32906
rect 17260 32908 17300 32948
rect 18604 32908 18644 32948
rect 18988 32908 19028 32948
rect 19372 32908 19412 32948
rect 20044 32908 20084 32948
rect 11980 32824 12020 32864
rect 13228 32824 13268 32864
rect 14860 32845 14900 32885
rect 16684 32824 16724 32864
rect 16780 32824 16820 32864
rect 17740 32824 17780 32864
rect 18220 32838 18260 32878
rect 7180 32740 7220 32780
rect 11788 32740 11828 32780
rect 18412 32740 18452 32780
rect 2860 32656 2900 32696
rect 9196 32656 9236 32696
rect 13420 32656 13460 32696
rect 15052 32656 15092 32696
rect 20236 32656 20276 32696
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 2668 32320 2708 32360
rect 4300 32320 4340 32360
rect 4972 32320 5012 32360
rect 8044 32320 8084 32360
rect 9868 32320 9908 32360
rect 11596 32320 11636 32360
rect 11980 32320 12020 32360
rect 12748 32320 12788 32360
rect 17164 32320 17204 32360
rect 20236 32320 20276 32360
rect 14956 32236 14996 32276
rect 16972 32236 17012 32276
rect 1228 32152 1268 32192
rect 2476 32152 2516 32192
rect 2860 32152 2900 32192
rect 4108 32152 4148 32192
rect 4492 32152 4532 32192
rect 4588 32152 4628 32192
rect 4780 32152 4820 32192
rect 5068 32152 5108 32192
rect 7756 32152 7796 32192
rect 7852 32152 7892 32192
rect 8428 32152 8468 32192
rect 9676 32152 9716 32192
rect 10156 32152 10196 32192
rect 11404 32152 11444 32192
rect 12460 32152 12500 32192
rect 12556 32152 12596 32192
rect 13228 32152 13268 32192
rect 13324 32152 13364 32192
rect 13708 32152 13748 32192
rect 13804 32152 13844 32192
rect 14284 32152 14324 32192
rect 14812 32142 14852 32182
rect 15244 32152 15284 32192
rect 15340 32152 15380 32192
rect 15724 32152 15764 32192
rect 15820 32152 15860 32192
rect 16300 32152 16340 32192
rect 16780 32138 16820 32178
rect 17356 32152 17396 32192
rect 18604 32152 18644 32192
rect 18796 32152 18836 32192
rect 20044 32152 20084 32192
rect 4492 31984 4532 32024
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 5452 31480 5492 31520
rect 13132 31480 13172 31520
rect 14764 31480 14804 31520
rect 16972 31480 17012 31520
rect 19948 31480 19988 31520
rect 2956 31396 2996 31436
rect 4300 31396 4340 31436
rect 11212 31396 11252 31436
rect 2380 31312 2420 31352
rect 2476 31312 2516 31352
rect 2860 31312 2900 31352
rect 3436 31312 3476 31352
rect 3964 31321 4004 31361
rect 4780 31312 4820 31352
rect 5068 31312 5108 31352
rect 5644 31312 5684 31352
rect 6892 31312 6932 31352
rect 7276 31312 7316 31352
rect 8524 31312 8564 31352
rect 8908 31312 8948 31352
rect 10156 31312 10196 31352
rect 10636 31312 10676 31352
rect 10732 31312 10772 31352
rect 12220 31354 12260 31394
rect 17740 31396 17780 31436
rect 19372 31396 19412 31436
rect 19756 31396 19796 31436
rect 11116 31312 11156 31352
rect 11692 31312 11732 31352
rect 13324 31312 13364 31352
rect 14572 31312 14612 31352
rect 15532 31312 15572 31352
rect 16780 31312 16820 31352
rect 17260 31312 17300 31352
rect 17356 31312 17396 31352
rect 17836 31312 17876 31352
rect 18316 31312 18356 31352
rect 18796 31317 18836 31357
rect 4108 31228 4148 31268
rect 5164 31228 5204 31268
rect 10348 31228 10388 31268
rect 4492 31144 4532 31184
rect 7084 31144 7124 31184
rect 8716 31144 8756 31184
rect 12364 31144 12404 31184
rect 13036 31144 13076 31184
rect 18988 31144 19028 31184
rect 19564 31144 19604 31184
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 1804 30808 1844 30848
rect 14764 30808 14804 30848
rect 16396 30808 16436 30848
rect 17356 30808 17396 30848
rect 19276 30808 19316 30848
rect 19660 30808 19700 30848
rect 6796 30724 6836 30764
rect 9388 30724 9428 30764
rect 12364 30724 12404 30764
rect 3340 30640 3380 30680
rect 4588 30640 4628 30680
rect 5068 30640 5108 30680
rect 5164 30640 5204 30680
rect 6124 30640 6164 30680
rect 6604 30626 6644 30666
rect 6988 30640 7028 30680
rect 7084 30640 7124 30680
rect 7180 30640 7220 30680
rect 7276 30640 7316 30680
rect 7660 30640 7700 30680
rect 7756 30621 7796 30661
rect 8140 30640 8180 30680
rect 8716 30640 8756 30680
rect 9196 30635 9236 30675
rect 10636 30640 10676 30680
rect 10732 30640 10772 30680
rect 11116 30640 11156 30680
rect 11212 30640 11252 30680
rect 11692 30640 11732 30680
rect 13324 30640 13364 30680
rect 14572 30640 14612 30680
rect 14956 30640 14996 30680
rect 16204 30640 16244 30680
rect 17836 30640 17876 30680
rect 19084 30640 19124 30680
rect 5548 30556 5588 30596
rect 5644 30556 5684 30596
rect 8236 30556 8276 30596
rect 12220 30598 12260 30638
rect 16780 30556 16820 30596
rect 17164 30556 17204 30596
rect 19468 30556 19508 30596
rect 19852 30556 19892 30596
rect 4780 30388 4820 30428
rect 16972 30388 17012 30428
rect 20044 30388 20084 30428
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 3436 30052 3476 30092
rect 6220 30052 6260 30092
rect 6412 30052 6452 30092
rect 10540 30052 10580 30092
rect 12460 30052 12500 30092
rect 19852 30052 19892 30092
rect 20236 30052 20276 30092
rect 1804 29968 1844 30008
rect 14860 29884 14900 29924
rect 16780 29884 16820 29924
rect 17164 29884 17204 29924
rect 18220 29884 18260 29924
rect 19660 29884 19700 29924
rect 20044 29884 20084 29924
rect 1996 29800 2036 29840
rect 3244 29800 3284 29840
rect 3724 29800 3764 29840
rect 3820 29800 3860 29840
rect 3916 29800 3956 29840
rect 4108 29800 4148 29840
rect 5356 29800 5396 29840
rect 5836 29800 5876 29840
rect 5932 29800 5972 29840
rect 6028 29800 6068 29840
rect 6508 29800 6548 29840
rect 7276 29800 7316 29840
rect 8524 29800 8564 29840
rect 9100 29800 9140 29840
rect 10348 29800 10388 29840
rect 11020 29800 11060 29840
rect 12268 29800 12308 29840
rect 13708 29800 13748 29840
rect 13804 29800 13844 29840
rect 13996 29800 14036 29840
rect 14284 29800 14324 29840
rect 14380 29800 14420 29840
rect 14764 29800 14804 29840
rect 15340 29800 15380 29840
rect 15820 29805 15860 29845
rect 17644 29800 17684 29840
rect 17740 29800 17780 29840
rect 18124 29800 18164 29840
rect 18700 29800 18740 29840
rect 19228 29809 19268 29849
rect 5548 29716 5588 29756
rect 13900 29716 13940 29756
rect 3628 29632 3668 29672
rect 8716 29632 8756 29672
rect 16012 29632 16052 29672
rect 16972 29632 17012 29672
rect 17356 29632 17396 29672
rect 19372 29632 19412 29672
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 1804 29296 1844 29336
rect 1996 29296 2036 29336
rect 4780 29296 4820 29336
rect 4972 29296 5012 29336
rect 11980 29296 12020 29336
rect 14188 29296 14228 29336
rect 15628 29296 15668 29336
rect 19852 29296 19892 29336
rect 6892 29212 6932 29252
rect 8908 29212 8948 29252
rect 14860 29212 14900 29252
rect 18220 29212 18260 29252
rect 2188 29128 2228 29168
rect 2320 29118 2360 29158
rect 2476 29128 2516 29168
rect 3724 29128 3764 29168
rect 4492 29128 4532 29168
rect 4588 29128 4628 29168
rect 5164 29128 5204 29168
rect 5260 29128 5300 29168
rect 5452 29128 5492 29168
rect 6700 29128 6740 29168
rect 7180 29128 7220 29168
rect 7276 29128 7316 29168
rect 7660 29128 7700 29168
rect 7756 29128 7796 29168
rect 8236 29128 8276 29168
rect 8716 29123 8756 29163
rect 10252 29128 10292 29168
rect 10348 29128 10388 29168
rect 10732 29128 10772 29168
rect 10828 29128 10868 29168
rect 11308 29128 11348 29168
rect 11788 29114 11828 29154
rect 12748 29128 12788 29168
rect 13996 29128 14036 29168
rect 14476 29128 14516 29168
rect 14764 29128 14804 29168
rect 16492 29128 16532 29168
rect 16588 29128 16628 29168
rect 17548 29128 17588 29168
rect 18028 29114 18068 29154
rect 18412 29128 18452 29168
rect 16972 29044 17012 29084
rect 19660 29086 19700 29126
rect 17068 29044 17108 29084
rect 20044 29044 20084 29084
rect 3916 28960 3956 29000
rect 15724 28960 15764 29000
rect 20236 28876 20276 28916
rect 15148 28834 15188 28874
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 11692 28540 11732 28580
rect 12172 28540 12212 28580
rect 15436 28540 15476 28580
rect 15916 28540 15956 28580
rect 18988 28540 19028 28580
rect 19756 28540 19796 28580
rect 20140 28540 20180 28580
rect 1804 28456 1844 28496
rect 15628 28456 15668 28496
rect 3532 28372 3572 28412
rect 19180 28372 19220 28412
rect 19564 28372 19604 28412
rect 19948 28372 19988 28412
rect 3052 28288 3092 28328
rect 3148 28288 3188 28328
rect 3628 28288 3668 28328
rect 4108 28288 4148 28328
rect 4588 28293 4628 28333
rect 5068 28288 5108 28328
rect 6316 28288 6356 28328
rect 6796 28288 6836 28328
rect 6892 28288 6932 28328
rect 7276 28288 7316 28328
rect 7372 28288 7412 28328
rect 7852 28288 7892 28328
rect 8332 28293 8372 28333
rect 10252 28288 10292 28328
rect 11500 28288 11540 28328
rect 11884 28288 11924 28328
rect 12172 28288 12212 28328
rect 12556 28288 12596 28328
rect 13804 28288 13844 28328
rect 13996 28288 14036 28328
rect 15244 28288 15284 28328
rect 16108 28288 16148 28328
rect 17356 28288 17396 28328
rect 17548 28288 17588 28328
rect 18796 28288 18836 28328
rect 4780 28204 4820 28244
rect 6508 28204 6548 28244
rect 1708 28120 1748 28160
rect 8524 28120 8564 28160
rect 12364 28120 12404 28160
rect 19372 28120 19412 28160
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 3148 27784 3188 27824
rect 8236 27784 8276 27824
rect 15436 27784 15476 27824
rect 16588 27784 16628 27824
rect 20044 27784 20084 27824
rect 6508 27700 6548 27740
rect 9868 27700 9908 27740
rect 11884 27700 11924 27740
rect 16012 27700 16052 27740
rect 17452 27700 17492 27740
rect 1708 27616 1748 27656
rect 2956 27616 2996 27656
rect 3340 27616 3380 27656
rect 3532 27616 3572 27656
rect 3724 27616 3764 27656
rect 4972 27616 5012 27656
rect 5452 27616 5492 27656
rect 5740 27616 5780 27656
rect 5836 27616 5876 27656
rect 6316 27616 6356 27656
rect 6412 27616 6452 27656
rect 6604 27616 6644 27656
rect 6796 27616 6836 27656
rect 8044 27616 8084 27656
rect 8428 27616 8468 27656
rect 9676 27616 9716 27656
rect 10156 27616 10196 27656
rect 10252 27616 10292 27656
rect 10732 27616 10772 27656
rect 11212 27616 11252 27656
rect 11692 27602 11732 27642
rect 12076 27616 12116 27656
rect 13324 27616 13364 27656
rect 13996 27616 14036 27656
rect 15244 27616 15284 27656
rect 15916 27616 15956 27656
rect 16108 27616 16148 27656
rect 16492 27605 16532 27645
rect 16684 27616 16724 27656
rect 16780 27616 16820 27656
rect 17644 27602 17684 27642
rect 18124 27616 18164 27656
rect 18604 27616 18644 27656
rect 18700 27616 18740 27656
rect 19084 27616 19124 27656
rect 19180 27616 19220 27656
rect 10636 27532 10676 27572
rect 17068 27532 17108 27572
rect 19468 27532 19508 27572
rect 19852 27532 19892 27572
rect 5164 27448 5204 27488
rect 15724 27448 15764 27488
rect 19660 27448 19700 27488
rect 3532 27364 3572 27404
rect 6124 27364 6164 27404
rect 13516 27364 13556 27404
rect 17260 27364 17300 27404
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 3436 27028 3476 27068
rect 5068 27028 5108 27068
rect 5644 27028 5684 27068
rect 11500 27028 11540 27068
rect 15436 27028 15476 27068
rect 1708 26944 1748 26984
rect 16972 26944 17012 26984
rect 8236 26860 8276 26900
rect 15244 26860 15284 26900
rect 19372 26860 19412 26900
rect 19756 26860 19796 26900
rect 1228 26776 1268 26816
rect 1324 26776 1364 26816
rect 1420 26776 1460 26816
rect 1516 26776 1556 26816
rect 1996 26776 2036 26816
rect 3244 26776 3284 26816
rect 3628 26776 3668 26816
rect 4876 26776 4916 26816
rect 5356 26776 5396 26816
rect 5644 26776 5684 26816
rect 6028 26776 6068 26816
rect 7276 26776 7316 26816
rect 7756 26776 7796 26816
rect 7852 26776 7892 26816
rect 8332 26776 8372 26816
rect 8812 26776 8852 26816
rect 9292 26781 9332 26821
rect 10060 26776 10100 26816
rect 11308 26776 11348 26816
rect 12844 26776 12884 26816
rect 12940 26776 12980 26816
rect 13324 26776 13364 26816
rect 13420 26776 13460 26816
rect 13900 26776 13940 26816
rect 14380 26790 14420 26830
rect 14764 26776 14804 26816
rect 14860 26776 14900 26816
rect 16300 26776 16340 26816
rect 16588 26776 16628 26816
rect 16684 26776 16724 26816
rect 17260 26776 17300 26816
rect 17356 26776 17396 26816
rect 17740 26776 17780 26816
rect 17836 26776 17876 26816
rect 18316 26776 18356 26816
rect 18796 26781 18836 26821
rect 7468 26692 7508 26732
rect 14572 26692 14612 26732
rect 1708 26608 1748 26648
rect 5068 26608 5108 26648
rect 9484 26608 9524 26648
rect 15052 26608 15092 26648
rect 15628 26608 15668 26648
rect 15916 26608 15956 26648
rect 18988 26608 19028 26648
rect 19564 26608 19604 26648
rect 19948 26608 19988 26648
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 1708 26272 1748 26312
rect 3436 26272 3476 26312
rect 3628 26272 3668 26312
rect 8524 26272 8564 26312
rect 10156 26272 10196 26312
rect 17068 26272 17108 26312
rect 18700 26272 18740 26312
rect 19180 26272 19220 26312
rect 1228 26188 1268 26228
rect 1324 26104 1364 26144
rect 1420 26104 1460 26144
rect 1516 26104 1556 26144
rect 1996 26104 2036 26144
rect 3244 26104 3284 26144
rect 3820 26104 3860 26144
rect 5068 26104 5108 26144
rect 5452 26104 5492 26144
rect 6700 26104 6740 26144
rect 7084 26104 7124 26144
rect 8332 26104 8372 26144
rect 8716 26104 8756 26144
rect 9964 26104 10004 26144
rect 12748 26104 12788 26144
rect 12844 26104 12884 26144
rect 13132 26104 13172 26144
rect 13420 26104 13460 26144
rect 13612 26104 13652 26144
rect 13804 26104 13844 26144
rect 15052 26104 15092 26144
rect 15628 26104 15668 26144
rect 16876 26104 16916 26144
rect 17260 26104 17300 26144
rect 18508 26104 18548 26144
rect 18892 26104 18932 26144
rect 18988 26104 19028 26144
rect 19756 26104 19796 26144
rect 19852 26104 19892 26144
rect 19948 26104 19988 26144
rect 20044 26104 20084 26144
rect 19372 26020 19412 26060
rect 6892 25852 6932 25892
rect 12460 25852 12500 25892
rect 13612 25852 13652 25892
rect 15244 25852 15284 25892
rect 19564 25852 19604 25892
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 1996 25516 2036 25556
rect 11596 25516 11636 25556
rect 17452 25516 17492 25556
rect 19084 25516 19124 25556
rect 1708 25432 1748 25472
rect 13036 25348 13076 25388
rect 1228 25264 1268 25304
rect 1420 25264 1460 25304
rect 1516 25264 1556 25304
rect 2188 25264 2228 25304
rect 3436 25264 3476 25304
rect 4012 25278 4052 25318
rect 4492 25264 4532 25304
rect 4972 25264 5012 25304
rect 5068 25264 5108 25304
rect 5452 25264 5492 25304
rect 5548 25264 5588 25304
rect 5836 25264 5876 25304
rect 5932 25264 5972 25304
rect 6988 25264 7028 25304
rect 7084 25264 7124 25304
rect 7468 25264 7508 25304
rect 7564 25264 7604 25304
rect 8044 25264 8084 25304
rect 8524 25269 8564 25309
rect 10156 25264 10196 25304
rect 11404 25264 11444 25304
rect 11980 25269 12020 25309
rect 12460 25264 12500 25304
rect 12940 25264 12980 25304
rect 13420 25264 13460 25304
rect 13516 25264 13556 25304
rect 13996 25264 14036 25304
rect 15244 25264 15284 25304
rect 16012 25264 16052 25304
rect 17260 25264 17300 25304
rect 17644 25264 17684 25304
rect 18892 25264 18932 25304
rect 19276 25243 19316 25283
rect 19372 25264 19412 25304
rect 19468 25243 19508 25283
rect 19564 25264 19604 25304
rect 19756 25264 19796 25304
rect 19852 25264 19892 25304
rect 3820 25180 3860 25220
rect 8716 25138 8756 25178
rect 11788 25180 11828 25220
rect 15436 25180 15476 25220
rect 1324 25096 1364 25136
rect 6124 25096 6164 25136
rect 15628 25096 15668 25136
rect 20044 25096 20084 25136
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 1420 24760 1460 24800
rect 1708 24760 1748 24800
rect 3436 24760 3476 24800
rect 7564 24760 7604 24800
rect 11404 24760 11444 24800
rect 13036 24760 13076 24800
rect 13324 24760 13364 24800
rect 13804 24760 13844 24800
rect 15436 24760 15476 24800
rect 3724 24676 3764 24716
rect 9580 24676 9620 24716
rect 17740 24676 17780 24716
rect 20236 24676 20276 24716
rect 1324 24592 1364 24632
rect 1516 24592 1556 24632
rect 1996 24592 2036 24632
rect 3244 24592 3284 24632
rect 3916 24587 3956 24627
rect 4396 24592 4436 24632
rect 5356 24592 5396 24632
rect 5452 24592 5492 24632
rect 6124 24592 6164 24632
rect 7372 24592 7412 24632
rect 7852 24592 7892 24632
rect 7948 24592 7988 24632
rect 8332 24592 8372 24632
rect 8908 24592 8948 24632
rect 9388 24578 9428 24618
rect 9964 24592 10004 24632
rect 11212 24592 11252 24632
rect 11596 24592 11636 24632
rect 12844 24592 12884 24632
rect 13228 24592 13268 24632
rect 13420 24592 13460 24632
rect 13516 24592 13556 24632
rect 13900 24613 13940 24653
rect 13996 24592 14036 24632
rect 14092 24592 14132 24632
rect 14284 24592 14324 24632
rect 14476 24592 14516 24632
rect 14572 24592 14612 24632
rect 14860 24592 14900 24632
rect 16012 24592 16052 24632
rect 16108 24592 16148 24632
rect 16492 24592 16532 24632
rect 17068 24592 17108 24632
rect 17548 24587 17588 24627
rect 17932 24592 17972 24632
rect 18124 24592 18164 24632
rect 18220 24592 18260 24632
rect 18508 24573 18548 24613
rect 18604 24592 18644 24632
rect 18988 24592 19028 24632
rect 19564 24592 19604 24632
rect 20044 24578 20084 24618
rect 4876 24508 4916 24548
rect 4972 24508 5012 24548
rect 8428 24508 8468 24548
rect 14764 24508 14804 24548
rect 15244 24508 15284 24548
rect 16588 24508 16628 24548
rect 19084 24508 19124 24548
rect 15628 24424 15668 24464
rect 17932 24340 17972 24380
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 3628 24004 3668 24044
rect 9388 24004 9428 24044
rect 1516 23920 1556 23960
rect 3436 23920 3476 23960
rect 4588 23920 4628 23960
rect 7468 23920 7508 23960
rect 17356 23920 17396 23960
rect 18124 23920 18164 23960
rect 1804 23836 1844 23876
rect 1996 23752 2036 23792
rect 3244 23752 3284 23792
rect 4012 23752 4052 23792
rect 4300 23752 4340 23792
rect 4588 23752 4628 23792
rect 4780 23752 4820 23792
rect 4876 23752 4916 23792
rect 5068 23752 5108 23792
rect 5164 23752 5204 23792
rect 6028 23752 6068 23792
rect 7276 23752 7316 23792
rect 7948 23752 7988 23792
rect 9196 23752 9236 23792
rect 9772 23752 9812 23792
rect 11020 23752 11060 23792
rect 11212 23752 11252 23792
rect 11308 23752 11348 23792
rect 11500 23752 11540 23792
rect 15916 23794 15956 23834
rect 11596 23752 11636 23792
rect 11697 23752 11737 23792
rect 13228 23752 13268 23792
rect 14476 23752 14516 23792
rect 17164 23752 17204 23792
rect 17548 23752 17588 23792
rect 17740 23752 17780 23792
rect 18316 23752 18356 23792
rect 19564 23752 19604 23792
rect 19948 23752 19988 23792
rect 20044 23752 20084 23792
rect 3916 23668 3956 23708
rect 5356 23584 5396 23624
rect 9580 23584 9620 23624
rect 11692 23584 11732 23624
rect 14668 23584 14708 23624
rect 15628 23584 15668 23624
rect 17644 23584 17684 23624
rect 19756 23584 19796 23624
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 4012 23248 4052 23288
rect 9292 23248 9332 23288
rect 9676 23248 9716 23288
rect 14860 23248 14900 23288
rect 18892 23248 18932 23288
rect 20140 23248 20180 23288
rect 3148 23164 3188 23204
rect 3628 23164 3668 23204
rect 5932 23164 5972 23204
rect 7564 23164 7604 23204
rect 12844 23164 12884 23204
rect 1708 23080 1748 23120
rect 2956 23080 2996 23120
rect 3340 23080 3380 23120
rect 3436 23080 3476 23120
rect 3532 23080 3572 23120
rect 3820 23080 3860 23120
rect 4108 23080 4148 23120
rect 4492 23080 4532 23120
rect 5740 23080 5780 23120
rect 6508 23080 6548 23120
rect 6796 23080 6836 23120
rect 6892 23080 6932 23120
rect 7468 23080 7508 23120
rect 7660 23080 7700 23120
rect 7756 23080 7796 23120
rect 7948 23080 7988 23120
rect 8140 23080 8180 23120
rect 8236 23080 8276 23120
rect 8716 23080 8756 23120
rect 8908 23080 8948 23120
rect 9004 23080 9044 23120
rect 9196 23080 9236 23120
rect 9388 23080 9428 23120
rect 9484 23080 9524 23120
rect 9868 23080 9908 23120
rect 11116 23080 11156 23120
rect 11404 23080 11444 23120
rect 12652 23080 12692 23120
rect 13132 23080 13172 23120
rect 13228 23080 13268 23120
rect 13612 23080 13652 23120
rect 14188 23080 14228 23120
rect 14668 23075 14708 23115
rect 15916 23080 15956 23120
rect 16012 23080 16052 23120
rect 16204 23080 16244 23120
rect 16588 23080 16628 23120
rect 16876 23080 16916 23120
rect 16972 23080 17012 23120
rect 17452 23080 17492 23120
rect 18700 23080 18740 23120
rect 19121 23080 19161 23120
rect 19276 23080 19316 23120
rect 19372 23080 19412 23120
rect 19564 23080 19604 23120
rect 19660 23080 19700 23120
rect 19852 23080 19892 23120
rect 19948 23080 19988 23120
rect 13708 22996 13748 23036
rect 15244 22996 15284 23036
rect 7948 22912 7988 22952
rect 9004 22912 9044 22952
rect 15628 22912 15668 22952
rect 17260 22912 17300 22952
rect 7180 22828 7220 22868
rect 15436 22828 15476 22868
rect 16204 22828 16244 22868
rect 19660 22828 19700 22868
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 2668 22492 2708 22532
rect 9580 22492 9620 22532
rect 18124 22492 18164 22532
rect 20044 22492 20084 22532
rect 5452 22408 5492 22448
rect 12364 22408 12404 22448
rect 13228 22324 13268 22364
rect 1228 22240 1268 22280
rect 2476 22240 2516 22280
rect 3052 22259 3092 22299
rect 3148 22240 3188 22280
rect 3532 22240 3572 22280
rect 3628 22240 3668 22280
rect 4108 22240 4148 22280
rect 4588 22254 4628 22294
rect 5260 22240 5300 22280
rect 5452 22240 5492 22280
rect 5836 22245 5876 22285
rect 6316 22240 6356 22280
rect 6796 22240 6836 22280
rect 6892 22240 6932 22280
rect 7276 22240 7316 22280
rect 7372 22259 7412 22299
rect 7852 22240 7892 22280
rect 7948 22240 7988 22280
rect 8140 22240 8180 22280
rect 9388 22240 9428 22280
rect 9772 22240 9812 22280
rect 9868 22240 9908 22280
rect 10060 22240 10100 22280
rect 10156 22240 10196 22280
rect 10257 22240 10297 22280
rect 10924 22240 10964 22280
rect 12172 22240 12212 22280
rect 12652 22240 12692 22280
rect 12748 22259 12788 22299
rect 13132 22240 13172 22280
rect 13708 22240 13748 22280
rect 14188 22245 14228 22285
rect 14572 22240 14612 22280
rect 14764 22240 14804 22280
rect 14860 22240 14900 22280
rect 15052 22240 15092 22280
rect 15148 22240 15188 22280
rect 16007 22240 16047 22280
rect 16108 22240 16148 22280
rect 16204 22240 16244 22280
rect 16396 22240 16436 22280
rect 16492 22240 16532 22280
rect 16684 22240 16724 22280
rect 17932 22240 17972 22280
rect 18604 22240 18644 22280
rect 19852 22240 19892 22280
rect 4780 22156 4820 22196
rect 5644 22156 5684 22196
rect 7660 22072 7700 22112
rect 10156 22072 10196 22112
rect 14380 22072 14420 22112
rect 14668 22072 14708 22112
rect 15340 22072 15380 22112
rect 15628 22072 15668 22112
rect 16108 22072 16148 22112
rect 18412 22072 18452 22112
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 2956 21736 2996 21776
rect 3436 21736 3476 21776
rect 3916 21736 3956 21776
rect 4684 21736 4724 21776
rect 6892 21736 6932 21776
rect 9484 21736 9524 21776
rect 9964 21736 10004 21776
rect 11308 21736 11348 21776
rect 14668 21736 14708 21776
rect 19084 21736 19124 21776
rect 19276 21736 19316 21776
rect 7564 21652 7604 21692
rect 13996 21652 14036 21692
rect 1516 21568 1556 21608
rect 2764 21568 2804 21608
rect 3628 21568 3668 21608
rect 3724 21568 3764 21608
rect 4012 21568 4052 21608
rect 4108 21568 4148 21608
rect 4204 21568 4244 21608
rect 4396 21568 4436 21608
rect 4492 21568 4532 21608
rect 5452 21568 5492 21608
rect 6700 21568 6740 21608
rect 7180 21568 7220 21608
rect 7468 21568 7508 21608
rect 8044 21568 8084 21608
rect 9292 21568 9332 21608
rect 9676 21568 9716 21608
rect 9772 21568 9812 21608
rect 11020 21568 11060 21608
rect 11116 21568 11156 21608
rect 12556 21568 12596 21608
rect 13804 21568 13844 21608
rect 14476 21568 14516 21608
rect 14572 21568 14612 21608
rect 14764 21568 14804 21608
rect 14860 21568 14900 21608
rect 15015 21568 15055 21608
rect 15244 21568 15284 21608
rect 15340 21568 15380 21608
rect 15532 21568 15572 21608
rect 16780 21568 16820 21608
rect 17164 21568 17204 21608
rect 17260 21568 17300 21608
rect 17452 21568 17492 21608
rect 17644 21568 17684 21608
rect 18892 21568 18932 21608
rect 19468 21568 19508 21608
rect 19564 21568 19604 21608
rect 19852 21568 19892 21608
rect 19948 21568 19988 21608
rect 20140 21568 20180 21608
rect 7852 21400 7892 21440
rect 17164 21400 17204 21440
rect 19852 21400 19892 21440
rect 16972 21316 17012 21356
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 2668 20980 2708 21020
rect 6892 20980 6932 21020
rect 14860 20980 14900 21020
rect 17068 20980 17108 21020
rect 17452 20980 17492 21020
rect 20236 20980 20276 21020
rect 11020 20896 11060 20936
rect 12940 20896 12980 20936
rect 13132 20896 13172 20936
rect 17644 20896 17684 20936
rect 3436 20812 3476 20852
rect 3532 20812 3572 20852
rect 17260 20812 17300 20852
rect 1228 20728 1268 20768
rect 2476 20728 2516 20768
rect 2956 20728 2996 20768
rect 3052 20728 3092 20768
rect 4012 20728 4052 20768
rect 4492 20733 4532 20773
rect 5452 20728 5492 20768
rect 6700 20728 6740 20768
rect 7084 20728 7124 20768
rect 8332 20728 8372 20768
rect 9580 20728 9620 20768
rect 10828 20728 10868 20768
rect 11212 20728 11252 20768
rect 11308 20728 11348 20768
rect 11500 20728 11540 20768
rect 11596 20728 11636 20768
rect 11753 20743 11793 20783
rect 11980 20728 12020 20768
rect 12076 20728 12116 20768
rect 12652 20728 12692 20768
rect 12844 20728 12884 20768
rect 12940 20728 12980 20768
rect 13420 20728 13460 20768
rect 14668 20728 14708 20768
rect 15340 20728 15380 20768
rect 15436 20728 15476 20768
rect 15628 20728 15668 20768
rect 16876 20728 16916 20768
rect 18023 20728 18063 20768
rect 18124 20728 18164 20768
rect 18220 20728 18260 20768
rect 18412 20728 18452 20768
rect 18508 20728 18548 20768
rect 18796 20728 18836 20768
rect 20044 20728 20084 20768
rect 4684 20644 4724 20684
rect 6892 20560 6932 20600
rect 8524 20560 8564 20600
rect 11404 20560 11444 20600
rect 12268 20560 12308 20600
rect 15148 20560 15188 20600
rect 17740 20560 17780 20600
rect 18028 20560 18068 20600
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 8812 20224 8852 20264
rect 9388 20224 9428 20264
rect 11500 20224 11540 20264
rect 13228 20224 13268 20264
rect 14956 20224 14996 20264
rect 18892 20224 18932 20264
rect 2668 20140 2708 20180
rect 6316 20140 6356 20180
rect 7276 20140 7316 20180
rect 11116 20140 11156 20180
rect 1228 20056 1268 20096
rect 2476 20056 2516 20096
rect 2860 20056 2900 20096
rect 4108 20056 4148 20096
rect 4588 20056 4628 20096
rect 4684 20056 4724 20096
rect 5164 20056 5204 20096
rect 5644 20056 5684 20096
rect 6124 20051 6164 20091
rect 7180 20056 7220 20096
rect 7852 20056 7892 20096
rect 8044 20056 8084 20096
rect 8140 20056 8180 20096
rect 8332 20056 8372 20096
rect 8428 20056 8468 20096
rect 8572 20041 8612 20081
rect 8716 20056 8756 20096
rect 8873 20041 8913 20081
rect 9100 20056 9140 20096
rect 9196 20056 9236 20096
rect 9676 20056 9716 20096
rect 10924 20056 10964 20096
rect 11308 20056 11348 20096
rect 11404 20056 11444 20096
rect 11596 20056 11636 20096
rect 11788 20056 11828 20096
rect 13036 20056 13076 20096
rect 13516 20056 13556 20096
rect 14764 20056 14804 20096
rect 15820 20056 15860 20096
rect 17068 20056 17108 20096
rect 17452 20056 17492 20096
rect 18700 20056 18740 20096
rect 19175 20056 19215 20096
rect 19276 20056 19316 20096
rect 19372 20056 19412 20096
rect 19564 20056 19604 20096
rect 19660 20056 19700 20096
rect 19852 20056 19892 20096
rect 19948 20056 19988 20096
rect 20044 20056 20084 20096
rect 20140 20051 20180 20091
rect 5068 19972 5108 20012
rect 4300 19888 4340 19928
rect 8140 19888 8180 19928
rect 17260 19888 17300 19928
rect 19660 19804 19700 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 2668 19468 2708 19508
rect 4492 19468 4532 19508
rect 6220 19468 6260 19508
rect 8236 19468 8276 19508
rect 10252 19468 10292 19508
rect 13132 19468 13172 19508
rect 17260 19468 17300 19508
rect 17548 19384 17588 19424
rect 19756 19384 19796 19424
rect 10060 19258 10100 19298
rect 1228 19216 1268 19256
rect 2476 19216 2516 19256
rect 3052 19216 3092 19256
rect 4300 19216 4340 19256
rect 4780 19216 4820 19256
rect 6028 19216 6068 19256
rect 6796 19216 6836 19256
rect 8044 19216 8084 19256
rect 8812 19216 8852 19256
rect 10540 19216 10580 19256
rect 10636 19216 10676 19256
rect 10828 19216 10868 19256
rect 10924 19216 10964 19256
rect 11081 19231 11121 19271
rect 11692 19216 11732 19256
rect 12940 19216 12980 19256
rect 13324 19216 13364 19256
rect 13420 19216 13460 19256
rect 13612 19216 13652 19256
rect 13708 19216 13748 19256
rect 13809 19216 13849 19256
rect 14092 19216 14132 19256
rect 14188 19216 14228 19256
rect 15820 19216 15860 19256
rect 17068 19216 17108 19256
rect 17836 19216 17876 19256
rect 19084 19216 19124 19256
rect 19660 19216 19700 19256
rect 19756 19216 19796 19256
rect 19948 19216 19988 19256
rect 19276 19132 19316 19172
rect 10732 19048 10772 19088
rect 13132 19048 13172 19088
rect 13708 19048 13748 19088
rect 14380 19048 14420 19088
rect 17260 19048 17300 19088
rect 17644 19048 17684 19088
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 2668 18712 2708 18752
rect 6124 18712 6164 18752
rect 8236 18712 8276 18752
rect 10828 18712 10868 18752
rect 19372 18754 19412 18794
rect 14668 18712 14708 18752
rect 16972 18712 17012 18752
rect 20236 18712 20276 18752
rect 5068 18628 5108 18668
rect 10156 18628 10196 18668
rect 16684 18628 16724 18668
rect 18892 18628 18932 18668
rect 1228 18544 1268 18584
rect 2476 18544 2516 18584
rect 3340 18544 3380 18584
rect 4588 18544 4628 18584
rect 4972 18544 5012 18584
rect 5164 18544 5204 18584
rect 5356 18544 5396 18584
rect 5644 18544 5684 18584
rect 5836 18544 5876 18584
rect 5932 18544 5972 18584
rect 6316 18544 6356 18584
rect 6501 18543 6541 18583
rect 6796 18544 6836 18584
rect 8044 18544 8084 18584
rect 8716 18544 8756 18584
rect 9964 18544 10004 18584
rect 10540 18544 10580 18584
rect 10636 18544 10676 18584
rect 11404 18544 11444 18584
rect 12652 18544 12692 18584
rect 13228 18544 13268 18584
rect 14476 18544 14516 18584
rect 14956 18544 14996 18584
rect 15052 18544 15092 18584
rect 15532 18544 15572 18584
rect 16012 18544 16052 18584
rect 16492 18530 16532 18570
rect 17164 18544 17204 18584
rect 17260 18544 17300 18584
rect 18700 18544 18740 18584
rect 19084 18544 19124 18584
rect 17452 18502 17492 18542
rect 19180 18544 19220 18584
rect 19564 18544 19604 18584
rect 19660 18544 19700 18584
rect 19852 18544 19892 18584
rect 15436 18460 15476 18500
rect 20044 18460 20084 18500
rect 3052 18376 3092 18416
rect 5644 18376 5684 18416
rect 19564 18376 19604 18416
rect 4780 18292 4820 18332
rect 6412 18292 6452 18332
rect 12844 18292 12884 18332
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 2092 17956 2132 17996
rect 16780 17956 16820 17996
rect 17164 17956 17204 17996
rect 18796 17956 18836 17996
rect 10444 17872 10484 17912
rect 12844 17872 12884 17912
rect 13804 17872 13844 17912
rect 2860 17788 2900 17828
rect 2956 17788 2996 17828
rect 16204 17788 16244 17828
rect 16588 17788 16628 17828
rect 16972 17788 17012 17828
rect 1804 17704 1844 17744
rect 1900 17717 1940 17757
rect 2092 17704 2132 17744
rect 2380 17704 2420 17744
rect 2476 17704 2516 17744
rect 3436 17704 3476 17744
rect 3916 17709 3956 17749
rect 4396 17704 4436 17744
rect 4588 17704 4628 17744
rect 4684 17704 4724 17744
rect 5068 17704 5108 17744
rect 5164 17704 5204 17744
rect 5356 17704 5396 17744
rect 6604 17704 6644 17744
rect 7084 17704 7124 17744
rect 7180 17704 7220 17744
rect 7564 17704 7604 17744
rect 7660 17704 7700 17744
rect 8140 17704 8180 17744
rect 8620 17718 8660 17758
rect 9196 17709 9236 17749
rect 9388 17704 9428 17744
rect 9484 17704 9524 17744
rect 9676 17704 9716 17744
rect 9772 17704 9812 17744
rect 10156 17704 10196 17744
rect 10348 17704 10388 17744
rect 10444 17704 10484 17744
rect 10636 17704 10676 17744
rect 10732 17704 10772 17744
rect 10924 17704 10964 17744
rect 12652 17746 12692 17786
rect 11020 17704 11060 17744
rect 11121 17704 11161 17744
rect 11404 17704 11444 17744
rect 13084 17715 13124 17755
rect 13228 17704 13268 17744
rect 13324 17719 13364 17759
rect 13516 17704 13556 17744
rect 13612 17704 13652 17744
rect 13804 17704 13844 17744
rect 13900 17704 13940 17744
rect 14092 17704 14132 17744
rect 14284 17704 14324 17744
rect 15532 17704 15572 17744
rect 17356 17704 17396 17744
rect 18604 17704 18644 17744
rect 19079 17704 19119 17744
rect 19180 17704 19220 17744
rect 19276 17704 19316 17744
rect 19468 17704 19508 17744
rect 19564 17704 19604 17744
rect 19756 17704 19796 17744
rect 19852 17704 19892 17744
rect 4108 17620 4148 17660
rect 6796 17620 6836 17660
rect 9292 17620 9332 17660
rect 4492 17536 4532 17576
rect 4876 17536 4916 17576
rect 9964 17536 10004 17576
rect 11116 17536 11156 17576
rect 13132 17536 13172 17576
rect 15724 17536 15764 17576
rect 8812 17494 8852 17534
rect 16396 17536 16436 17576
rect 19084 17536 19124 17576
rect 20044 17536 20084 17576
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 3532 17200 3572 17240
rect 3916 17200 3956 17240
rect 9484 17200 9524 17240
rect 16588 17200 16628 17240
rect 17164 17200 17204 17240
rect 19084 17200 19124 17240
rect 19852 17200 19892 17240
rect 20236 17200 20276 17240
rect 7276 17116 7316 17156
rect 9292 17116 9332 17156
rect 12748 17116 12788 17156
rect 14764 17116 14804 17156
rect 1228 17032 1268 17072
rect 2476 17032 2516 17072
rect 2956 17032 2996 17072
rect 3239 17032 3279 17072
rect 3340 17032 3380 17072
rect 3436 17032 3476 17072
rect 3628 17032 3668 17072
rect 3724 17032 3764 17072
rect 4108 17032 4148 17072
rect 5356 17032 5396 17072
rect 5836 17032 5876 17072
rect 7084 17032 7124 17072
rect 7564 17032 7604 17072
rect 7660 17032 7700 17072
rect 8620 17032 8660 17072
rect 9100 17018 9140 17058
rect 9676 17032 9716 17072
rect 10924 17032 10964 17072
rect 11308 17032 11348 17072
rect 12556 17032 12596 17072
rect 13036 17032 13076 17072
rect 13132 17052 13172 17092
rect 14092 17032 14132 17072
rect 15148 17032 15188 17072
rect 16396 17032 16436 17072
rect 17644 17032 17684 17072
rect 18892 17032 18932 17072
rect 8044 16948 8084 16988
rect 8140 16948 8180 16988
rect 13516 16948 13556 16988
rect 13612 16948 13652 16988
rect 14620 16990 14660 17030
rect 16972 16948 17012 16988
rect 19276 16948 19316 16988
rect 19660 16948 19700 16988
rect 20044 16948 20084 16988
rect 2668 16864 2708 16904
rect 2860 16864 2900 16904
rect 19468 16780 19508 16820
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 5260 16444 5300 16484
rect 9100 16444 9140 16484
rect 9388 16444 9428 16484
rect 14860 16444 14900 16484
rect 15436 16360 15476 16400
rect 17452 16360 17492 16400
rect 17836 16360 17876 16400
rect 15244 16276 15284 16316
rect 17260 16276 17300 16316
rect 17644 16276 17684 16316
rect 2284 16192 2324 16232
rect 3532 16192 3572 16232
rect 4108 16192 4148 16232
rect 4204 16192 4244 16232
rect 4588 16192 4628 16232
rect 4876 16192 4916 16232
rect 5548 16192 5588 16232
rect 6796 16192 6836 16232
rect 7660 16192 7700 16232
rect 8908 16192 8948 16232
rect 9580 16192 9620 16232
rect 10828 16192 10868 16232
rect 12844 16192 12884 16232
rect 12940 16192 12980 16232
rect 13420 16192 13460 16232
rect 14668 16192 14708 16232
rect 15628 16192 15668 16232
rect 16876 16192 16916 16232
rect 18028 16192 18068 16232
rect 18220 16192 18260 16232
rect 18515 16197 18555 16237
rect 18700 16192 18740 16232
rect 18796 16192 18836 16232
rect 18988 16192 19028 16232
rect 19084 16192 19124 16232
rect 19276 16192 19316 16232
rect 19372 16192 19412 16232
rect 19527 16192 19567 16232
rect 19756 16192 19796 16232
rect 19852 16192 19892 16232
rect 3724 16108 3764 16148
rect 4972 16108 5012 16148
rect 3916 16024 3956 16064
rect 6988 16024 7028 16064
rect 13132 16024 13172 16064
rect 17068 16024 17108 16064
rect 18124 16024 18164 16064
rect 18604 16024 18644 16064
rect 19180 16024 19220 16064
rect 20044 16024 20084 16064
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 3052 15688 3092 15728
rect 3628 15688 3668 15728
rect 16972 15688 17012 15728
rect 19084 15688 19124 15728
rect 19468 15688 19508 15728
rect 19852 15688 19892 15728
rect 20236 15688 20276 15728
rect 5644 15604 5684 15644
rect 8620 15604 8660 15644
rect 1612 15520 1652 15560
rect 2860 15520 2900 15560
rect 3916 15520 3956 15560
rect 4012 15520 4052 15560
rect 4492 15520 4532 15560
rect 4972 15520 5012 15560
rect 5452 15506 5492 15546
rect 6892 15520 6932 15560
rect 6988 15520 7028 15560
rect 7948 15520 7988 15560
rect 8428 15506 8468 15546
rect 8908 15520 8948 15560
rect 10156 15520 10196 15560
rect 10540 15520 10580 15560
rect 10732 15520 10772 15560
rect 11596 15520 11636 15560
rect 12844 15520 12884 15560
rect 13708 15520 13748 15560
rect 14956 15520 14996 15560
rect 15532 15520 15572 15560
rect 16780 15520 16820 15560
rect 17164 15520 17204 15560
rect 17260 15520 17300 15560
rect 17452 15520 17492 15560
rect 17644 15520 17684 15560
rect 18892 15520 18932 15560
rect 3436 15436 3476 15476
rect 4396 15436 4436 15476
rect 7372 15436 7412 15476
rect 7468 15436 7508 15476
rect 19276 15436 19316 15476
rect 19660 15436 19700 15476
rect 20044 15436 20084 15476
rect 13420 15352 13460 15392
rect 10348 15268 10388 15308
rect 10636 15268 10676 15308
rect 13036 15268 13076 15308
rect 15148 15268 15188 15308
rect 17452 15268 17492 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 2668 14932 2708 14972
rect 5452 14932 5492 14972
rect 8140 14932 8180 14972
rect 17260 14932 17300 14972
rect 19180 14932 19220 14972
rect 20044 14932 20084 14972
rect 3628 14848 3668 14888
rect 9196 14848 9236 14888
rect 9580 14848 9620 14888
rect 19852 14764 19892 14804
rect 1228 14680 1268 14720
rect 2476 14680 2516 14720
rect 3052 14680 3092 14720
rect 3340 14680 3380 14720
rect 3532 14680 3572 14720
rect 3724 14680 3764 14720
rect 3820 14680 3860 14720
rect 4012 14680 4052 14720
rect 5260 14680 5300 14720
rect 5644 14680 5684 14720
rect 5836 14680 5876 14720
rect 5932 14680 5972 14720
rect 6700 14680 6740 14720
rect 7948 14680 7988 14720
rect 8524 14680 8564 14720
rect 8812 14680 8852 14720
rect 9388 14680 9428 14720
rect 9580 14680 9620 14720
rect 9772 14680 9812 14720
rect 10060 14680 10100 14720
rect 10348 14680 10388 14720
rect 10444 14680 10484 14720
rect 10828 14680 10868 14720
rect 10924 14680 10964 14720
rect 11404 14680 11444 14720
rect 11884 14685 11924 14725
rect 13420 14680 13460 14720
rect 13516 14680 13556 14720
rect 13900 14680 13940 14720
rect 13996 14680 14036 14720
rect 14476 14680 14516 14720
rect 15004 14689 15044 14729
rect 15532 14680 15572 14720
rect 16780 14680 16820 14720
rect 16972 14680 17012 14720
rect 17068 14680 17108 14720
rect 17260 14680 17300 14720
rect 17452 14680 17492 14720
rect 17548 14680 17588 14720
rect 17740 14680 17780 14720
rect 18988 14680 19028 14720
rect 19372 14680 19412 14720
rect 19468 14680 19508 14720
rect 19660 14680 19700 14720
rect 3244 14596 3284 14636
rect 8908 14596 8948 14636
rect 12076 14596 12116 14636
rect 15340 14596 15380 14636
rect 5740 14512 5780 14552
rect 9964 14512 10004 14552
rect 15148 14512 15188 14552
rect 19564 14512 19604 14552
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 3148 14176 3188 14216
rect 5356 14176 5396 14216
rect 5836 14176 5876 14216
rect 8044 14176 8084 14216
rect 8236 14176 8276 14216
rect 11404 14176 11444 14216
rect 13036 14176 13076 14216
rect 17548 14176 17588 14216
rect 18028 14176 18068 14216
rect 20236 14176 20276 14216
rect 15148 14092 15188 14132
rect 1708 14008 1748 14048
rect 2956 14008 2996 14048
rect 3532 14008 3572 14048
rect 3628 14008 3668 14048
rect 3724 14008 3764 14048
rect 3820 14008 3860 14048
rect 4012 14008 4052 14048
rect 4396 14008 4436 14048
rect 4876 14008 4916 14048
rect 4972 14008 5012 14048
rect 5164 14008 5204 14048
rect 5260 14008 5300 14048
rect 5417 13993 5457 14033
rect 6028 14008 6068 14048
rect 6124 14008 6164 14048
rect 6412 14008 6452 14048
rect 6604 14008 6644 14048
rect 7852 14008 7892 14048
rect 8428 14008 8468 14048
rect 9676 14008 9716 14048
rect 9964 14008 10004 14048
rect 11212 14008 11252 14048
rect 11596 14008 11636 14048
rect 12844 14008 12884 14048
rect 13420 14008 13460 14048
rect 13516 14008 13556 14048
rect 14476 14008 14516 14048
rect 14956 14003 14996 14043
rect 15820 14008 15860 14048
rect 15916 14008 15956 14048
rect 16876 14008 16916 14048
rect 17356 14003 17396 14043
rect 17740 14008 17780 14048
rect 17836 14008 17876 14048
rect 18412 14008 18452 14048
rect 19660 14008 19700 14048
rect 4108 13924 4148 13964
rect 4300 13924 4340 13964
rect 6316 13924 6356 13964
rect 13900 13924 13940 13964
rect 13996 13924 14036 13964
rect 16300 13924 16340 13964
rect 16396 13924 16436 13964
rect 20044 13924 20084 13964
rect 4204 13840 4244 13880
rect 4684 13840 4724 13880
rect 8044 13756 8084 13796
rect 8236 13756 8276 13796
rect 19852 13756 19892 13796
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 3148 13420 3188 13460
rect 7180 13420 7220 13460
rect 15916 13420 15956 13460
rect 16876 13420 16916 13460
rect 20236 13420 20276 13460
rect 3628 13336 3668 13376
rect 4684 13336 4724 13376
rect 11596 13336 11636 13376
rect 19084 13336 19124 13376
rect 20044 13252 20084 13292
rect 1708 13168 1748 13208
rect 2956 13168 2996 13208
rect 3916 13168 3956 13208
rect 4012 13168 4052 13208
rect 4300 13168 4340 13208
rect 5164 13168 5204 13208
rect 5260 13168 5300 13208
rect 5644 13168 5684 13208
rect 5740 13168 5780 13208
rect 6220 13168 6260 13208
rect 6700 13182 6740 13222
rect 7084 13157 7124 13197
rect 7564 13168 7604 13208
rect 7660 13168 7700 13208
rect 7852 13168 7892 13208
rect 7948 13168 7988 13208
rect 8140 13168 8180 13208
rect 8332 13168 8372 13208
rect 9580 13168 9620 13208
rect 9964 13168 10004 13208
rect 11212 13168 11252 13208
rect 12940 13168 12980 13208
rect 13036 13168 13076 13208
rect 13420 13168 13460 13208
rect 13516 13168 13556 13208
rect 13996 13168 14036 13208
rect 14476 13173 14516 13213
rect 15244 13168 15284 13208
rect 15532 13168 15572 13208
rect 15628 13168 15668 13208
rect 16204 13168 16244 13208
rect 16492 13168 16532 13208
rect 16588 13168 16628 13208
rect 17356 13168 17396 13208
rect 18604 13168 18644 13208
rect 19372 13168 19412 13208
rect 19468 13168 19508 13208
rect 19756 13168 19796 13208
rect 6892 13084 6932 13124
rect 11404 13084 11444 13124
rect 14668 13084 14708 13124
rect 3148 13000 3188 13040
rect 7372 13000 7412 13040
rect 8140 13000 8180 13040
rect 9772 13000 9812 13040
rect 18796 13000 18836 13040
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 10540 12664 10580 12704
rect 14476 12664 14516 12704
rect 17356 12664 17396 12704
rect 17932 12664 17972 12704
rect 3628 12580 3668 12620
rect 4876 12580 4916 12620
rect 6988 12580 7028 12620
rect 9004 12580 9044 12620
rect 12556 12580 12596 12620
rect 15340 12580 15380 12620
rect 20236 12580 20276 12620
rect 1228 12496 1268 12536
rect 1420 12496 1460 12536
rect 1516 12496 1556 12536
rect 1708 12496 1748 12536
rect 2956 12496 2996 12536
rect 3340 12496 3380 12536
rect 3436 12496 3476 12536
rect 3532 12496 3572 12536
rect 3820 12496 3860 12536
rect 3916 12496 3956 12536
rect 4012 12496 4052 12536
rect 4108 12496 4148 12536
rect 4972 12496 5012 12536
rect 5260 12496 5300 12536
rect 5644 12496 5684 12536
rect 5740 12496 5780 12536
rect 5932 12496 5972 12536
rect 6124 12496 6164 12536
rect 6412 12496 6452 12536
rect 7276 12496 7316 12536
rect 7372 12496 7412 12536
rect 7852 12496 7892 12536
rect 8332 12496 8372 12536
rect 8812 12482 8852 12522
rect 10252 12496 10292 12536
rect 10348 12496 10388 12536
rect 10828 12496 10868 12536
rect 10924 12496 10964 12536
rect 11404 12496 11444 12536
rect 11884 12496 11924 12536
rect 12364 12482 12404 12522
rect 13036 12496 13076 12536
rect 14284 12496 14324 12536
rect 14860 12496 14900 12536
rect 14956 12496 14996 12536
rect 15148 12496 15188 12536
rect 15532 12482 15572 12522
rect 16012 12496 16052 12536
rect 16492 12496 16532 12536
rect 16972 12496 17012 12536
rect 17068 12496 17108 12536
rect 17644 12496 17684 12536
rect 17740 12496 17780 12536
rect 18508 12496 18548 12536
rect 18604 12496 18644 12536
rect 19564 12496 19604 12536
rect 20044 12491 20084 12531
rect 7756 12412 7796 12452
rect 11308 12412 11348 12452
rect 16588 12412 16628 12452
rect 18988 12412 19028 12452
rect 19084 12412 19124 12452
rect 1420 12328 1460 12368
rect 4588 12328 4628 12368
rect 5932 12328 5972 12368
rect 6604 12328 6644 12368
rect 9196 12328 9236 12368
rect 15148 12328 15188 12368
rect 3148 12244 3188 12284
rect 6124 12244 6164 12284
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 3148 11908 3188 11948
rect 6412 11908 6452 11948
rect 6892 11908 6932 11948
rect 9004 11908 9044 11948
rect 10636 11908 10676 11948
rect 12268 11908 12308 11948
rect 17932 11908 17972 11948
rect 20140 11908 20180 11948
rect 3436 11824 3476 11864
rect 3724 11824 3764 11864
rect 4300 11824 4340 11864
rect 4684 11824 4724 11864
rect 1228 11656 1268 11696
rect 1420 11656 1460 11696
rect 1516 11656 1556 11696
rect 1708 11656 1748 11696
rect 2956 11656 2996 11696
rect 3340 11656 3380 11696
rect 3628 11656 3668 11696
rect 3724 11656 3764 11696
rect 3916 11656 3956 11696
rect 4108 11656 4148 11696
rect 4204 11656 4244 11696
rect 4396 11656 4436 11696
rect 4972 11656 5012 11696
rect 6220 11656 6260 11696
rect 6604 11656 6644 11696
rect 6892 11656 6932 11696
rect 7084 11656 7124 11696
rect 7564 11656 7604 11696
rect 8812 11656 8852 11696
rect 10060 11656 10100 11696
rect 10156 11656 10196 11696
rect 10348 11656 10388 11696
rect 10636 11656 10676 11696
rect 10828 11656 10868 11696
rect 12076 11656 12116 11696
rect 13900 11656 13940 11696
rect 15148 11656 15188 11696
rect 15724 11656 15764 11696
rect 16972 11656 17012 11696
rect 17164 11656 17204 11696
rect 17260 11656 17300 11696
rect 17356 11656 17396 11696
rect 17932 11656 17972 11696
rect 18220 11656 18260 11696
rect 18700 11656 18740 11696
rect 19948 11656 19988 11696
rect 9196 11572 9236 11612
rect 15340 11572 15380 11612
rect 1324 11488 1364 11528
rect 6700 11488 6740 11528
rect 9868 11488 9908 11528
rect 15532 11488 15572 11528
rect 17452 11488 17492 11528
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 13036 11194 13076 11234
rect 2668 11152 2708 11192
rect 4684 11152 4724 11192
rect 6124 11152 6164 11192
rect 16972 11152 17012 11192
rect 17740 11152 17780 11192
rect 8620 11068 8660 11108
rect 11020 11068 11060 11108
rect 15052 11068 15092 11108
rect 20140 11068 20180 11108
rect 1228 10984 1268 11024
rect 2476 10984 2516 11024
rect 2860 10984 2900 11024
rect 4108 10984 4148 11024
rect 5164 10984 5204 11024
rect 5452 10984 5492 11024
rect 5644 10984 5684 11024
rect 5836 10984 5876 11024
rect 5932 10984 5972 11024
rect 6316 10984 6356 11024
rect 6412 10984 6452 11024
rect 6700 10984 6740 11024
rect 7180 10984 7220 11024
rect 8428 10984 8468 11024
rect 9196 10984 9236 11024
rect 9388 10984 9428 11024
rect 9580 10984 9620 11024
rect 10828 10984 10868 11024
rect 11308 10984 11348 11024
rect 11404 10984 11444 11024
rect 11884 10984 11924 11024
rect 12364 10984 12404 11024
rect 12844 10970 12884 11010
rect 13324 10984 13364 11024
rect 13420 10984 13460 11024
rect 13804 10984 13844 11024
rect 14380 10984 14420 11024
rect 14860 10970 14900 11010
rect 15436 10984 15476 11024
rect 15628 10984 15668 11024
rect 15916 10984 15956 11024
rect 16204 10984 16244 11024
rect 16300 10984 16340 11024
rect 16780 10984 16820 11024
rect 16876 10984 16916 11024
rect 17068 10984 17108 11024
rect 17260 10984 17300 11024
rect 17356 10984 17396 11024
rect 17452 10984 17492 11024
rect 17548 10984 17588 11024
rect 17932 10984 17972 11024
rect 18028 10984 18068 11024
rect 18412 10984 18452 11024
rect 18508 10984 18548 11024
rect 18892 10984 18932 11024
rect 19468 10984 19508 11024
rect 11788 10900 11828 10940
rect 13900 10900 13940 10940
rect 18988 10900 19028 10940
rect 19996 10942 20036 10982
rect 5452 10816 5492 10856
rect 6892 10816 6932 10856
rect 15436 10816 15476 10856
rect 16588 10816 16628 10856
rect 4300 10732 4340 10772
rect 5644 10732 5684 10772
rect 6604 10732 6644 10772
rect 9292 10732 9332 10772
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 2668 10396 2708 10436
rect 3436 10396 3476 10436
rect 12844 10396 12884 10436
rect 14764 10396 14804 10436
rect 17164 10396 17204 10436
rect 3820 10312 3860 10352
rect 4588 10312 4628 10352
rect 6988 10312 7028 10352
rect 9196 10312 9236 10352
rect 10828 10312 10868 10352
rect 3724 10228 3764 10268
rect 3916 10228 3956 10268
rect 18316 10228 18356 10268
rect 1228 10144 1268 10184
rect 2476 10144 2516 10184
rect 2860 10144 2900 10184
rect 3148 10144 3188 10184
rect 3436 10144 3476 10184
rect 3628 10144 3668 10184
rect 4012 10144 4052 10184
rect 4204 10144 4244 10184
rect 4396 10144 4436 10184
rect 4588 10144 4628 10184
rect 4780 10144 4820 10184
rect 4876 10144 4916 10184
rect 5159 10144 5199 10184
rect 5260 10144 5300 10184
rect 5356 10144 5396 10184
rect 5548 10144 5588 10184
rect 5644 10144 5684 10184
rect 6028 10144 6068 10184
rect 6316 10144 6356 10184
rect 6988 10144 7028 10184
rect 7084 10144 7124 10184
rect 7276 10144 7316 10184
rect 7564 10144 7604 10184
rect 8812 10144 8852 10184
rect 9484 10144 9524 10184
rect 9580 10144 9620 10184
rect 9772 10144 9812 10184
rect 10156 10144 10196 10184
rect 10444 10144 10484 10184
rect 10540 10144 10580 10184
rect 11020 10144 11060 10184
rect 11212 10144 11252 10184
rect 11404 10144 11444 10184
rect 12652 10144 12692 10184
rect 13324 10144 13364 10184
rect 14572 10144 14612 10184
rect 14956 10144 14996 10184
rect 15052 10144 15092 10184
rect 15724 10144 15764 10184
rect 16972 10144 17012 10184
rect 17740 10144 17780 10184
rect 17836 10144 17876 10184
rect 17932 10144 17972 10184
rect 18028 10144 18068 10184
rect 18220 10144 18260 10184
rect 18509 10129 18549 10169
rect 18700 10144 18740 10184
rect 19948 10144 19988 10184
rect 2956 10060 2996 10100
rect 4300 10060 4340 10100
rect 9004 10060 9044 10100
rect 11116 10060 11156 10100
rect 20140 10060 20180 10100
rect 5356 9976 5396 10016
rect 6124 9976 6164 10016
rect 6700 9976 6740 10016
rect 9772 9976 9812 10016
rect 15244 9976 15284 10016
rect 17356 9976 17396 10016
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 3052 9640 3092 9680
rect 4684 9682 4724 9722
rect 5644 9640 5684 9680
rect 6700 9640 6740 9680
rect 8716 9640 8756 9680
rect 9196 9640 9236 9680
rect 13132 9640 13172 9680
rect 14476 9640 14516 9680
rect 16780 9640 16820 9680
rect 19084 9640 19124 9680
rect 1612 9472 1652 9512
rect 2860 9472 2900 9512
rect 3716 9471 3756 9511
rect 4012 9472 4052 9512
rect 4300 9472 4340 9512
rect 4396 9472 4436 9512
rect 4876 9472 4916 9512
rect 4972 9472 5012 9512
rect 5068 9472 5108 9512
rect 5164 9472 5204 9512
rect 5548 9472 5588 9512
rect 5836 9472 5876 9512
rect 6028 9472 6068 9512
rect 6220 9458 6260 9498
rect 6316 9472 6356 9512
rect 6988 9472 7028 9512
rect 7084 9472 7124 9512
rect 7468 9430 7508 9470
rect 7564 9472 7604 9512
rect 8044 9472 8084 9512
rect 8524 9458 8564 9498
rect 9676 9472 9716 9512
rect 10924 9472 10964 9512
rect 11692 9472 11732 9512
rect 12940 9472 12980 9512
rect 13612 9472 13652 9512
rect 13708 9472 13748 9512
rect 13804 9472 13844 9512
rect 13900 9472 13940 9512
rect 14284 9472 14324 9512
rect 14380 9472 14420 9512
rect 14572 9472 14612 9512
rect 14668 9472 14708 9512
rect 14823 9472 14863 9512
rect 15340 9472 15380 9512
rect 16588 9472 16628 9512
rect 17644 9472 17684 9512
rect 18892 9472 18932 9512
rect 19367 9472 19407 9512
rect 19468 9472 19508 9512
rect 19564 9472 19604 9512
rect 19756 9472 19796 9512
rect 19852 9472 19892 9512
rect 20044 9472 20084 9512
rect 20236 9472 20276 9512
rect 20140 9388 20180 9428
rect 3628 9304 3668 9344
rect 6028 9304 6068 9344
rect 15052 9304 15092 9344
rect 17356 9304 17396 9344
rect 3052 9220 3092 9260
rect 11116 9220 11156 9260
rect 19084 9220 19124 9260
rect 19852 9220 19892 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 3916 8884 3956 8924
rect 6316 8884 6356 8924
rect 8332 8884 8372 8924
rect 14764 8884 14804 8924
rect 19084 8884 19124 8924
rect 3340 8800 3380 8840
rect 15340 8800 15380 8840
rect 20236 8800 20276 8840
rect 4492 8716 4532 8756
rect 9292 8716 9332 8756
rect 20044 8716 20084 8756
rect 1900 8632 1940 8672
rect 3148 8632 3188 8672
rect 3916 8632 3956 8672
rect 4108 8632 4148 8672
rect 4204 8632 4244 8672
rect 4396 8632 4436 8672
rect 4684 8632 4724 8672
rect 4876 8632 4916 8672
rect 6124 8632 6164 8672
rect 6892 8632 6932 8672
rect 8140 8632 8180 8672
rect 8716 8632 8756 8672
rect 8812 8632 8852 8672
rect 9196 8632 9236 8672
rect 9772 8632 9812 8672
rect 10300 8641 10340 8681
rect 10732 8632 10772 8672
rect 10828 8632 10868 8672
rect 11212 8632 11252 8672
rect 12460 8632 12500 8672
rect 13324 8632 13364 8672
rect 14572 8632 14612 8672
rect 15436 8632 15476 8672
rect 16876 8632 16916 8672
rect 16972 8632 17012 8672
rect 17644 8632 17684 8672
rect 18892 8632 18932 8672
rect 19276 8632 19316 8672
rect 19372 8632 19412 8672
rect 19564 8632 19604 8672
rect 19660 8632 19700 8672
rect 19817 8647 19857 8687
rect 6604 8464 6644 8504
rect 10444 8464 10484 8504
rect 11020 8464 11060 8504
rect 12652 8464 12692 8504
rect 15052 8464 15092 8504
rect 17164 8464 17204 8504
rect 17356 8464 17396 8504
rect 19084 8464 19124 8504
rect 19756 8464 19796 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 3628 8128 3668 8168
rect 3916 8128 3956 8168
rect 8620 8128 8660 8168
rect 10348 8128 10388 8168
rect 14860 8128 14900 8168
rect 19756 8128 19796 8168
rect 20140 8128 20180 8168
rect 12748 8044 12788 8084
rect 2956 7960 2996 8000
rect 3052 7960 3092 8000
rect 3148 7960 3188 8000
rect 3244 7960 3284 8000
rect 3436 7960 3476 8000
rect 3532 7960 3572 8000
rect 3724 7960 3764 8000
rect 3916 7960 3956 8000
rect 4108 7960 4148 8000
rect 4204 7960 4244 8000
rect 4684 7960 4724 8000
rect 4780 7960 4820 8000
rect 4972 7960 5012 8000
rect 7180 7960 7220 8000
rect 8428 7960 8468 8000
rect 8908 7960 8948 8000
rect 10156 7960 10196 8000
rect 11020 7960 11060 8000
rect 11116 7960 11156 8000
rect 12076 7960 12116 8000
rect 12604 7950 12644 7990
rect 13420 7960 13460 8000
rect 14668 7960 14708 8000
rect 17644 7960 17684 8000
rect 18892 7960 18932 8000
rect 19468 7960 19508 8000
rect 19564 7960 19604 8000
rect 19948 7960 19988 8000
rect 20044 7960 20084 8000
rect 20236 7960 20276 8000
rect 11500 7876 11540 7916
rect 11596 7876 11636 7916
rect 4684 7792 4724 7832
rect 6316 7792 6356 7832
rect 6604 7792 6644 7832
rect 15052 7792 15092 7832
rect 17356 7792 17396 7832
rect 19084 7708 19124 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 4492 7372 4532 7412
rect 20236 7372 20276 7412
rect 12364 7288 12404 7328
rect 15052 7288 15092 7328
rect 18796 7288 18836 7328
rect 19276 7288 19316 7328
rect 8812 7204 8852 7244
rect 13132 7204 13172 7244
rect 13228 7204 13268 7244
rect 16012 7204 16052 7244
rect 20044 7204 20084 7244
rect 4204 7120 4244 7160
rect 4492 7120 4532 7160
rect 6508 7120 6548 7160
rect 7756 7120 7796 7160
rect 8236 7120 8276 7160
rect 8332 7120 8372 7160
rect 8716 7120 8756 7160
rect 9292 7120 9332 7160
rect 9820 7129 9860 7169
rect 10924 7120 10964 7160
rect 12172 7120 12212 7160
rect 12652 7120 12692 7160
rect 12748 7120 12788 7160
rect 13708 7120 13748 7160
rect 14188 7125 14228 7165
rect 15436 7120 15476 7160
rect 15532 7120 15572 7160
rect 15916 7120 15956 7160
rect 16492 7120 16532 7160
rect 16972 7125 17012 7165
rect 17356 7120 17396 7160
rect 18604 7120 18644 7160
rect 18988 7120 19028 7160
rect 19180 7120 19220 7160
rect 19276 7120 19316 7160
rect 19756 7120 19796 7160
rect 19852 7120 19892 7160
rect 7948 7036 7988 7076
rect 17164 7036 17204 7076
rect 9964 6952 10004 6992
rect 14380 6952 14420 6992
rect 19564 6952 19604 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 6604 6616 6644 6656
rect 9868 6616 9908 6656
rect 14188 6616 14228 6656
rect 16492 6616 16532 6656
rect 20140 6616 20180 6656
rect 8428 6448 8468 6488
rect 9676 6448 9716 6488
rect 12748 6448 12788 6488
rect 13996 6448 14036 6488
rect 15052 6448 15092 6488
rect 16300 6448 16340 6488
rect 18700 6448 18740 6488
rect 19948 6448 19988 6488
rect 10156 6364 10196 6404
rect 11692 6364 11732 6404
rect 11500 6280 11540 6320
rect 17356 6280 17396 6320
rect 10348 6196 10388 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 14860 5860 14900 5900
rect 6604 5776 6644 5816
rect 15052 5776 15092 5816
rect 13420 5608 13460 5648
rect 14668 5608 14708 5648
rect 19660 5608 19700 5648
rect 19756 5608 19796 5648
rect 17356 5440 17396 5480
rect 19468 5440 19508 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 6604 5104 6644 5144
rect 15052 5104 15092 5144
rect 17356 4768 17396 4808
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 6604 4264 6644 4304
rect 15052 4264 15092 4304
rect 17356 3928 17396 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 6604 3592 6644 3632
rect 15052 3592 15092 3632
rect 17356 3592 17396 3632
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 6892 2836 6932 2876
rect 15052 2752 15092 2792
rect 7084 2668 7124 2708
rect 11404 2668 11444 2708
rect 13804 2668 13844 2708
rect 14380 2668 14420 2708
rect 11596 2416 11636 2456
rect 13996 2416 14036 2456
rect 14572 2416 14612 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 5740 2080 5780 2120
rect 6124 2080 6164 2120
rect 6508 2080 6548 2120
rect 6892 2080 6932 2120
rect 7276 2080 7316 2120
rect 7660 2080 7700 2120
rect 13900 2080 13940 2120
rect 15244 2080 15284 2120
rect 17260 2080 17300 2120
rect 17644 2080 17684 2120
rect 18028 2080 18068 2120
rect 18412 2080 18452 2120
rect 18796 2080 18836 2120
rect 19180 2080 19220 2120
rect 19564 2080 19604 2120
rect 19948 2080 19988 2120
rect 5932 1828 5972 1868
rect 6316 1828 6356 1868
rect 6700 1828 6740 1868
rect 7084 1828 7124 1868
rect 7468 1828 7508 1868
rect 7852 1828 7892 1868
rect 8140 1828 8180 1868
rect 8620 1828 8660 1868
rect 9004 1828 9044 1868
rect 9580 1828 9620 1868
rect 9772 1828 9812 1868
rect 10156 1841 10196 1881
rect 10540 1828 10580 1868
rect 10924 1828 10964 1868
rect 11500 1828 11540 1868
rect 11692 1828 11732 1868
rect 12076 1828 12116 1868
rect 12748 1828 12788 1868
rect 13324 1828 13364 1868
rect 14284 1828 14324 1868
rect 14668 1828 14708 1868
rect 15628 1828 15668 1868
rect 16012 1828 16052 1868
rect 16396 1828 16436 1868
rect 16780 1828 16820 1868
rect 17452 1828 17492 1868
rect 17836 1828 17876 1868
rect 18220 1828 18260 1868
rect 18604 1828 18644 1868
rect 18988 1828 19028 1868
rect 19372 1828 19412 1868
rect 19756 1828 19796 1868
rect 20121 1825 20161 1865
rect 9196 1744 9236 1784
rect 15436 1744 15476 1784
rect 8332 1660 8372 1700
rect 8812 1660 8852 1700
rect 9388 1660 9428 1700
rect 9964 1660 10004 1700
rect 10348 1660 10388 1700
rect 10732 1660 10772 1700
rect 11116 1660 11156 1700
rect 11308 1660 11348 1700
rect 11884 1660 11924 1700
rect 12268 1660 12308 1700
rect 12940 1660 12980 1700
rect 13132 1660 13172 1700
rect 14092 1660 14132 1700
rect 14476 1660 14516 1700
rect 15820 1660 15860 1700
rect 16204 1660 16244 1700
rect 16588 1660 16628 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 6508 1240 6548 1280
rect 14188 1240 14228 1280
rect 18028 1240 18068 1280
rect 18412 1240 18452 1280
rect 18796 1240 18836 1280
rect 6700 1156 6740 1196
rect 6892 1156 6932 1196
rect 9388 1156 9428 1196
rect 10348 1156 10388 1196
rect 11116 1156 11156 1196
rect 11596 1156 11636 1196
rect 13036 1156 13076 1196
rect 13420 1156 13460 1196
rect 13804 1156 13844 1196
rect 14572 1156 14612 1196
rect 14956 1156 14996 1196
rect 15340 1156 15380 1196
rect 15724 1156 15764 1196
rect 16108 1156 16148 1196
rect 18220 1156 18260 1196
rect 18604 1156 18644 1196
rect 18988 1156 19028 1196
rect 19372 1156 19412 1196
rect 7084 904 7124 944
rect 9196 904 9236 944
rect 10540 904 10580 944
rect 11308 904 11348 944
rect 11788 904 11828 944
rect 13228 904 13268 944
rect 13612 904 13652 944
rect 14380 904 14420 944
rect 14764 904 14804 944
rect 15148 904 15188 944
rect 15532 904 15572 944
rect 15916 904 15956 944
rect 19180 904 19220 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal2 >>
rect 1784 85936 1864 86016
rect 1976 85936 2056 86016
rect 2168 85936 2248 86016
rect 2360 85936 2440 86016
rect 2552 85936 2632 86016
rect 2744 85936 2824 86016
rect 2936 85936 3016 86016
rect 3128 85936 3208 86016
rect 3320 85936 3400 86016
rect 3512 85936 3592 86016
rect 3704 85936 3784 86016
rect 3896 85936 3976 86016
rect 4088 85936 4168 86016
rect 4280 85936 4360 86016
rect 4472 85936 4552 86016
rect 4664 85936 4744 86016
rect 4856 85936 4936 86016
rect 5048 85936 5128 86016
rect 5240 85936 5320 86016
rect 5432 85936 5512 86016
rect 5624 85936 5704 86016
rect 5816 85936 5896 86016
rect 6008 85936 6088 86016
rect 6200 85936 6280 86016
rect 6392 85936 6472 86016
rect 6584 85936 6664 86016
rect 6776 85936 6856 86016
rect 6968 85936 7048 86016
rect 7160 85936 7240 86016
rect 7352 85936 7432 86016
rect 7544 85936 7624 86016
rect 7736 85936 7816 86016
rect 7928 85936 8008 86016
rect 8120 85936 8200 86016
rect 8312 85936 8392 86016
rect 8504 85936 8584 86016
rect 8696 85936 8776 86016
rect 8888 85936 8968 86016
rect 9080 85936 9160 86016
rect 9272 85936 9352 86016
rect 9464 85936 9544 86016
rect 9656 85936 9736 86016
rect 9848 85936 9928 86016
rect 10040 85936 10120 86016
rect 10232 85936 10312 86016
rect 10424 85936 10504 86016
rect 10616 85936 10696 86016
rect 10808 85936 10888 86016
rect 11000 85936 11080 86016
rect 11192 85936 11272 86016
rect 11384 85936 11464 86016
rect 11576 85936 11656 86016
rect 11768 85936 11848 86016
rect 11960 85936 12040 86016
rect 12152 85936 12232 86016
rect 12344 85936 12424 86016
rect 12536 85936 12616 86016
rect 12728 85936 12808 86016
rect 12920 85936 13000 86016
rect 13112 85936 13192 86016
rect 13304 85936 13384 86016
rect 13496 85936 13576 86016
rect 13688 85936 13768 86016
rect 13880 85936 13960 86016
rect 14072 85936 14152 86016
rect 14264 85936 14344 86016
rect 14456 85936 14536 86016
rect 14648 85936 14728 86016
rect 14840 85936 14920 86016
rect 15032 85936 15112 86016
rect 15224 85936 15304 86016
rect 15416 85936 15496 86016
rect 15608 85936 15688 86016
rect 15800 85936 15880 86016
rect 15992 85936 16072 86016
rect 16184 85936 16264 86016
rect 16376 85936 16456 86016
rect 16568 85936 16648 86016
rect 16760 85936 16840 86016
rect 16952 85936 17032 86016
rect 17144 85936 17224 86016
rect 17336 85936 17416 86016
rect 17528 85936 17608 86016
rect 17720 85936 17800 86016
rect 17912 85936 17992 86016
rect 18104 85936 18184 86016
rect 18296 85936 18376 86016
rect 18488 85936 18568 86016
rect 18680 85936 18760 86016
rect 18872 85936 18952 86016
rect 19064 85952 19144 86016
rect 19064 85936 19084 85952
rect 1035 85112 1077 85121
rect 1035 85072 1036 85112
rect 1076 85072 1077 85112
rect 1035 85063 1077 85072
rect 171 78560 213 78569
rect 171 78520 172 78560
rect 212 78520 213 78560
rect 171 78511 213 78520
rect 75 66464 117 66473
rect 75 66424 76 66464
rect 116 66424 117 66464
rect 75 66415 117 66424
rect 76 36653 116 66415
rect 172 59837 212 78511
rect 267 73856 309 73865
rect 267 73816 268 73856
rect 308 73816 309 73856
rect 267 73807 309 73816
rect 268 61013 308 73807
rect 843 70496 885 70505
rect 843 70456 844 70496
rect 884 70456 885 70496
rect 843 70447 885 70456
rect 844 65549 884 70447
rect 843 65540 885 65549
rect 843 65500 844 65540
rect 884 65500 885 65540
rect 843 65491 885 65500
rect 747 65120 789 65129
rect 747 65080 748 65120
rect 788 65080 789 65120
rect 747 65071 789 65080
rect 267 61004 309 61013
rect 267 60964 268 61004
rect 308 60964 309 61004
rect 267 60955 309 60964
rect 171 59828 213 59837
rect 171 59788 172 59828
rect 212 59788 213 59828
rect 171 59779 213 59788
rect 363 59744 405 59753
rect 363 59704 364 59744
rect 404 59704 405 59744
rect 363 59695 405 59704
rect 171 59072 213 59081
rect 171 59032 172 59072
rect 212 59032 213 59072
rect 171 59023 213 59032
rect 172 46649 212 59023
rect 171 46640 213 46649
rect 171 46600 172 46640
rect 212 46600 213 46640
rect 171 46591 213 46600
rect 364 44465 404 59695
rect 748 50420 788 65071
rect 939 60416 981 60425
rect 939 60376 940 60416
rect 980 60376 981 60416
rect 939 60367 981 60376
rect 940 50420 980 60367
rect 1036 54209 1076 85063
rect 1708 83768 1748 83777
rect 1804 83768 1844 85936
rect 1748 83728 1844 83768
rect 1900 83768 1940 83777
rect 1996 83768 2036 85936
rect 1940 83728 2036 83768
rect 1708 83719 1748 83728
rect 1900 83719 1940 83728
rect 2188 83609 2228 85936
rect 2284 83768 2324 83777
rect 2380 83768 2420 85936
rect 2324 83728 2420 83768
rect 2284 83719 2324 83728
rect 2187 83600 2229 83609
rect 2187 83560 2188 83600
rect 2228 83560 2229 83600
rect 2187 83551 2229 83560
rect 1515 83516 1557 83525
rect 1515 83476 1516 83516
rect 1556 83476 1557 83516
rect 1515 83467 1557 83476
rect 2091 83516 2133 83525
rect 2476 83516 2516 83525
rect 2091 83476 2092 83516
rect 2132 83476 2133 83516
rect 2091 83467 2133 83476
rect 2284 83476 2476 83516
rect 1516 83382 1556 83467
rect 2092 83382 2132 83467
rect 2284 76880 2324 83476
rect 2476 83467 2516 83476
rect 2572 82844 2612 85936
rect 2668 83768 2708 83777
rect 2764 83768 2804 85936
rect 2708 83728 2804 83768
rect 2668 83719 2708 83728
rect 2667 83600 2709 83609
rect 2667 83560 2668 83600
rect 2708 83560 2709 83600
rect 2956 83600 2996 85936
rect 3052 83768 3092 83777
rect 3148 83768 3188 85936
rect 3340 83861 3380 85936
rect 3435 84860 3477 84869
rect 3435 84820 3436 84860
rect 3476 84820 3477 84860
rect 3435 84811 3477 84820
rect 3436 84449 3476 84811
rect 3435 84440 3477 84449
rect 3435 84400 3436 84440
rect 3476 84400 3477 84440
rect 3435 84391 3477 84400
rect 3339 83852 3381 83861
rect 3339 83812 3340 83852
rect 3380 83812 3381 83852
rect 3339 83803 3381 83812
rect 3092 83728 3188 83768
rect 3436 83768 3476 83777
rect 3532 83768 3572 85936
rect 3724 84869 3764 85936
rect 3723 84860 3765 84869
rect 3723 84820 3724 84860
rect 3764 84820 3765 84860
rect 3916 84860 3956 85936
rect 4108 85037 4148 85936
rect 4107 85028 4149 85037
rect 4107 84988 4108 85028
rect 4148 84988 4149 85028
rect 4107 84979 4149 84988
rect 3916 84820 4148 84860
rect 3723 84811 3765 84820
rect 3688 84692 4056 84701
rect 3728 84652 3770 84692
rect 3810 84652 3852 84692
rect 3892 84652 3934 84692
rect 3974 84652 4016 84692
rect 3688 84643 4056 84652
rect 4108 84524 4148 84820
rect 4300 84692 4340 85936
rect 4395 85028 4437 85037
rect 4395 84988 4396 85028
rect 4436 84988 4437 85028
rect 4395 84979 4437 84988
rect 3476 83728 3572 83768
rect 3820 84484 4148 84524
rect 4204 84652 4340 84692
rect 3820 83768 3860 84484
rect 4107 83852 4149 83861
rect 4107 83812 4108 83852
rect 4148 83812 4149 83852
rect 4107 83803 4149 83812
rect 3052 83719 3092 83728
rect 3436 83719 3476 83728
rect 3820 83719 3860 83728
rect 3148 83644 3380 83684
rect 3148 83600 3188 83644
rect 2956 83560 3188 83600
rect 3340 83600 3380 83644
rect 3340 83560 3476 83600
rect 2667 83551 2709 83560
rect 2668 83012 2708 83551
rect 2859 83516 2901 83525
rect 2859 83476 2860 83516
rect 2900 83476 2901 83516
rect 2859 83467 2901 83476
rect 3244 83516 3284 83525
rect 3284 83476 3380 83516
rect 3244 83467 3284 83476
rect 2860 83382 2900 83467
rect 3052 83012 3092 83021
rect 2668 82963 2708 82972
rect 2764 82972 3052 83012
rect 2764 82844 2804 82972
rect 3052 82963 3092 82972
rect 2572 82804 2804 82844
rect 2859 82844 2901 82853
rect 2859 82804 2860 82844
rect 2900 82804 2901 82844
rect 2859 82795 2901 82804
rect 3243 82844 3285 82853
rect 3243 82804 3244 82844
rect 3284 82804 3285 82844
rect 3243 82795 3285 82804
rect 2860 82710 2900 82795
rect 3244 82710 3284 82795
rect 2379 81164 2421 81173
rect 2379 81124 2380 81164
rect 2420 81124 2421 81164
rect 2379 81115 2421 81124
rect 1612 76840 2324 76880
rect 1515 72764 1557 72773
rect 1515 72724 1516 72764
rect 1556 72724 1557 72764
rect 1515 72715 1557 72724
rect 1323 72344 1365 72353
rect 1323 72304 1324 72344
rect 1364 72304 1365 72344
rect 1323 72295 1365 72304
rect 1228 72176 1268 72185
rect 1324 72176 1364 72295
rect 1268 72136 1364 72176
rect 1228 72127 1268 72136
rect 1516 71504 1556 72715
rect 1516 71455 1556 71464
rect 1323 70412 1365 70421
rect 1323 70372 1324 70412
rect 1364 70372 1365 70412
rect 1323 70363 1365 70372
rect 1228 69992 1268 70001
rect 1324 69992 1364 70363
rect 1268 69952 1364 69992
rect 1515 69992 1557 70001
rect 1515 69952 1516 69992
rect 1556 69952 1557 69992
rect 1228 69943 1268 69952
rect 1515 69943 1557 69952
rect 1516 68480 1556 69943
rect 1324 67640 1364 67649
rect 1324 67397 1364 67600
rect 1323 67388 1365 67397
rect 1323 67348 1324 67388
rect 1364 67348 1365 67388
rect 1323 67339 1365 67348
rect 1227 66968 1269 66977
rect 1227 66928 1228 66968
rect 1268 66928 1269 66968
rect 1227 66919 1269 66928
rect 1228 66834 1268 66919
rect 1419 66128 1461 66137
rect 1419 66088 1420 66128
rect 1460 66088 1461 66128
rect 1419 66079 1461 66088
rect 1420 65994 1460 66079
rect 1131 64448 1173 64457
rect 1131 64408 1132 64448
rect 1172 64408 1173 64448
rect 1131 64399 1173 64408
rect 1035 54200 1077 54209
rect 1035 54160 1036 54200
rect 1076 54160 1077 54200
rect 1035 54151 1077 54160
rect 748 50380 884 50420
rect 940 50380 1076 50420
rect 363 44456 405 44465
rect 363 44416 364 44456
rect 404 44416 405 44456
rect 363 44407 405 44416
rect 747 41768 789 41777
rect 747 41728 748 41768
rect 788 41728 789 41768
rect 747 41719 789 41728
rect 171 38492 213 38501
rect 171 38452 172 38492
rect 212 38452 213 38492
rect 171 38443 213 38452
rect 75 36644 117 36653
rect 75 36604 76 36644
rect 116 36604 117 36644
rect 75 36595 117 36604
rect 75 35552 117 35561
rect 75 35512 76 35552
rect 116 35512 117 35552
rect 75 35503 117 35512
rect 76 10361 116 35503
rect 172 17417 212 38443
rect 651 37316 693 37325
rect 651 37276 652 37316
rect 692 37276 693 37316
rect 651 37267 693 37276
rect 652 31529 692 37267
rect 748 33797 788 41719
rect 844 40433 884 50380
rect 939 41432 981 41441
rect 939 41392 940 41432
rect 980 41392 981 41432
rect 939 41383 981 41392
rect 843 40424 885 40433
rect 843 40384 844 40424
rect 884 40384 885 40424
rect 843 40375 885 40384
rect 843 39920 885 39929
rect 843 39880 844 39920
rect 884 39880 885 39920
rect 843 39871 885 39880
rect 747 33788 789 33797
rect 747 33748 748 33788
rect 788 33748 789 33788
rect 747 33739 789 33748
rect 651 31520 693 31529
rect 651 31480 652 31520
rect 692 31480 693 31520
rect 651 31471 693 31480
rect 267 29252 309 29261
rect 267 29212 268 29252
rect 308 29212 309 29252
rect 267 29203 309 29212
rect 268 20105 308 29203
rect 267 20096 309 20105
rect 267 20056 268 20096
rect 308 20056 309 20096
rect 267 20047 309 20056
rect 459 19592 501 19601
rect 459 19552 460 19592
rect 500 19552 501 19592
rect 459 19543 501 19552
rect 171 17408 213 17417
rect 171 17368 172 17408
rect 212 17368 213 17408
rect 171 17359 213 17368
rect 363 16568 405 16577
rect 363 16528 364 16568
rect 404 16528 405 16568
rect 363 16519 405 16528
rect 75 10352 117 10361
rect 75 10312 76 10352
rect 116 10312 117 10352
rect 75 10303 117 10312
rect 364 8681 404 16519
rect 460 11369 500 19543
rect 844 15065 884 39871
rect 940 15485 980 41383
rect 1036 35888 1076 50380
rect 1132 38240 1172 64399
rect 1228 62432 1268 62441
rect 1228 62348 1268 62392
rect 1323 62348 1365 62357
rect 1228 62308 1324 62348
rect 1364 62308 1365 62348
rect 1323 62299 1365 62308
rect 1516 61517 1556 68440
rect 1612 61937 1652 76840
rect 1995 74528 2037 74537
rect 1995 74488 1996 74528
rect 2036 74488 2037 74528
rect 1995 74479 2037 74488
rect 1899 73184 1941 73193
rect 1899 73144 1900 73184
rect 1940 73144 1941 73184
rect 1899 73135 1941 73144
rect 1803 65540 1845 65549
rect 1803 65500 1804 65540
rect 1844 65500 1845 65540
rect 1803 65491 1845 65500
rect 1707 64112 1749 64121
rect 1707 64072 1708 64112
rect 1748 64072 1749 64112
rect 1707 64063 1749 64072
rect 1708 63944 1748 64063
rect 1708 63895 1748 63904
rect 1707 62852 1749 62861
rect 1707 62812 1708 62852
rect 1748 62812 1749 62852
rect 1707 62803 1749 62812
rect 1708 62357 1748 62803
rect 1707 62348 1749 62357
rect 1707 62308 1708 62348
rect 1748 62308 1749 62348
rect 1707 62299 1749 62308
rect 1611 61928 1653 61937
rect 1611 61888 1612 61928
rect 1652 61888 1653 61928
rect 1611 61879 1653 61888
rect 1515 61508 1557 61517
rect 1515 61468 1516 61508
rect 1556 61468 1557 61508
rect 1515 61459 1557 61468
rect 1420 60920 1460 60929
rect 1420 60593 1460 60880
rect 1419 60584 1461 60593
rect 1419 60544 1420 60584
rect 1460 60544 1461 60584
rect 1419 60535 1461 60544
rect 1228 60080 1268 60089
rect 1268 60040 1364 60080
rect 1228 60031 1268 60040
rect 1324 59417 1364 60040
rect 1323 59408 1365 59417
rect 1323 59368 1324 59408
rect 1364 59368 1365 59408
rect 1323 59359 1365 59368
rect 1516 59240 1556 61459
rect 1611 60836 1653 60845
rect 1611 60796 1612 60836
rect 1652 60796 1653 60836
rect 1611 60787 1653 60796
rect 1324 59200 1556 59240
rect 1324 57896 1364 59200
rect 1612 59072 1652 60787
rect 1420 59032 1652 59072
rect 1420 58568 1460 59032
rect 1420 57980 1460 58528
rect 1420 57940 1652 57980
rect 1324 57847 1364 57856
rect 1515 57644 1557 57653
rect 1515 57604 1516 57644
rect 1556 57604 1557 57644
rect 1515 57595 1557 57604
rect 1324 57056 1364 57065
rect 1324 56645 1364 57016
rect 1323 56636 1365 56645
rect 1323 56596 1324 56636
rect 1364 56596 1365 56636
rect 1323 56587 1365 56596
rect 1324 55721 1364 56587
rect 1419 56048 1461 56057
rect 1419 56008 1420 56048
rect 1460 56008 1461 56048
rect 1419 55999 1461 56008
rect 1323 55712 1365 55721
rect 1323 55672 1324 55712
rect 1364 55672 1365 55712
rect 1323 55663 1365 55672
rect 1324 55544 1364 55553
rect 1324 55460 1364 55504
rect 1420 55460 1460 55999
rect 1324 55420 1460 55460
rect 1324 54284 1364 55420
rect 1419 54956 1461 54965
rect 1419 54916 1420 54956
rect 1460 54916 1461 54956
rect 1419 54907 1461 54916
rect 1420 54872 1460 54907
rect 1420 54377 1460 54832
rect 1419 54368 1461 54377
rect 1419 54328 1420 54368
rect 1460 54328 1461 54368
rect 1419 54319 1461 54328
rect 1228 54244 1364 54284
rect 1228 53705 1268 54244
rect 1516 54200 1556 57595
rect 1612 57476 1652 57940
rect 1708 57653 1748 62299
rect 1707 57644 1749 57653
rect 1707 57604 1708 57644
rect 1748 57604 1749 57644
rect 1707 57595 1749 57604
rect 1612 57436 1748 57476
rect 1611 56552 1653 56561
rect 1611 56512 1612 56552
rect 1652 56512 1653 56552
rect 1611 56503 1653 56512
rect 1612 56384 1652 56503
rect 1612 55049 1652 56344
rect 1611 55040 1653 55049
rect 1611 55000 1612 55040
rect 1652 55000 1653 55040
rect 1611 54991 1653 55000
rect 1324 54160 1556 54200
rect 1227 53696 1269 53705
rect 1227 53656 1228 53696
rect 1268 53656 1269 53696
rect 1227 53647 1269 53656
rect 1324 53369 1364 54160
rect 1420 54032 1460 54041
rect 1460 53992 1652 54032
rect 1420 53983 1460 53992
rect 1228 53360 1268 53369
rect 1323 53360 1365 53369
rect 1268 53320 1324 53360
rect 1364 53320 1365 53360
rect 1228 53311 1268 53320
rect 1323 53311 1365 53320
rect 1324 53226 1364 53311
rect 1515 52856 1557 52865
rect 1515 52816 1516 52856
rect 1556 52816 1557 52856
rect 1515 52807 1557 52816
rect 1419 52604 1461 52613
rect 1419 52564 1420 52604
rect 1460 52564 1461 52604
rect 1419 52555 1461 52564
rect 1420 52520 1460 52555
rect 1420 52469 1460 52480
rect 1419 51848 1461 51857
rect 1419 51808 1420 51848
rect 1460 51808 1461 51848
rect 1419 51799 1461 51808
rect 1228 51008 1268 51017
rect 1228 50924 1268 50968
rect 1323 50924 1365 50933
rect 1228 50884 1324 50924
rect 1364 50884 1365 50924
rect 1323 50875 1365 50884
rect 1420 50261 1460 51799
rect 1419 50252 1461 50261
rect 1419 50212 1420 50252
rect 1460 50212 1461 50252
rect 1419 50203 1461 50212
rect 1419 49664 1461 49673
rect 1419 49624 1420 49664
rect 1460 49624 1461 49664
rect 1419 49615 1461 49624
rect 1323 48992 1365 49001
rect 1323 48952 1324 48992
rect 1364 48952 1365 48992
rect 1323 48943 1365 48952
rect 1324 48824 1364 48943
rect 1324 48775 1364 48784
rect 1323 48236 1365 48245
rect 1420 48236 1460 49615
rect 1516 49001 1556 52807
rect 1612 50177 1652 53992
rect 1708 50345 1748 57436
rect 1707 50336 1749 50345
rect 1707 50296 1708 50336
rect 1748 50296 1749 50336
rect 1707 50287 1749 50296
rect 1611 50168 1653 50177
rect 1611 50128 1612 50168
rect 1652 50128 1653 50168
rect 1611 50119 1653 50128
rect 1515 48992 1557 49001
rect 1515 48952 1516 48992
rect 1556 48952 1557 48992
rect 1515 48943 1557 48952
rect 1323 48196 1324 48236
rect 1364 48196 1460 48236
rect 1323 48187 1365 48196
rect 1228 47984 1268 47993
rect 1324 47984 1364 48187
rect 1268 47944 1364 47984
rect 1228 47935 1268 47944
rect 1612 46985 1652 50119
rect 1708 47993 1748 50287
rect 1707 47984 1749 47993
rect 1707 47944 1708 47984
rect 1748 47944 1749 47984
rect 1707 47935 1749 47944
rect 1611 46976 1653 46985
rect 1611 46936 1612 46976
rect 1652 46936 1653 46976
rect 1611 46927 1653 46936
rect 1419 46808 1461 46817
rect 1419 46768 1420 46808
rect 1460 46768 1461 46808
rect 1419 46759 1461 46768
rect 1323 46640 1365 46649
rect 1323 46600 1324 46640
rect 1364 46600 1365 46640
rect 1323 46591 1365 46600
rect 1228 46472 1268 46481
rect 1228 45641 1268 46432
rect 1227 45632 1269 45641
rect 1227 45592 1228 45632
rect 1268 45592 1269 45632
rect 1227 45583 1269 45592
rect 1324 42776 1364 46591
rect 1420 45800 1460 46759
rect 1707 46640 1749 46649
rect 1707 46600 1708 46640
rect 1748 46600 1749 46640
rect 1707 46591 1749 46600
rect 1420 45751 1460 45760
rect 1420 42776 1460 42785
rect 1324 42736 1420 42776
rect 1323 41516 1365 41525
rect 1323 41476 1324 41516
rect 1364 41476 1365 41516
rect 1323 41467 1365 41476
rect 1228 39752 1268 39761
rect 1324 39752 1364 41467
rect 1268 39712 1364 39752
rect 1228 39703 1268 39712
rect 1228 38240 1268 38249
rect 1132 38200 1228 38240
rect 1228 37913 1268 38200
rect 1227 37904 1269 37913
rect 1227 37864 1228 37904
rect 1268 37864 1269 37904
rect 1227 37855 1269 37864
rect 1323 37232 1365 37241
rect 1323 37192 1324 37232
rect 1364 37192 1365 37232
rect 1323 37183 1365 37192
rect 1227 36728 1269 36737
rect 1227 36688 1228 36728
rect 1268 36688 1269 36728
rect 1227 36679 1269 36688
rect 1228 36594 1268 36679
rect 1228 35888 1268 35897
rect 1036 35848 1228 35888
rect 1228 35477 1268 35848
rect 1227 35468 1269 35477
rect 1227 35428 1228 35468
rect 1268 35428 1269 35468
rect 1227 35419 1269 35428
rect 1227 34376 1269 34385
rect 1227 34336 1228 34376
rect 1268 34336 1269 34376
rect 1227 34327 1269 34336
rect 1228 34242 1268 34327
rect 1035 33788 1077 33797
rect 1035 33748 1036 33788
rect 1076 33748 1077 33788
rect 1035 33739 1077 33748
rect 939 15476 981 15485
rect 939 15436 940 15476
rect 980 15436 981 15476
rect 939 15427 981 15436
rect 843 15056 885 15065
rect 843 15016 844 15056
rect 884 15016 885 15056
rect 843 15007 885 15016
rect 1036 13721 1076 33739
rect 1228 33704 1268 33713
rect 1324 33704 1364 37183
rect 1420 34469 1460 42736
rect 1708 37577 1748 46591
rect 1804 41945 1844 65491
rect 1900 61181 1940 73135
rect 1996 62693 2036 74479
rect 2283 70832 2325 70841
rect 2283 70792 2284 70832
rect 2324 70792 2325 70832
rect 2283 70783 2325 70792
rect 2091 67808 2133 67817
rect 2091 67768 2092 67808
rect 2132 67768 2133 67808
rect 2091 67759 2133 67768
rect 1995 62684 2037 62693
rect 1995 62644 1996 62684
rect 2036 62644 2037 62684
rect 1995 62635 2037 62644
rect 1899 61172 1941 61181
rect 1899 61132 1900 61172
rect 1940 61132 1941 61172
rect 1899 61123 1941 61132
rect 1995 60584 2037 60593
rect 1995 60544 1996 60584
rect 2036 60544 2037 60584
rect 1995 60535 2037 60544
rect 1899 57056 1941 57065
rect 1899 57016 1900 57056
rect 1940 57016 1941 57056
rect 1899 57007 1941 57016
rect 1900 46817 1940 57007
rect 1996 51857 2036 60535
rect 2092 58661 2132 67759
rect 2284 66977 2324 70783
rect 2380 70664 2420 81115
rect 2475 72428 2517 72437
rect 2475 72388 2476 72428
rect 2516 72388 2517 72428
rect 2475 72379 2517 72388
rect 2476 72176 2516 72379
rect 2516 72136 2612 72176
rect 2476 72127 2516 72136
rect 2572 71504 2612 72136
rect 2668 72008 2708 72017
rect 2708 71968 2900 72008
rect 2668 71959 2708 71968
rect 2764 71504 2804 71513
rect 2572 71464 2764 71504
rect 2283 66968 2325 66977
rect 2283 66928 2284 66968
rect 2324 66928 2325 66968
rect 2283 66919 2325 66928
rect 2380 66142 2420 70624
rect 2475 70076 2517 70085
rect 2475 70036 2476 70076
rect 2516 70036 2517 70076
rect 2475 70027 2517 70036
rect 2476 69992 2516 70027
rect 2476 68228 2516 69952
rect 2668 69740 2708 69749
rect 2476 68188 2612 68228
rect 2475 67640 2517 67649
rect 2475 67600 2476 67640
rect 2516 67600 2517 67640
rect 2475 67591 2517 67600
rect 2572 67640 2612 68188
rect 2476 66968 2516 67591
rect 2572 67481 2612 67600
rect 2571 67472 2613 67481
rect 2571 67432 2572 67472
rect 2612 67432 2613 67472
rect 2571 67423 2613 67432
rect 2668 67304 2708 69700
rect 2764 68480 2804 71464
rect 2860 69152 2900 71968
rect 2956 71252 2996 71261
rect 2996 71212 3284 71252
rect 2956 71203 2996 71212
rect 2955 70748 2997 70757
rect 2955 70708 2956 70748
rect 2996 70708 2997 70748
rect 2955 70699 2997 70708
rect 2956 69992 2996 70699
rect 2956 69943 2996 69952
rect 2860 69103 2900 69112
rect 2955 69152 2997 69161
rect 2955 69112 2956 69152
rect 2996 69112 2997 69152
rect 2955 69103 2997 69112
rect 2956 69018 2996 69103
rect 3244 68480 3284 71212
rect 3340 69404 3380 83476
rect 3436 83012 3476 83560
rect 3628 83516 3668 83525
rect 3628 83357 3668 83476
rect 4011 83516 4053 83525
rect 4011 83476 4012 83516
rect 4052 83476 4053 83516
rect 4011 83467 4053 83476
rect 4012 83382 4052 83467
rect 3627 83348 3669 83357
rect 3627 83308 3628 83348
rect 3668 83308 3669 83348
rect 3627 83299 3669 83308
rect 3688 83180 4056 83189
rect 3728 83140 3770 83180
rect 3810 83140 3852 83180
rect 3892 83140 3934 83180
rect 3974 83140 4016 83180
rect 3688 83131 4056 83140
rect 3436 82963 3476 82972
rect 3916 83012 3956 83021
rect 4108 83012 4148 83803
rect 4204 83768 4244 84652
rect 4299 84440 4341 84449
rect 4299 84400 4300 84440
rect 4340 84400 4341 84440
rect 4299 84391 4341 84400
rect 4300 84306 4340 84391
rect 4204 83719 4244 83728
rect 4396 83684 4436 84979
rect 4492 84692 4532 85936
rect 4492 84652 4628 84692
rect 4491 84356 4533 84365
rect 4491 84316 4492 84356
rect 4532 84316 4533 84356
rect 4491 84307 4533 84316
rect 4492 84222 4532 84307
rect 4588 83768 4628 84652
rect 4684 83768 4724 85936
rect 4876 84113 4916 85936
rect 5068 84701 5108 85936
rect 5067 84692 5109 84701
rect 5067 84652 5068 84692
rect 5108 84652 5109 84692
rect 5067 84643 5109 84652
rect 5260 84617 5300 85936
rect 5452 84692 5492 85936
rect 5644 85205 5684 85936
rect 5643 85196 5685 85205
rect 5643 85156 5644 85196
rect 5684 85156 5685 85196
rect 5643 85147 5685 85156
rect 5452 84652 5684 84692
rect 5259 84608 5301 84617
rect 5259 84568 5260 84608
rect 5300 84568 5301 84608
rect 5259 84559 5301 84568
rect 4875 84104 4917 84113
rect 4875 84064 4876 84104
rect 4916 84064 4917 84104
rect 4875 84055 4917 84064
rect 5355 84104 5397 84113
rect 5355 84064 5356 84104
rect 5396 84064 5397 84104
rect 5355 84055 5397 84064
rect 4928 83936 5296 83945
rect 4968 83896 5010 83936
rect 5050 83896 5092 83936
rect 5132 83896 5174 83936
rect 5214 83896 5256 83936
rect 4928 83887 5296 83896
rect 4972 83768 5012 83777
rect 4684 83728 4972 83768
rect 4588 83719 4628 83728
rect 4972 83719 5012 83728
rect 5356 83768 5396 84055
rect 5644 83768 5684 84652
rect 5836 84449 5876 85936
rect 6028 85121 6068 85936
rect 6027 85112 6069 85121
rect 6027 85072 6028 85112
rect 6068 85072 6069 85112
rect 6027 85063 6069 85072
rect 6220 84449 6260 85936
rect 6412 85625 6452 85936
rect 6411 85616 6453 85625
rect 6411 85576 6412 85616
rect 6452 85576 6453 85616
rect 6411 85567 6453 85576
rect 6604 84533 6644 85936
rect 6603 84524 6645 84533
rect 6603 84484 6604 84524
rect 6644 84484 6645 84524
rect 6603 84475 6645 84484
rect 6796 84449 6836 85936
rect 5835 84440 5877 84449
rect 5835 84400 5836 84440
rect 5876 84400 5877 84440
rect 5835 84391 5877 84400
rect 6219 84440 6261 84449
rect 6219 84400 6220 84440
rect 6260 84400 6261 84440
rect 6219 84391 6261 84400
rect 6795 84440 6837 84449
rect 6795 84400 6796 84440
rect 6836 84400 6837 84440
rect 6795 84391 6837 84400
rect 6603 83852 6645 83861
rect 6603 83812 6604 83852
rect 6644 83812 6645 83852
rect 6603 83803 6645 83812
rect 5932 83768 5972 83777
rect 5644 83728 5932 83768
rect 5356 83719 5396 83728
rect 5932 83719 5972 83728
rect 5547 83684 5589 83693
rect 4396 83644 4532 83684
rect 4396 83516 4436 83525
rect 4396 83357 4436 83476
rect 4395 83348 4437 83357
rect 4395 83308 4396 83348
rect 4436 83308 4437 83348
rect 4395 83299 4437 83308
rect 3956 82972 4148 83012
rect 4492 83012 4532 83644
rect 5547 83644 5548 83684
rect 5588 83644 5589 83684
rect 5547 83635 5589 83644
rect 4780 83516 4820 83525
rect 4780 83189 4820 83476
rect 5164 83516 5204 83525
rect 5164 83273 5204 83476
rect 5548 83516 5588 83635
rect 5548 83467 5588 83476
rect 6123 83516 6165 83525
rect 6123 83476 6124 83516
rect 6164 83476 6165 83516
rect 6123 83467 6165 83476
rect 6508 83516 6548 83525
rect 6124 83382 6164 83467
rect 5163 83264 5205 83273
rect 5163 83224 5164 83264
rect 5204 83224 5205 83264
rect 5163 83215 5205 83224
rect 6508 83189 6548 83476
rect 4779 83180 4821 83189
rect 4779 83140 4780 83180
rect 4820 83140 4821 83180
rect 4779 83131 4821 83140
rect 5547 83180 5589 83189
rect 5547 83140 5548 83180
rect 5588 83140 5589 83180
rect 5547 83131 5589 83140
rect 6507 83180 6549 83189
rect 6507 83140 6508 83180
rect 6548 83140 6549 83180
rect 6507 83131 6549 83140
rect 4588 83012 4628 83021
rect 4492 82972 4588 83012
rect 3916 82963 3956 82972
rect 4588 82963 4628 82972
rect 3627 82844 3669 82853
rect 3627 82804 3628 82844
rect 3668 82804 3669 82844
rect 3627 82795 3669 82804
rect 4107 82844 4149 82853
rect 4107 82804 4108 82844
rect 4148 82804 4149 82844
rect 4107 82795 4149 82804
rect 4779 82844 4821 82853
rect 4779 82804 4780 82844
rect 4820 82804 4821 82844
rect 4779 82795 4821 82804
rect 3628 82710 3668 82795
rect 4108 82710 4148 82795
rect 4780 82710 4820 82795
rect 4928 82424 5296 82433
rect 4968 82384 5010 82424
rect 5050 82384 5092 82424
rect 5132 82384 5174 82424
rect 5214 82384 5256 82424
rect 4928 82375 5296 82384
rect 3688 81668 4056 81677
rect 3728 81628 3770 81668
rect 3810 81628 3852 81668
rect 3892 81628 3934 81668
rect 3974 81628 4016 81668
rect 3688 81619 4056 81628
rect 5451 81248 5493 81257
rect 5451 81208 5452 81248
rect 5492 81208 5493 81248
rect 5451 81199 5493 81208
rect 4928 80912 5296 80921
rect 4968 80872 5010 80912
rect 5050 80872 5092 80912
rect 5132 80872 5174 80912
rect 5214 80872 5256 80912
rect 4928 80863 5296 80872
rect 3688 80156 4056 80165
rect 3728 80116 3770 80156
rect 3810 80116 3852 80156
rect 3892 80116 3934 80156
rect 3974 80116 4016 80156
rect 3688 80107 4056 80116
rect 3531 79484 3573 79493
rect 3531 79444 3532 79484
rect 3572 79444 3573 79484
rect 3531 79435 3573 79444
rect 3532 73688 3572 79435
rect 4928 79400 5296 79409
rect 4968 79360 5010 79400
rect 5050 79360 5092 79400
rect 5132 79360 5174 79400
rect 5214 79360 5256 79400
rect 4928 79351 5296 79360
rect 5355 78812 5397 78821
rect 5355 78772 5356 78812
rect 5396 78772 5397 78812
rect 5355 78763 5397 78772
rect 3688 78644 4056 78653
rect 3728 78604 3770 78644
rect 3810 78604 3852 78644
rect 3892 78604 3934 78644
rect 3974 78604 4016 78644
rect 3688 78595 4056 78604
rect 4928 77888 5296 77897
rect 4968 77848 5010 77888
rect 5050 77848 5092 77888
rect 5132 77848 5174 77888
rect 5214 77848 5256 77888
rect 4928 77839 5296 77848
rect 3688 77132 4056 77141
rect 3728 77092 3770 77132
rect 3810 77092 3852 77132
rect 3892 77092 3934 77132
rect 3974 77092 4016 77132
rect 3688 77083 4056 77092
rect 4299 76796 4341 76805
rect 4299 76756 4300 76796
rect 4340 76756 4341 76796
rect 4299 76747 4341 76756
rect 3688 75620 4056 75629
rect 3728 75580 3770 75620
rect 3810 75580 3852 75620
rect 3892 75580 3934 75620
rect 3974 75580 4016 75620
rect 3688 75571 4056 75580
rect 3688 74108 4056 74117
rect 3728 74068 3770 74108
rect 3810 74068 3852 74108
rect 3892 74068 3934 74108
rect 3974 74068 4016 74108
rect 3688 74059 4056 74068
rect 3724 73688 3764 73697
rect 3532 73648 3724 73688
rect 3435 72428 3477 72437
rect 3435 72388 3436 72428
rect 3476 72388 3477 72428
rect 3435 72379 3477 72388
rect 3436 70496 3476 72379
rect 3532 70673 3572 73648
rect 3724 73639 3764 73648
rect 3916 73016 3956 73025
rect 3916 72773 3956 72976
rect 3915 72764 3957 72773
rect 3915 72724 3916 72764
rect 3956 72724 3957 72764
rect 3915 72715 3957 72724
rect 4107 72764 4149 72773
rect 4107 72724 4108 72764
rect 4148 72724 4149 72764
rect 4107 72715 4149 72724
rect 3688 72596 4056 72605
rect 3728 72556 3770 72596
rect 3810 72556 3852 72596
rect 3892 72556 3934 72596
rect 3974 72556 4016 72596
rect 3688 72547 4056 72556
rect 3688 71084 4056 71093
rect 3728 71044 3770 71084
rect 3810 71044 3852 71084
rect 3892 71044 3934 71084
rect 3974 71044 4016 71084
rect 3688 71035 4056 71044
rect 4011 70748 4053 70757
rect 4011 70708 4012 70748
rect 4052 70708 4053 70748
rect 4011 70699 4053 70708
rect 3531 70664 3573 70673
rect 3531 70624 3532 70664
rect 3572 70624 3573 70664
rect 3531 70615 3573 70624
rect 3628 70664 3668 70673
rect 3628 70496 3668 70624
rect 4012 70664 4052 70699
rect 4012 70613 4052 70624
rect 3820 70505 3860 70590
rect 3436 70456 3668 70496
rect 3628 70337 3668 70456
rect 3819 70496 3861 70505
rect 3819 70456 3820 70496
rect 3860 70456 3861 70496
rect 3819 70447 3861 70456
rect 3627 70328 3669 70337
rect 3627 70288 3628 70328
rect 3668 70288 3669 70328
rect 3627 70279 3669 70288
rect 3688 69572 4056 69581
rect 3728 69532 3770 69572
rect 3810 69532 3852 69572
rect 3892 69532 3934 69572
rect 3974 69532 4016 69572
rect 3688 69523 4056 69532
rect 3340 69364 3668 69404
rect 3340 69152 3380 69161
rect 3340 68741 3380 69112
rect 3436 69152 3476 69163
rect 3436 69077 3476 69112
rect 3531 69152 3573 69161
rect 3531 69112 3532 69152
rect 3572 69112 3573 69152
rect 3531 69103 3573 69112
rect 3435 69068 3477 69077
rect 3435 69028 3436 69068
rect 3476 69028 3477 69068
rect 3435 69019 3477 69028
rect 3339 68732 3381 68741
rect 3339 68692 3340 68732
rect 3380 68692 3381 68732
rect 3339 68683 3381 68692
rect 3436 68480 3476 68489
rect 3244 68440 3436 68480
rect 2764 67649 2804 68440
rect 3436 68431 3476 68440
rect 3532 68480 3572 69103
rect 2956 68228 2996 68237
rect 2956 67817 2996 68188
rect 3532 67976 3572 68440
rect 3628 68237 3668 69364
rect 3915 69152 3957 69161
rect 3915 69112 3916 69152
rect 3956 69112 3957 69152
rect 3915 69103 3957 69112
rect 3916 69018 3956 69103
rect 4011 69068 4053 69077
rect 4011 69028 4012 69068
rect 4052 69028 4053 69068
rect 4011 69019 4053 69028
rect 3915 68732 3957 68741
rect 3915 68692 3916 68732
rect 3956 68692 3957 68732
rect 3915 68683 3957 68692
rect 3916 68405 3956 68683
rect 4012 68480 4052 69019
rect 4108 68564 4148 72715
rect 4300 72176 4340 76747
rect 4928 76376 5296 76385
rect 4968 76336 5010 76376
rect 5050 76336 5092 76376
rect 5132 76336 5174 76376
rect 5214 76336 5256 76376
rect 4928 76327 5296 76336
rect 4928 74864 5296 74873
rect 4968 74824 5010 74864
rect 5050 74824 5092 74864
rect 5132 74824 5174 74864
rect 5214 74824 5256 74864
rect 4928 74815 5296 74824
rect 5356 74705 5396 78763
rect 5355 74696 5397 74705
rect 5164 74656 5356 74696
rect 5396 74656 5397 74696
rect 4971 74528 5013 74537
rect 4971 74488 4972 74528
rect 5012 74488 5013 74528
rect 4971 74479 5013 74488
rect 5164 74528 5204 74656
rect 5355 74647 5397 74656
rect 5356 74562 5396 74647
rect 5164 74479 5204 74488
rect 4972 73688 5012 74479
rect 5452 73865 5492 81199
rect 5451 73856 5493 73865
rect 5451 73816 5452 73856
rect 5492 73816 5493 73856
rect 5451 73807 5493 73816
rect 4972 73604 5012 73648
rect 5452 73688 5492 73699
rect 5452 73613 5492 73648
rect 5548 73688 5588 83131
rect 6315 82004 6357 82013
rect 6315 81964 6316 82004
rect 6356 81964 6357 82004
rect 6315 81955 6357 81964
rect 6123 79148 6165 79157
rect 6123 79108 6124 79148
rect 6164 79108 6165 79148
rect 6123 79099 6165 79108
rect 5643 74696 5685 74705
rect 5643 74656 5644 74696
rect 5684 74656 5685 74696
rect 5643 74647 5685 74656
rect 4780 73564 5012 73604
rect 5163 73604 5205 73613
rect 5163 73564 5164 73604
rect 5204 73564 5205 73604
rect 4780 73100 4820 73564
rect 5163 73555 5205 73564
rect 5451 73604 5493 73613
rect 5451 73564 5452 73604
rect 5492 73564 5493 73604
rect 5451 73555 5493 73564
rect 5164 73470 5204 73555
rect 4928 73352 5296 73361
rect 4968 73312 5010 73352
rect 5050 73312 5092 73352
rect 5132 73312 5174 73352
rect 5214 73312 5256 73352
rect 4928 73303 5296 73312
rect 5548 73100 5588 73648
rect 4492 73060 4820 73100
rect 5452 73060 5588 73100
rect 4340 72136 4436 72176
rect 4300 72127 4340 72136
rect 4299 70496 4341 70505
rect 4299 70456 4300 70496
rect 4340 70456 4341 70496
rect 4299 70447 4341 70456
rect 4203 70328 4245 70337
rect 4203 70288 4204 70328
rect 4244 70288 4245 70328
rect 4203 70279 4245 70288
rect 4204 69992 4244 70279
rect 4204 69943 4244 69952
rect 4300 69572 4340 70447
rect 4396 70421 4436 72136
rect 4395 70412 4437 70421
rect 4395 70372 4396 70412
rect 4436 70372 4437 70412
rect 4395 70363 4437 70372
rect 4396 70169 4436 70363
rect 4492 70253 4532 73060
rect 5164 73016 5204 73025
rect 5164 72017 5204 72976
rect 5356 72764 5396 72773
rect 5163 72008 5205 72017
rect 5163 71968 5164 72008
rect 5204 71968 5205 72008
rect 5163 71959 5205 71968
rect 4928 71840 5296 71849
rect 4968 71800 5010 71840
rect 5050 71800 5092 71840
rect 5132 71800 5174 71840
rect 5214 71800 5256 71840
rect 4928 71791 5296 71800
rect 5067 71588 5109 71597
rect 5067 71548 5068 71588
rect 5108 71548 5109 71588
rect 5067 71539 5109 71548
rect 4587 71504 4629 71513
rect 4587 71464 4588 71504
rect 4628 71464 4629 71504
rect 4587 71455 4629 71464
rect 4684 71504 4724 71513
rect 4588 71370 4628 71455
rect 4587 70412 4629 70421
rect 4587 70372 4588 70412
rect 4628 70372 4629 70412
rect 4587 70363 4629 70372
rect 4491 70244 4533 70253
rect 4491 70204 4492 70244
rect 4532 70204 4533 70244
rect 4491 70195 4533 70204
rect 4395 70160 4437 70169
rect 4395 70120 4396 70160
rect 4436 70120 4437 70160
rect 4395 70111 4437 70120
rect 4588 70034 4628 70363
rect 4491 69992 4533 70001
rect 4588 69992 4628 69994
rect 4491 69952 4492 69992
rect 4532 69952 4628 69992
rect 4491 69943 4533 69952
rect 4396 69740 4436 69749
rect 4436 69700 4628 69740
rect 4396 69691 4436 69700
rect 4300 69532 4436 69572
rect 4396 69166 4436 69532
rect 4396 69117 4436 69126
rect 4491 69152 4533 69161
rect 4491 69112 4492 69152
rect 4532 69112 4533 69152
rect 4588 69152 4628 69700
rect 4684 69329 4724 71464
rect 5068 71504 5108 71539
rect 5356 71513 5396 72724
rect 5068 70505 5108 71464
rect 5355 71504 5397 71513
rect 5355 71464 5356 71504
rect 5396 71464 5397 71504
rect 5355 71455 5397 71464
rect 5164 71420 5204 71429
rect 5164 71261 5204 71380
rect 5259 71420 5301 71429
rect 5259 71380 5260 71420
rect 5300 71380 5301 71420
rect 5259 71371 5301 71380
rect 5163 71252 5205 71261
rect 5163 71212 5164 71252
rect 5204 71212 5205 71252
rect 5163 71203 5205 71212
rect 5260 70664 5300 71371
rect 5452 71168 5492 73060
rect 5547 72176 5589 72185
rect 5547 72136 5548 72176
rect 5588 72136 5589 72176
rect 5547 72127 5589 72136
rect 5548 72042 5588 72127
rect 5644 71672 5684 74647
rect 5931 73856 5973 73865
rect 5931 73816 5932 73856
rect 5972 73816 5973 73856
rect 5931 73807 5973 73816
rect 5932 73772 5972 73807
rect 5932 73721 5972 73732
rect 6027 73688 6069 73697
rect 6027 73648 6028 73688
rect 6068 73648 6069 73688
rect 6027 73639 6069 73648
rect 6028 73554 6068 73639
rect 5932 72176 5972 72185
rect 6124 72176 6164 79099
rect 6316 73100 6356 81955
rect 6604 81920 6644 83803
rect 6699 83768 6741 83777
rect 6699 83728 6700 83768
rect 6740 83728 6741 83768
rect 6699 83719 6741 83728
rect 6700 83634 6740 83719
rect 6988 83684 7028 85936
rect 7180 85877 7220 85936
rect 7179 85868 7221 85877
rect 7179 85828 7180 85868
rect 7220 85828 7221 85868
rect 7179 85819 7221 85828
rect 7372 84692 7412 85936
rect 7564 84776 7604 85936
rect 7756 84869 7796 85936
rect 7755 84860 7797 84869
rect 7755 84820 7756 84860
rect 7796 84820 7797 84860
rect 7755 84811 7797 84820
rect 7180 84652 7412 84692
rect 7468 84736 7604 84776
rect 7180 83768 7220 84652
rect 7468 83777 7508 84736
rect 7755 84524 7797 84533
rect 7755 84484 7756 84524
rect 7796 84484 7797 84524
rect 7755 84475 7797 84484
rect 7563 84020 7605 84029
rect 7563 83980 7564 84020
rect 7604 83980 7605 84020
rect 7563 83971 7605 83980
rect 7180 83719 7220 83728
rect 7467 83768 7509 83777
rect 7467 83728 7468 83768
rect 7508 83728 7509 83768
rect 7467 83719 7509 83728
rect 7564 83768 7604 83971
rect 7564 83719 7604 83728
rect 7756 83768 7796 84475
rect 7851 83936 7893 83945
rect 7851 83896 7852 83936
rect 7892 83896 7893 83936
rect 7851 83887 7893 83896
rect 7756 83719 7796 83728
rect 6988 83644 7124 83684
rect 6987 83516 7029 83525
rect 6987 83476 6988 83516
rect 7028 83476 7029 83516
rect 6987 83467 7029 83476
rect 6988 83382 7028 83467
rect 6508 81880 6644 81920
rect 6411 74528 6453 74537
rect 6411 74488 6412 74528
rect 6452 74488 6453 74528
rect 6411 74479 6453 74488
rect 6412 74394 6452 74479
rect 6508 73688 6548 81880
rect 6700 76712 6740 76721
rect 6700 76385 6740 76672
rect 6699 76376 6741 76385
rect 6699 76336 6700 76376
rect 6740 76336 6741 76376
rect 6699 76327 6741 76336
rect 6700 76040 6740 76049
rect 6740 76000 6932 76040
rect 6700 75991 6740 76000
rect 6795 75452 6837 75461
rect 6795 75412 6796 75452
rect 6836 75412 6837 75452
rect 6795 75403 6837 75412
rect 6700 75200 6740 75209
rect 6700 74705 6740 75160
rect 6699 74696 6741 74705
rect 6699 74656 6700 74696
rect 6740 74656 6741 74696
rect 6699 74647 6741 74656
rect 6796 74528 6836 75403
rect 6796 74479 6836 74488
rect 6603 74276 6645 74285
rect 6603 74236 6604 74276
rect 6644 74236 6645 74276
rect 6603 74227 6645 74236
rect 6604 74142 6644 74227
rect 6508 73639 6548 73648
rect 6316 73060 6548 73100
rect 5972 72136 6164 72176
rect 5932 72127 5972 72136
rect 5260 70589 5300 70624
rect 5356 71128 5492 71168
rect 5548 71632 5684 71672
rect 5740 72008 5780 72017
rect 5259 70580 5301 70589
rect 5259 70540 5260 70580
rect 5300 70540 5301 70580
rect 5259 70531 5301 70540
rect 5067 70496 5109 70505
rect 5260 70500 5300 70531
rect 5067 70456 5068 70496
rect 5108 70456 5109 70496
rect 5067 70447 5109 70456
rect 4928 70328 5296 70337
rect 4968 70288 5010 70328
rect 5050 70288 5092 70328
rect 5132 70288 5174 70328
rect 5214 70288 5256 70328
rect 4928 70279 5296 70288
rect 4971 70160 5013 70169
rect 4971 70120 4972 70160
rect 5012 70120 5013 70160
rect 4971 70111 5013 70120
rect 4683 69320 4725 69329
rect 4683 69280 4684 69320
rect 4724 69280 4725 69320
rect 4683 69271 4725 69280
rect 4972 69161 5012 70111
rect 4779 69152 4821 69161
rect 4588 69112 4724 69152
rect 4491 69103 4533 69112
rect 4108 68524 4340 68564
rect 4052 68440 4148 68480
rect 4012 68431 4052 68440
rect 3915 68396 3957 68405
rect 3915 68356 3916 68396
rect 3956 68356 3957 68396
rect 3915 68347 3957 68356
rect 3916 68262 3956 68347
rect 3627 68228 3669 68237
rect 3627 68188 3628 68228
rect 3668 68188 3669 68228
rect 3627 68179 3669 68188
rect 3688 68060 4056 68069
rect 3728 68020 3770 68060
rect 3810 68020 3852 68060
rect 3892 68020 3934 68060
rect 3974 68020 4016 68060
rect 3688 68011 4056 68020
rect 3436 67936 3572 67976
rect 2955 67808 2997 67817
rect 2955 67768 2956 67808
rect 2996 67768 2997 67808
rect 2955 67759 2997 67768
rect 2763 67640 2805 67649
rect 2763 67600 2764 67640
rect 2804 67600 2805 67640
rect 2763 67591 2805 67600
rect 2956 67640 2996 67651
rect 2956 67565 2996 67600
rect 2955 67556 2997 67565
rect 2955 67516 2956 67556
rect 2996 67516 2997 67556
rect 2955 67507 2997 67516
rect 2764 67472 2804 67481
rect 3051 67472 3093 67481
rect 2804 67432 2900 67472
rect 2764 67423 2804 67432
rect 2668 67264 2804 67304
rect 2516 66928 2612 66968
rect 2476 66919 2516 66928
rect 2187 66128 2229 66137
rect 2187 66088 2188 66128
rect 2228 66088 2229 66128
rect 2187 66079 2229 66088
rect 2284 66102 2420 66142
rect 2572 66128 2612 66928
rect 2668 66725 2708 66810
rect 2667 66716 2709 66725
rect 2667 66676 2668 66716
rect 2708 66676 2709 66716
rect 2667 66667 2709 66676
rect 2668 66128 2708 66137
rect 2091 58652 2133 58661
rect 2091 58612 2092 58652
rect 2132 58612 2133 58652
rect 2091 58603 2133 58612
rect 2188 56057 2228 66079
rect 2284 60845 2324 66102
rect 2572 66088 2668 66128
rect 2668 64793 2708 66088
rect 2764 65456 2804 67264
rect 2860 66137 2900 67432
rect 3051 67432 3052 67472
rect 3092 67432 3093 67472
rect 3051 67423 3093 67432
rect 2955 66716 2997 66725
rect 2955 66676 2956 66716
rect 2996 66676 2997 66716
rect 2955 66667 2997 66676
rect 2859 66128 2901 66137
rect 2859 66088 2860 66128
rect 2900 66088 2901 66128
rect 2859 66079 2901 66088
rect 2860 65960 2900 65969
rect 2860 65633 2900 65920
rect 2859 65624 2901 65633
rect 2859 65584 2860 65624
rect 2900 65584 2901 65624
rect 2859 65575 2901 65584
rect 2764 65407 2804 65416
rect 2859 65456 2901 65465
rect 2859 65416 2860 65456
rect 2900 65416 2901 65456
rect 2859 65407 2901 65416
rect 2860 65322 2900 65407
rect 2667 64784 2709 64793
rect 2667 64744 2668 64784
rect 2708 64744 2709 64784
rect 2667 64735 2709 64744
rect 2571 64616 2613 64625
rect 2571 64576 2572 64616
rect 2612 64576 2613 64616
rect 2571 64567 2613 64576
rect 2572 64482 2612 64567
rect 2956 64280 2996 66667
rect 2860 64240 2996 64280
rect 2763 64112 2805 64121
rect 2763 64072 2764 64112
rect 2804 64072 2805 64112
rect 2763 64063 2805 64072
rect 2571 62768 2613 62777
rect 2571 62728 2572 62768
rect 2612 62728 2613 62768
rect 2571 62719 2613 62728
rect 2476 62432 2516 62441
rect 2572 62432 2612 62719
rect 2516 62392 2612 62432
rect 2476 62383 2516 62392
rect 2475 62264 2517 62273
rect 2475 62224 2476 62264
rect 2516 62224 2517 62264
rect 2475 62215 2517 62224
rect 2283 60836 2325 60845
rect 2283 60796 2284 60836
rect 2324 60796 2325 60836
rect 2283 60787 2325 60796
rect 2476 60080 2516 62215
rect 2572 60929 2612 62392
rect 2764 62264 2804 64063
rect 2860 63104 2900 64240
rect 2955 63944 2997 63953
rect 2955 63904 2956 63944
rect 2996 63904 2997 63944
rect 2955 63895 2997 63904
rect 2956 63810 2996 63895
rect 2860 63055 2900 63064
rect 2955 63104 2997 63113
rect 2955 63064 2956 63104
rect 2996 63064 2997 63104
rect 2955 63055 2997 63064
rect 2956 62970 2996 63055
rect 3052 62777 3092 67423
rect 3340 66968 3380 66977
rect 3244 66928 3340 66968
rect 3244 66305 3284 66928
rect 3340 66919 3380 66928
rect 3436 66389 3476 67936
rect 3531 67808 3573 67817
rect 3531 67768 3532 67808
rect 3572 67768 3573 67808
rect 3531 67759 3573 67768
rect 3435 66380 3477 66389
rect 3435 66340 3436 66380
rect 3476 66340 3477 66380
rect 3435 66331 3477 66340
rect 3243 66296 3285 66305
rect 3243 66256 3244 66296
rect 3284 66256 3285 66296
rect 3243 66247 3285 66256
rect 3532 66128 3572 67759
rect 4108 67472 4148 68440
rect 4204 67649 4244 67734
rect 4203 67640 4245 67649
rect 4203 67600 4204 67640
rect 4244 67600 4245 67640
rect 4203 67591 4245 67600
rect 4108 67432 4244 67472
rect 3688 66548 4056 66557
rect 3728 66508 3770 66548
rect 3810 66508 3852 66548
rect 3892 66508 3934 66548
rect 3974 66508 4016 66548
rect 3688 66499 4056 66508
rect 3723 66380 3765 66389
rect 3723 66340 3724 66380
rect 3764 66340 3765 66380
rect 3723 66331 3765 66340
rect 3628 66128 3668 66137
rect 3532 66088 3628 66128
rect 3628 66079 3668 66088
rect 3724 66128 3764 66331
rect 4204 66212 4244 67432
rect 4300 67061 4340 68524
rect 4492 68480 4532 69103
rect 4587 68984 4629 68993
rect 4587 68944 4588 68984
rect 4628 68944 4629 68984
rect 4587 68935 4629 68944
rect 4588 68850 4628 68935
rect 4684 68648 4724 69112
rect 4779 69112 4780 69152
rect 4820 69112 4821 69152
rect 4779 69103 4821 69112
rect 4971 69152 5013 69161
rect 4971 69112 4972 69152
rect 5012 69112 5013 69152
rect 4971 69103 5013 69112
rect 4780 69018 4820 69103
rect 4928 68816 5296 68825
rect 4968 68776 5010 68816
rect 5050 68776 5092 68816
rect 5132 68776 5174 68816
rect 5214 68776 5256 68816
rect 4928 68767 5296 68776
rect 5356 68741 5396 71128
rect 5451 71000 5493 71009
rect 5451 70960 5452 71000
rect 5492 70960 5493 71000
rect 5451 70951 5493 70960
rect 5452 70916 5492 70951
rect 5452 70865 5492 70876
rect 5451 70748 5493 70757
rect 5451 70708 5452 70748
rect 5492 70708 5493 70748
rect 5451 70699 5493 70708
rect 5355 68732 5397 68741
rect 5355 68692 5356 68732
rect 5396 68692 5397 68732
rect 5355 68683 5397 68692
rect 4684 68608 5012 68648
rect 4532 68440 4724 68480
rect 4492 68431 4532 68440
rect 4588 67640 4628 67649
rect 4492 67600 4588 67640
rect 4396 67472 4436 67481
rect 4299 67052 4341 67061
rect 4299 67012 4300 67052
rect 4340 67012 4341 67052
rect 4299 67003 4341 67012
rect 4396 66221 4436 67432
rect 3243 66044 3285 66053
rect 3243 66004 3244 66044
rect 3284 66004 3285 66044
rect 3243 65995 3285 66004
rect 3147 65540 3189 65549
rect 3147 65500 3148 65540
rect 3188 65500 3189 65540
rect 3147 65491 3189 65500
rect 3148 65129 3188 65491
rect 3244 65456 3284 65995
rect 3627 65624 3669 65633
rect 3627 65584 3628 65624
rect 3668 65584 3669 65624
rect 3627 65575 3669 65584
rect 3628 65456 3668 65575
rect 3724 65465 3764 66088
rect 4108 66128 4148 66139
rect 4108 66053 4148 66088
rect 4107 66044 4149 66053
rect 4107 66004 4108 66044
rect 4148 66004 4149 66044
rect 4107 65995 4149 66004
rect 3915 65708 3957 65717
rect 3915 65668 3916 65708
rect 3956 65668 3957 65708
rect 3915 65659 3957 65668
rect 3819 65540 3861 65549
rect 3819 65500 3820 65540
rect 3860 65500 3861 65540
rect 3819 65491 3861 65500
rect 3244 65407 3284 65416
rect 3340 65416 3668 65456
rect 3723 65456 3765 65465
rect 3723 65416 3724 65456
rect 3764 65416 3765 65456
rect 3340 65414 3380 65416
rect 3723 65407 3765 65416
rect 3820 65456 3860 65491
rect 3820 65405 3860 65416
rect 3147 65120 3189 65129
rect 3147 65080 3148 65120
rect 3188 65080 3189 65120
rect 3147 65071 3189 65080
rect 3147 64784 3189 64793
rect 3147 64744 3148 64784
rect 3188 64744 3189 64784
rect 3147 64735 3189 64744
rect 3148 63953 3188 64735
rect 3243 64280 3285 64289
rect 3243 64240 3244 64280
rect 3284 64240 3285 64280
rect 3243 64231 3285 64240
rect 3147 63944 3189 63953
rect 3147 63904 3148 63944
rect 3188 63904 3189 63944
rect 3147 63895 3189 63904
rect 3147 63692 3189 63701
rect 3147 63652 3148 63692
rect 3188 63652 3189 63692
rect 3147 63643 3189 63652
rect 3148 63558 3188 63643
rect 3147 63440 3189 63449
rect 3147 63400 3148 63440
rect 3188 63400 3189 63440
rect 3147 63391 3189 63400
rect 3148 63113 3188 63391
rect 3147 63104 3189 63113
rect 3147 63064 3148 63104
rect 3188 63064 3189 63104
rect 3147 63055 3189 63064
rect 3051 62768 3093 62777
rect 3051 62728 3052 62768
rect 3092 62728 3093 62768
rect 3051 62719 3093 62728
rect 2956 62441 2996 62526
rect 2955 62432 2997 62441
rect 2955 62392 2956 62432
rect 2996 62392 2997 62432
rect 2955 62383 2997 62392
rect 2764 62224 3092 62264
rect 2668 62180 2708 62189
rect 2668 61601 2708 62140
rect 2763 61760 2805 61769
rect 2763 61720 2764 61760
rect 2804 61720 2805 61760
rect 2763 61711 2805 61720
rect 2667 61592 2709 61601
rect 2667 61552 2668 61592
rect 2708 61552 2709 61592
rect 2667 61543 2709 61552
rect 2571 60920 2613 60929
rect 2668 60920 2708 60929
rect 2571 60880 2572 60920
rect 2612 60880 2668 60920
rect 2571 60871 2613 60880
rect 2668 60871 2708 60880
rect 2572 60786 2612 60871
rect 2667 60752 2709 60761
rect 2667 60712 2668 60752
rect 2708 60712 2709 60752
rect 2667 60703 2709 60712
rect 2668 60332 2708 60703
rect 2668 60283 2708 60292
rect 2283 59408 2325 59417
rect 2283 59368 2284 59408
rect 2324 59368 2325 59408
rect 2283 59359 2325 59368
rect 2187 56048 2229 56057
rect 2187 56008 2188 56048
rect 2228 56008 2229 56048
rect 2187 55999 2229 56008
rect 2284 53957 2324 59359
rect 2283 53948 2325 53957
rect 2283 53908 2284 53948
rect 2324 53908 2325 53948
rect 2283 53899 2325 53908
rect 2284 53612 2324 53899
rect 2092 53572 2324 53612
rect 1995 51848 2037 51857
rect 1995 51808 1996 51848
rect 2036 51808 2037 51848
rect 1995 51799 2037 51808
rect 2092 50933 2132 53572
rect 2187 53360 2229 53369
rect 2187 53320 2188 53360
rect 2228 53320 2229 53360
rect 2187 53311 2229 53320
rect 2476 53360 2516 60040
rect 2764 59417 2804 61711
rect 2859 61592 2901 61601
rect 2859 61552 2860 61592
rect 2900 61552 2901 61592
rect 2859 61543 2901 61552
rect 2956 61592 2996 61601
rect 2860 61458 2900 61543
rect 2956 61256 2996 61552
rect 3052 61433 3092 62224
rect 3051 61424 3093 61433
rect 3051 61384 3052 61424
rect 3092 61384 3093 61424
rect 3051 61375 3093 61384
rect 3148 61256 3188 63055
rect 2956 61216 3188 61256
rect 2859 61088 2901 61097
rect 2859 61048 2860 61088
rect 2900 61048 2901 61088
rect 2859 61039 2901 61048
rect 2860 60954 2900 61039
rect 2956 60668 2996 61216
rect 3244 61088 3284 64231
rect 3340 63281 3380 65374
rect 3916 65288 3956 65659
rect 4204 65633 4244 66172
rect 4395 66212 4437 66221
rect 4395 66172 4396 66212
rect 4436 66172 4437 66212
rect 4395 66163 4437 66172
rect 4299 66128 4341 66137
rect 4299 66088 4300 66128
rect 4340 66088 4341 66128
rect 4299 66079 4341 66088
rect 4203 65624 4245 65633
rect 4203 65584 4204 65624
rect 4244 65584 4245 65624
rect 4203 65575 4245 65584
rect 4300 65451 4340 66079
rect 4492 66044 4532 67600
rect 4588 67591 4628 67600
rect 4587 66968 4629 66977
rect 4587 66928 4588 66968
rect 4628 66928 4629 66968
rect 4587 66919 4629 66928
rect 4588 66834 4628 66919
rect 4587 66128 4629 66137
rect 4587 66088 4588 66128
rect 4628 66088 4629 66128
rect 4587 66079 4629 66088
rect 4684 66128 4724 68440
rect 4972 68475 5012 68608
rect 5164 68564 5204 68573
rect 5204 68524 5396 68564
rect 5164 68515 5204 68524
rect 4972 68426 5012 68435
rect 4928 67304 5296 67313
rect 4968 67264 5010 67304
rect 5050 67264 5092 67304
rect 5132 67264 5174 67304
rect 5214 67264 5256 67304
rect 4928 67255 5296 67264
rect 4971 67052 5013 67061
rect 4971 67012 4972 67052
rect 5012 67012 5013 67052
rect 4971 67003 5013 67012
rect 4972 66968 5012 67003
rect 4972 66917 5012 66928
rect 5356 66893 5396 68524
rect 5355 66884 5397 66893
rect 5355 66844 5356 66884
rect 5396 66844 5397 66884
rect 5355 66835 5397 66844
rect 4779 66800 4821 66809
rect 4779 66760 4780 66800
rect 4820 66760 4821 66800
rect 4779 66751 4821 66760
rect 4780 66666 4820 66751
rect 5163 66212 5205 66221
rect 5163 66172 5164 66212
rect 5204 66172 5205 66212
rect 5163 66163 5205 66172
rect 4396 66004 4532 66044
rect 4396 65465 4436 66004
rect 4492 65540 4532 65549
rect 4300 65402 4340 65411
rect 4395 65456 4437 65465
rect 4395 65416 4396 65456
rect 4436 65416 4437 65456
rect 4395 65407 4437 65416
rect 3532 65248 3956 65288
rect 4299 65288 4341 65297
rect 4299 65248 4300 65288
rect 4340 65248 4341 65288
rect 3435 65120 3477 65129
rect 3435 65080 3436 65120
rect 3476 65080 3477 65120
rect 3435 65071 3477 65080
rect 3436 63944 3476 65071
rect 3532 64121 3572 65248
rect 4299 65239 4341 65248
rect 3688 65036 4056 65045
rect 3728 64996 3770 65036
rect 3810 64996 3852 65036
rect 3892 64996 3934 65036
rect 3974 64996 4016 65036
rect 3688 64987 4056 64996
rect 3819 64784 3861 64793
rect 3819 64744 3820 64784
rect 3860 64744 3861 64784
rect 3819 64735 3861 64744
rect 3820 64616 3860 64735
rect 3820 64567 3860 64576
rect 4204 64616 4244 64644
rect 4300 64616 4340 65239
rect 4396 64625 4436 65407
rect 4492 65297 4532 65500
rect 4491 65288 4533 65297
rect 4491 65248 4492 65288
rect 4532 65248 4533 65288
rect 4491 65239 4533 65248
rect 4244 64576 4340 64616
rect 4204 64567 4244 64576
rect 4012 64448 4052 64457
rect 4052 64408 4148 64448
rect 4012 64399 4052 64408
rect 4011 64196 4053 64205
rect 4011 64156 4012 64196
rect 4052 64156 4053 64196
rect 4011 64147 4053 64156
rect 3531 64112 3573 64121
rect 3531 64072 3532 64112
rect 3572 64072 3573 64112
rect 3531 64063 3573 64072
rect 3436 63895 3476 63904
rect 3532 63944 3572 63953
rect 3435 63776 3477 63785
rect 3435 63736 3436 63776
rect 3476 63736 3477 63776
rect 3435 63727 3477 63736
rect 3339 63272 3381 63281
rect 3339 63232 3340 63272
rect 3380 63232 3381 63272
rect 3339 63223 3381 63232
rect 3436 63188 3476 63727
rect 3532 63449 3572 63904
rect 4012 63944 4052 64147
rect 4108 64121 4148 64408
rect 4107 64112 4149 64121
rect 4107 64072 4108 64112
rect 4148 64072 4149 64112
rect 4107 64063 4149 64072
rect 3916 63860 3956 63871
rect 4012 63869 4052 63904
rect 3916 63785 3956 63820
rect 4011 63860 4053 63869
rect 4011 63820 4012 63860
rect 4052 63820 4053 63860
rect 4011 63811 4053 63820
rect 3915 63776 3957 63785
rect 4012 63780 4052 63811
rect 3915 63736 3916 63776
rect 3956 63736 3957 63776
rect 3915 63727 3957 63736
rect 4203 63776 4245 63785
rect 4203 63736 4204 63776
rect 4244 63736 4245 63776
rect 4203 63727 4245 63736
rect 3688 63524 4056 63533
rect 3728 63484 3770 63524
rect 3810 63484 3852 63524
rect 3892 63484 3934 63524
rect 3974 63484 4016 63524
rect 3688 63475 4056 63484
rect 3531 63440 3573 63449
rect 3531 63400 3532 63440
rect 3572 63400 3573 63440
rect 3531 63391 3573 63400
rect 3915 63356 3957 63365
rect 3915 63316 3916 63356
rect 3956 63316 3957 63356
rect 3915 63307 3957 63316
rect 3531 63272 3573 63281
rect 3531 63232 3532 63272
rect 3572 63232 3573 63272
rect 3531 63223 3573 63232
rect 3339 63104 3381 63113
rect 3339 63064 3340 63104
rect 3380 63064 3381 63104
rect 3339 63055 3381 63064
rect 3340 61601 3380 63055
rect 3436 61685 3476 63148
rect 3435 61676 3477 61685
rect 3435 61636 3436 61676
rect 3476 61636 3477 61676
rect 3435 61627 3477 61636
rect 3339 61592 3381 61601
rect 3339 61552 3340 61592
rect 3380 61552 3381 61592
rect 3339 61543 3381 61552
rect 3340 61458 3380 61543
rect 3436 61542 3476 61627
rect 3435 61424 3477 61433
rect 3435 61384 3436 61424
rect 3476 61384 3477 61424
rect 3435 61375 3477 61384
rect 3244 61048 3380 61088
rect 3148 60929 3188 61014
rect 3147 60920 3189 60929
rect 3147 60880 3148 60920
rect 3188 60880 3189 60920
rect 3147 60871 3189 60880
rect 3244 60920 3284 60929
rect 3244 60668 3284 60880
rect 2956 60628 3284 60668
rect 3051 60080 3093 60089
rect 3051 60040 3052 60080
rect 3092 60040 3093 60080
rect 3051 60031 3093 60040
rect 3052 59946 3092 60031
rect 3244 59585 3284 60628
rect 3243 59576 3285 59585
rect 3243 59536 3244 59576
rect 3284 59536 3285 59576
rect 3243 59527 3285 59536
rect 2763 59408 2805 59417
rect 2763 59368 2764 59408
rect 2804 59368 2805 59408
rect 2763 59359 2805 59368
rect 3148 59408 3188 59417
rect 3148 59324 3188 59368
rect 3243 59408 3285 59417
rect 3243 59368 3244 59408
rect 3284 59368 3285 59408
rect 3243 59359 3285 59368
rect 3052 59284 3188 59324
rect 2764 59240 2804 59251
rect 2764 59165 2804 59200
rect 2763 59156 2805 59165
rect 2763 59116 2764 59156
rect 2804 59116 2805 59156
rect 2763 59107 2805 59116
rect 2667 58820 2709 58829
rect 2667 58780 2668 58820
rect 2708 58780 2709 58820
rect 2667 58771 2709 58780
rect 2668 58568 2708 58771
rect 2668 58519 2708 58528
rect 2860 58400 2900 58409
rect 3052 58400 3092 59284
rect 3147 59156 3189 59165
rect 3147 59116 3148 59156
rect 3188 59116 3189 59156
rect 3147 59107 3189 59116
rect 3148 58736 3188 59107
rect 3148 58687 3188 58696
rect 2900 58360 3092 58400
rect 2860 58351 2900 58360
rect 3244 58073 3284 59359
rect 3340 58232 3380 61048
rect 3436 58568 3476 61375
rect 3532 60248 3572 63223
rect 3916 63104 3956 63307
rect 4204 63113 4244 63727
rect 4203 63104 4245 63113
rect 3956 63064 4148 63104
rect 3916 63055 3956 63064
rect 3688 62012 4056 62021
rect 3728 61972 3770 62012
rect 3810 61972 3852 62012
rect 3892 61972 3934 62012
rect 3974 61972 4016 62012
rect 3688 61963 4056 61972
rect 3723 61676 3765 61685
rect 3723 61636 3724 61676
rect 3764 61636 3765 61676
rect 3723 61627 3765 61636
rect 3724 60920 3764 61627
rect 3916 61592 3956 61601
rect 4108 61592 4148 63064
rect 4203 63064 4204 63104
rect 4244 63064 4245 63104
rect 4203 63055 4245 63064
rect 4203 62432 4245 62441
rect 4203 62392 4204 62432
rect 4244 62392 4245 62432
rect 4203 62383 4245 62392
rect 4300 62432 4340 64576
rect 4395 64616 4437 64625
rect 4395 64576 4396 64616
rect 4436 64576 4437 64616
rect 4395 64567 4437 64576
rect 4492 64373 4532 65239
rect 4491 64364 4533 64373
rect 4491 64324 4492 64364
rect 4532 64324 4533 64364
rect 4491 64315 4533 64324
rect 4492 63944 4532 63953
rect 4588 63944 4628 66079
rect 4684 65549 4724 66088
rect 5164 66142 5204 66163
rect 5164 66077 5204 66102
rect 4779 66044 4821 66053
rect 4779 66004 4780 66044
rect 4820 66004 4821 66044
rect 4779 65995 4821 66004
rect 4683 65540 4725 65549
rect 4683 65500 4684 65540
rect 4724 65500 4725 65540
rect 4683 65491 4725 65500
rect 4532 63904 4628 63944
rect 4395 63692 4437 63701
rect 4395 63652 4396 63692
rect 4436 63652 4437 63692
rect 4395 63643 4437 63652
rect 4396 63118 4436 63643
rect 4492 63365 4532 63904
rect 4491 63356 4533 63365
rect 4491 63316 4492 63356
rect 4532 63316 4533 63356
rect 4491 63307 4533 63316
rect 4587 63272 4629 63281
rect 4587 63232 4588 63272
rect 4628 63232 4629 63272
rect 4587 63223 4629 63232
rect 4396 63069 4436 63078
rect 4588 63020 4628 63223
rect 4588 62971 4628 62980
rect 4683 63020 4725 63029
rect 4683 62980 4684 63020
rect 4724 62980 4725 63020
rect 4683 62971 4725 62980
rect 4588 62432 4628 62441
rect 4300 62392 4588 62432
rect 4204 62298 4244 62383
rect 3956 61552 4148 61592
rect 3916 61543 3956 61552
rect 4108 60920 4148 61552
rect 4204 60920 4244 60929
rect 4108 60880 4204 60920
rect 3628 60836 3668 60847
rect 3628 60761 3668 60796
rect 3627 60752 3669 60761
rect 3627 60712 3628 60752
rect 3668 60712 3669 60752
rect 3627 60703 3669 60712
rect 3724 60677 3764 60880
rect 4204 60871 4244 60880
rect 3723 60668 3765 60677
rect 3723 60628 3724 60668
rect 3764 60628 3765 60668
rect 3723 60619 3765 60628
rect 4107 60668 4149 60677
rect 4107 60628 4108 60668
rect 4148 60628 4149 60668
rect 4107 60619 4149 60628
rect 3688 60500 4056 60509
rect 3728 60460 3770 60500
rect 3810 60460 3852 60500
rect 3892 60460 3934 60500
rect 3974 60460 4016 60500
rect 3688 60451 4056 60460
rect 3532 60208 3764 60248
rect 3724 59417 3764 60208
rect 3723 59408 3765 59417
rect 3723 59368 3724 59408
rect 3764 59368 3765 59408
rect 3723 59359 3765 59368
rect 3628 59324 3668 59333
rect 3628 59165 3668 59284
rect 3724 59274 3764 59359
rect 3627 59156 3669 59165
rect 3627 59116 3628 59156
rect 3668 59116 3669 59156
rect 3627 59107 3669 59116
rect 3688 58988 4056 58997
rect 3728 58948 3770 58988
rect 3810 58948 3852 58988
rect 3892 58948 3934 58988
rect 3974 58948 4016 58988
rect 3688 58939 4056 58948
rect 4108 58745 4148 60619
rect 4300 60584 4340 62392
rect 4588 62383 4628 62392
rect 4684 62264 4724 62971
rect 4588 62224 4724 62264
rect 4396 62180 4436 62189
rect 4396 61769 4436 62140
rect 4395 61760 4437 61769
rect 4395 61720 4396 61760
rect 4436 61720 4437 61760
rect 4395 61711 4437 61720
rect 4396 61597 4436 61606
rect 4396 61097 4436 61557
rect 4588 61424 4628 62224
rect 4683 61760 4725 61769
rect 4683 61720 4684 61760
rect 4724 61720 4725 61760
rect 4683 61711 4725 61720
rect 4395 61088 4437 61097
rect 4395 61048 4396 61088
rect 4436 61048 4437 61088
rect 4395 61039 4437 61048
rect 4588 60920 4628 61384
rect 4204 60544 4340 60584
rect 4396 60880 4628 60920
rect 4684 60915 4724 61711
rect 4204 60089 4244 60544
rect 4203 60080 4245 60089
rect 4203 60040 4204 60080
rect 4244 60040 4245 60080
rect 4203 60031 4245 60040
rect 4300 60080 4340 60089
rect 4203 59660 4245 59669
rect 4203 59620 4204 59660
rect 4244 59620 4245 59660
rect 4203 59611 4245 59620
rect 4204 59408 4244 59611
rect 4204 59249 4244 59368
rect 4203 59240 4245 59249
rect 4203 59200 4204 59240
rect 4244 59200 4245 59240
rect 4203 59191 4245 59200
rect 4300 58829 4340 60040
rect 4299 58820 4341 58829
rect 4299 58780 4300 58820
rect 4340 58780 4341 58820
rect 4299 58771 4341 58780
rect 4107 58736 4149 58745
rect 4107 58696 4108 58736
rect 4148 58696 4149 58736
rect 4107 58687 4149 58696
rect 3531 58568 3573 58577
rect 3436 58528 3532 58568
rect 3572 58528 3573 58568
rect 3531 58519 3573 58528
rect 3532 58434 3572 58519
rect 3340 58192 3572 58232
rect 3243 58064 3285 58073
rect 3243 58024 3244 58064
rect 3284 58024 3285 58064
rect 3243 58015 3285 58024
rect 3435 58064 3477 58073
rect 3435 58024 3436 58064
rect 3476 58024 3477 58064
rect 3435 58015 3477 58024
rect 2572 57896 2612 57905
rect 3148 57896 3188 57905
rect 3340 57896 3380 57905
rect 2612 57856 2708 57896
rect 2572 57847 2612 57856
rect 2571 57056 2613 57065
rect 2571 57016 2572 57056
rect 2612 57016 2613 57056
rect 2571 57007 2613 57016
rect 2572 55544 2612 57007
rect 2668 56729 2708 57856
rect 3188 57856 3284 57896
rect 3148 57847 3188 57856
rect 3244 57737 3284 57856
rect 3340 57821 3380 57856
rect 3436 57896 3476 58015
rect 3436 57847 3476 57856
rect 3339 57812 3381 57821
rect 3339 57772 3340 57812
rect 3380 57772 3381 57812
rect 3339 57763 3381 57772
rect 3243 57728 3285 57737
rect 3243 57688 3244 57728
rect 3284 57688 3285 57728
rect 3243 57679 3285 57688
rect 2764 57644 2804 57653
rect 2804 57604 3092 57644
rect 2764 57595 2804 57604
rect 2763 57308 2805 57317
rect 2763 57268 2764 57308
rect 2804 57268 2805 57308
rect 2763 57259 2805 57268
rect 2764 57174 2804 57259
rect 2859 57056 2901 57065
rect 2859 57016 2860 57056
rect 2900 57016 2901 57056
rect 2859 57007 2901 57016
rect 3052 57056 3092 57604
rect 3052 57007 3092 57016
rect 3148 57056 3188 57065
rect 2667 56720 2709 56729
rect 2667 56680 2668 56720
rect 2708 56680 2709 56720
rect 2667 56671 2709 56680
rect 2860 56384 2900 57007
rect 3051 56888 3093 56897
rect 3051 56848 3052 56888
rect 3092 56848 3093 56888
rect 3051 56839 3093 56848
rect 3052 56552 3092 56839
rect 3052 56503 3092 56512
rect 2860 56335 2900 56344
rect 3148 56300 3188 57016
rect 3244 56897 3284 57679
rect 3340 57317 3380 57763
rect 3436 57728 3476 57737
rect 3436 57653 3476 57688
rect 3436 57644 3484 57653
rect 3436 57604 3443 57644
rect 3483 57604 3484 57644
rect 3442 57595 3484 57604
rect 3339 57308 3381 57317
rect 3339 57268 3340 57308
rect 3380 57268 3381 57308
rect 3339 57259 3381 57268
rect 3532 57224 3572 58192
rect 4108 58064 4148 58073
rect 4148 58024 4340 58064
rect 4108 58015 4148 58024
rect 3628 57896 3668 57905
rect 3628 57653 3668 57856
rect 3723 57896 3765 57905
rect 3723 57856 3724 57896
rect 3764 57856 3765 57896
rect 3723 57847 3765 57856
rect 3916 57896 3956 57907
rect 3724 57762 3764 57847
rect 3916 57821 3956 57856
rect 4012 57896 4052 57905
rect 3915 57812 3957 57821
rect 3915 57772 3916 57812
rect 3956 57772 3957 57812
rect 3915 57763 3957 57772
rect 4012 57653 4052 57856
rect 4113 57896 4153 57905
rect 4113 57737 4153 57856
rect 4112 57728 4154 57737
rect 4112 57688 4113 57728
rect 4153 57688 4154 57728
rect 4112 57679 4154 57688
rect 3627 57644 3669 57653
rect 3627 57604 3628 57644
rect 3668 57604 3669 57644
rect 3627 57595 3669 57604
rect 4011 57644 4053 57653
rect 4011 57604 4012 57644
rect 4052 57604 4053 57644
rect 4011 57595 4053 57604
rect 3688 57476 4056 57485
rect 3728 57436 3770 57476
rect 3810 57436 3852 57476
rect 3892 57436 3934 57476
rect 3974 57436 4016 57476
rect 3688 57427 4056 57436
rect 3532 57184 3668 57224
rect 3628 57140 3668 57184
rect 3532 57056 3572 57065
rect 3243 56888 3285 56897
rect 3243 56848 3244 56888
rect 3284 56848 3285 56888
rect 3243 56839 3285 56848
rect 3435 56384 3477 56393
rect 3435 56344 3436 56384
rect 3476 56344 3477 56384
rect 3435 56335 3477 56344
rect 2956 56260 3188 56300
rect 2764 55712 2804 55721
rect 2612 55504 2708 55544
rect 2572 55495 2612 55504
rect 2668 54872 2708 55504
rect 2764 55385 2804 55672
rect 2763 55376 2805 55385
rect 2763 55336 2764 55376
rect 2804 55336 2805 55376
rect 2763 55327 2805 55336
rect 2091 50924 2133 50933
rect 2091 50884 2092 50924
rect 2132 50884 2133 50924
rect 2091 50875 2133 50884
rect 1899 46808 1941 46817
rect 1899 46768 1900 46808
rect 1940 46768 1941 46808
rect 1899 46759 1941 46768
rect 1996 44960 2036 44969
rect 1996 44045 2036 44920
rect 1995 44036 2037 44045
rect 1995 43996 1996 44036
rect 2036 43996 2037 44036
rect 1995 43987 2037 43996
rect 1803 41936 1845 41945
rect 1803 41896 1804 41936
rect 1844 41896 1845 41936
rect 1803 41887 1845 41896
rect 1803 41264 1845 41273
rect 1803 41224 1804 41264
rect 1844 41224 1845 41264
rect 1803 41215 1845 41224
rect 1804 41130 1844 41215
rect 1899 40424 1941 40433
rect 1899 40384 1900 40424
rect 1940 40384 1941 40424
rect 1899 40375 1941 40384
rect 1707 37568 1749 37577
rect 1707 37528 1708 37568
rect 1748 37528 1749 37568
rect 1707 37519 1749 37528
rect 1515 36728 1557 36737
rect 1515 36688 1516 36728
rect 1556 36688 1557 36728
rect 1515 36679 1557 36688
rect 1419 34460 1461 34469
rect 1419 34420 1420 34460
rect 1460 34420 1461 34460
rect 1419 34411 1461 34420
rect 1268 33664 1364 33704
rect 1228 33655 1268 33664
rect 1228 32822 1268 32831
rect 1227 32782 1228 32789
rect 1268 32782 1269 32789
rect 1227 32780 1269 32782
rect 1227 32740 1228 32780
rect 1268 32740 1269 32780
rect 1227 32731 1269 32740
rect 1228 32687 1268 32731
rect 1516 32453 1556 36679
rect 1900 36056 1940 40375
rect 1996 36905 2036 43987
rect 2092 42953 2132 50875
rect 2188 47069 2228 53311
rect 2476 52520 2516 53320
rect 2572 54832 2668 54872
rect 2572 53201 2612 54832
rect 2668 54823 2708 54832
rect 2667 54704 2709 54713
rect 2667 54664 2668 54704
rect 2708 54664 2709 54704
rect 2667 54655 2709 54664
rect 2668 54032 2708 54655
rect 2668 53983 2708 53992
rect 2764 53360 2804 55327
rect 2859 55124 2901 55133
rect 2859 55084 2860 55124
rect 2900 55084 2901 55124
rect 2859 55075 2901 55084
rect 2860 55040 2900 55075
rect 2860 54989 2900 55000
rect 2956 54200 2996 56260
rect 3436 56250 3476 56335
rect 3532 55973 3572 57016
rect 3628 56225 3668 57100
rect 4108 57056 4148 57065
rect 4300 57056 4340 58024
rect 4148 57016 4340 57056
rect 3627 56216 3669 56225
rect 3627 56176 3628 56216
rect 3668 56176 3669 56216
rect 3627 56167 3669 56176
rect 3531 55964 3573 55973
rect 3531 55924 3532 55964
rect 3572 55924 3573 55964
rect 3531 55915 3573 55924
rect 3688 55964 4056 55973
rect 3728 55924 3770 55964
rect 3810 55924 3852 55964
rect 3892 55924 3934 55964
rect 3974 55924 4016 55964
rect 3688 55915 4056 55924
rect 3052 55756 3572 55796
rect 3052 55040 3092 55756
rect 3244 55553 3284 55638
rect 3148 55544 3188 55553
rect 3148 55040 3188 55504
rect 3243 55544 3285 55553
rect 3243 55504 3244 55544
rect 3284 55504 3285 55544
rect 3243 55495 3285 55504
rect 3436 55544 3476 55553
rect 3436 55460 3476 55504
rect 3532 55544 3572 55756
rect 4011 55712 4053 55721
rect 4011 55672 4012 55712
rect 4052 55672 4053 55712
rect 4011 55663 4053 55672
rect 3916 55553 3956 55638
rect 3633 55544 3673 55553
rect 3532 55495 3572 55504
rect 3628 55504 3633 55544
rect 3628 55495 3673 55504
rect 3915 55544 3957 55553
rect 3915 55504 3916 55544
rect 3956 55504 3957 55544
rect 3915 55495 3957 55504
rect 4012 55544 4052 55663
rect 4012 55495 4052 55504
rect 3340 55420 3476 55460
rect 3340 55133 3380 55420
rect 3628 55385 3668 55495
rect 3532 55376 3572 55385
rect 3339 55124 3381 55133
rect 3339 55084 3340 55124
rect 3380 55084 3476 55124
rect 3339 55075 3381 55084
rect 3148 55000 3284 55040
rect 3052 54991 3092 55000
rect 3148 54872 3188 54883
rect 3148 54797 3188 54832
rect 3147 54788 3189 54797
rect 3147 54748 3148 54788
rect 3188 54748 3189 54788
rect 3147 54739 3189 54748
rect 3244 54704 3284 55000
rect 3340 54881 3380 54966
rect 3339 54872 3381 54881
rect 3339 54832 3340 54872
rect 3380 54832 3381 54872
rect 3339 54823 3381 54832
rect 3244 54664 3380 54704
rect 2956 54160 3284 54200
rect 3148 54032 3188 54041
rect 2860 53948 2900 53957
rect 3148 53948 3188 53992
rect 2900 53908 3188 53948
rect 3244 54032 3284 54160
rect 2860 53899 2900 53908
rect 3244 53705 3284 53992
rect 3243 53696 3285 53705
rect 3243 53656 3244 53696
rect 3284 53656 3285 53696
rect 3243 53647 3285 53656
rect 3052 53528 3092 53537
rect 3340 53528 3380 54664
rect 3092 53488 3380 53528
rect 3052 53479 3092 53488
rect 2956 53360 2996 53369
rect 2764 53320 2956 53360
rect 2956 53311 2996 53320
rect 3148 53360 3188 53369
rect 2571 53192 2613 53201
rect 2571 53152 2572 53192
rect 2612 53152 2613 53192
rect 2571 53143 2613 53152
rect 2955 53192 2997 53201
rect 2955 53152 2956 53192
rect 2996 53152 2997 53192
rect 2955 53143 2997 53152
rect 2668 53108 2708 53117
rect 2668 52940 2708 53068
rect 2668 52900 2804 52940
rect 2668 52520 2708 52529
rect 2476 52480 2668 52520
rect 2668 51848 2708 52480
rect 2572 51808 2668 51848
rect 2475 51344 2517 51353
rect 2475 51304 2476 51344
rect 2516 51304 2517 51344
rect 2475 51295 2517 51304
rect 2476 51008 2516 51295
rect 2283 50756 2325 50765
rect 2283 50716 2284 50756
rect 2324 50716 2325 50756
rect 2283 50707 2325 50716
rect 2284 48329 2324 50707
rect 2476 50420 2516 50968
rect 2572 50588 2612 51808
rect 2668 51799 2708 51808
rect 2764 51101 2804 52900
rect 2859 52352 2901 52361
rect 2859 52312 2860 52352
rect 2900 52312 2901 52352
rect 2859 52303 2901 52312
rect 2860 51857 2900 52303
rect 2859 51848 2901 51857
rect 2859 51808 2860 51848
rect 2900 51808 2901 51848
rect 2859 51799 2901 51808
rect 2859 51680 2901 51689
rect 2859 51640 2860 51680
rect 2900 51640 2901 51680
rect 2859 51631 2901 51640
rect 2763 51092 2805 51101
rect 2763 51052 2764 51092
rect 2804 51052 2805 51092
rect 2763 51043 2805 51052
rect 2860 51017 2900 51631
rect 2859 51008 2901 51017
rect 2859 50968 2860 51008
rect 2900 50968 2901 51008
rect 2859 50959 2901 50968
rect 2667 50840 2709 50849
rect 2860 50840 2900 50849
rect 2667 50800 2668 50840
rect 2708 50800 2709 50840
rect 2667 50791 2709 50800
rect 2764 50800 2860 50840
rect 2668 50706 2708 50791
rect 2572 50548 2708 50588
rect 2476 50380 2612 50420
rect 2572 50336 2612 50380
rect 2572 50287 2612 50296
rect 2668 50168 2708 50548
rect 2572 50128 2708 50168
rect 2379 50084 2421 50093
rect 2379 50044 2380 50084
rect 2420 50044 2421 50084
rect 2379 50035 2421 50044
rect 2380 49950 2420 50035
rect 2572 49160 2612 50128
rect 2667 49412 2709 49421
rect 2667 49372 2668 49412
rect 2708 49372 2709 49412
rect 2667 49363 2709 49372
rect 2668 49278 2708 49363
rect 2572 49120 2708 49160
rect 2572 48824 2612 48833
rect 2476 48784 2572 48824
rect 2283 48320 2325 48329
rect 2283 48280 2284 48320
rect 2324 48280 2325 48320
rect 2283 48271 2325 48280
rect 2476 48077 2516 48784
rect 2572 48775 2612 48784
rect 2668 48656 2708 49120
rect 2764 48749 2804 50800
rect 2860 50791 2900 50800
rect 2859 50084 2901 50093
rect 2859 50044 2860 50084
rect 2900 50044 2901 50084
rect 2859 50035 2901 50044
rect 2860 49510 2900 50035
rect 2860 49461 2900 49470
rect 2859 49328 2901 49337
rect 2859 49288 2860 49328
rect 2900 49288 2901 49328
rect 2859 49279 2901 49288
rect 2763 48740 2805 48749
rect 2763 48700 2764 48740
rect 2804 48700 2805 48740
rect 2763 48691 2805 48700
rect 2572 48616 2708 48656
rect 2475 48068 2517 48077
rect 2475 48028 2476 48068
rect 2516 48028 2517 48068
rect 2475 48019 2517 48028
rect 2476 47984 2516 48019
rect 2476 47933 2516 47944
rect 2379 47900 2421 47909
rect 2379 47860 2380 47900
rect 2420 47860 2421 47900
rect 2379 47851 2421 47860
rect 2187 47060 2229 47069
rect 2187 47020 2188 47060
rect 2228 47020 2229 47060
rect 2187 47011 2229 47020
rect 2188 46649 2228 47011
rect 2187 46640 2229 46649
rect 2187 46600 2188 46640
rect 2228 46600 2229 46640
rect 2187 46591 2229 46600
rect 2380 46472 2420 47851
rect 2475 47816 2517 47825
rect 2475 47776 2476 47816
rect 2516 47776 2517 47816
rect 2475 47767 2517 47776
rect 2476 47312 2516 47767
rect 2572 47741 2612 48616
rect 2763 48572 2805 48581
rect 2763 48532 2764 48572
rect 2804 48532 2805 48572
rect 2763 48523 2805 48532
rect 2764 48438 2804 48523
rect 2860 48320 2900 49279
rect 2956 48413 2996 53143
rect 3148 53108 3188 53320
rect 3243 53360 3285 53369
rect 3243 53320 3244 53360
rect 3284 53320 3285 53360
rect 3243 53311 3285 53320
rect 3244 53226 3284 53311
rect 3436 53108 3476 55084
rect 3148 53068 3476 53108
rect 3532 52688 3572 55336
rect 3627 55376 3669 55385
rect 3627 55336 3628 55376
rect 3668 55336 3669 55376
rect 3627 55327 3669 55336
rect 3688 54452 4056 54461
rect 3728 54412 3770 54452
rect 3810 54412 3852 54452
rect 3892 54412 3934 54452
rect 3974 54412 4016 54452
rect 3688 54403 4056 54412
rect 3723 54284 3765 54293
rect 3723 54244 3724 54284
rect 3764 54244 3765 54284
rect 3723 54235 3765 54244
rect 3724 54116 3764 54235
rect 3724 54067 3764 54076
rect 3628 54032 3668 54043
rect 4108 54032 4148 57016
rect 4203 55628 4245 55637
rect 4203 55588 4204 55628
rect 4244 55588 4245 55628
rect 4203 55579 4245 55588
rect 4204 55376 4244 55579
rect 4204 55327 4244 55336
rect 4204 54032 4244 54041
rect 4108 53992 4204 54032
rect 3628 53957 3668 53992
rect 4204 53983 4244 53992
rect 3627 53948 3669 53957
rect 3627 53908 3628 53948
rect 3668 53908 3669 53948
rect 3627 53899 3669 53908
rect 4299 53864 4341 53873
rect 4299 53824 4300 53864
rect 4340 53824 4341 53864
rect 4299 53815 4341 53824
rect 4107 53780 4149 53789
rect 4107 53740 4108 53780
rect 4148 53740 4149 53780
rect 4107 53731 4149 53740
rect 3688 52940 4056 52949
rect 3728 52900 3770 52940
rect 3810 52900 3852 52940
rect 3892 52900 3934 52940
rect 3974 52900 4016 52940
rect 3688 52891 4056 52900
rect 3724 52688 3764 52697
rect 3532 52648 3668 52688
rect 3052 52520 3092 52529
rect 3052 52016 3092 52480
rect 3340 52520 3380 52529
rect 3244 52352 3284 52361
rect 3052 51967 3092 51976
rect 3148 52312 3244 52352
rect 3051 51764 3093 51773
rect 3051 51724 3052 51764
rect 3092 51724 3093 51764
rect 3051 51715 3093 51724
rect 3052 51176 3092 51715
rect 3052 51127 3092 51136
rect 3052 51008 3092 51017
rect 3148 51008 3188 52312
rect 3244 52303 3284 52312
rect 3243 51848 3285 51857
rect 3243 51803 3244 51848
rect 3284 51803 3285 51848
rect 3243 51799 3285 51803
rect 3244 51713 3284 51799
rect 3340 51689 3380 52480
rect 3532 52520 3572 52529
rect 3532 52361 3572 52480
rect 3531 52352 3573 52361
rect 3531 52312 3532 52352
rect 3572 52312 3573 52352
rect 3531 52303 3573 52312
rect 3628 52100 3668 52648
rect 3764 52648 3956 52688
rect 3724 52639 3764 52648
rect 3436 52060 3668 52100
rect 3724 52520 3764 52529
rect 3339 51680 3381 51689
rect 3339 51640 3340 51680
rect 3380 51640 3381 51680
rect 3339 51631 3381 51640
rect 3339 51092 3381 51101
rect 3339 51052 3340 51092
rect 3380 51052 3381 51092
rect 3339 51043 3381 51052
rect 3092 50968 3188 51008
rect 3340 51008 3380 51043
rect 3052 50959 3092 50968
rect 3340 50957 3380 50968
rect 3243 50084 3285 50093
rect 3243 50044 3244 50084
rect 3284 50044 3285 50084
rect 3243 50035 3285 50044
rect 3051 48992 3093 49001
rect 3051 48952 3052 48992
rect 3092 48952 3093 48992
rect 3051 48943 3093 48952
rect 2955 48404 2997 48413
rect 2955 48364 2956 48404
rect 2996 48364 2997 48404
rect 2955 48355 2997 48364
rect 2764 48280 2900 48320
rect 2668 47816 2708 47825
rect 2571 47732 2613 47741
rect 2571 47692 2572 47732
rect 2612 47692 2613 47732
rect 2571 47683 2613 47692
rect 2476 47263 2516 47272
rect 2572 47396 2612 47405
rect 2476 46472 2516 46481
rect 2380 46432 2476 46472
rect 2476 46423 2516 46432
rect 2187 44792 2229 44801
rect 2187 44752 2188 44792
rect 2228 44752 2229 44792
rect 2187 44743 2229 44752
rect 2091 42944 2133 42953
rect 2091 42904 2092 42944
rect 2132 42904 2133 42944
rect 2091 42895 2133 42904
rect 2091 37736 2133 37745
rect 2091 37696 2092 37736
rect 2132 37696 2133 37736
rect 2091 37687 2133 37696
rect 1995 36896 2037 36905
rect 1995 36856 1996 36896
rect 2036 36856 2037 36896
rect 1995 36847 2037 36856
rect 1995 36056 2037 36065
rect 1900 36016 1996 36056
rect 2036 36016 2037 36056
rect 1995 36007 2037 36016
rect 1899 34964 1941 34973
rect 1899 34924 1900 34964
rect 1940 34924 1941 34964
rect 1899 34915 1941 34924
rect 1900 34830 1940 34915
rect 1515 32444 1557 32453
rect 1515 32404 1516 32444
rect 1556 32404 1557 32444
rect 1515 32395 1557 32404
rect 1323 32360 1365 32369
rect 1323 32320 1324 32360
rect 1364 32320 1365 32360
rect 1323 32311 1365 32320
rect 1131 32276 1173 32285
rect 1131 32236 1132 32276
rect 1172 32236 1173 32276
rect 1131 32227 1173 32236
rect 1132 30857 1172 32227
rect 1228 32192 1268 32201
rect 1324 32192 1364 32311
rect 1268 32152 1364 32192
rect 1228 32143 1268 32152
rect 1899 32108 1941 32117
rect 1899 32068 1900 32108
rect 1940 32068 1941 32108
rect 1899 32059 1941 32068
rect 1131 30848 1173 30857
rect 1131 30808 1132 30848
rect 1172 30808 1173 30848
rect 1131 30799 1173 30808
rect 1804 30848 1844 30859
rect 1804 30773 1844 30808
rect 1803 30764 1845 30773
rect 1803 30724 1804 30764
rect 1844 30724 1845 30764
rect 1803 30715 1845 30724
rect 1804 30008 1844 30715
rect 1419 29672 1461 29681
rect 1419 29632 1420 29672
rect 1460 29632 1461 29672
rect 1419 29623 1461 29632
rect 1227 28160 1269 28169
rect 1227 28120 1228 28160
rect 1268 28120 1269 28160
rect 1227 28111 1269 28120
rect 1228 27665 1268 28111
rect 1227 27656 1269 27665
rect 1227 27616 1228 27656
rect 1268 27616 1269 27656
rect 1227 27607 1269 27616
rect 1323 26984 1365 26993
rect 1323 26944 1324 26984
rect 1364 26944 1365 26984
rect 1323 26935 1365 26944
rect 1227 26816 1269 26825
rect 1227 26776 1228 26816
rect 1268 26776 1269 26816
rect 1227 26767 1269 26776
rect 1324 26816 1364 26935
rect 1324 26767 1364 26776
rect 1420 26816 1460 29623
rect 1804 29336 1844 29968
rect 1804 28496 1844 29296
rect 1804 28447 1844 28456
rect 1708 28160 1748 28169
rect 1515 27908 1557 27917
rect 1515 27868 1516 27908
rect 1556 27868 1557 27908
rect 1515 27859 1557 27868
rect 1420 26767 1460 26776
rect 1516 26816 1556 27859
rect 1708 27656 1748 28120
rect 1900 27992 1940 32059
rect 1996 30101 2036 36007
rect 2092 35132 2132 37687
rect 2092 35083 2132 35092
rect 2091 32780 2133 32789
rect 2091 32740 2092 32780
rect 2132 32740 2133 32780
rect 2091 32731 2133 32740
rect 2092 31604 2132 32731
rect 2188 32201 2228 44743
rect 2572 44129 2612 47356
rect 2668 47312 2708 47776
rect 2668 47144 2708 47272
rect 2764 47312 2804 48280
rect 2764 47263 2804 47272
rect 2860 47984 2900 47993
rect 2860 47144 2900 47944
rect 3052 47984 3092 48943
rect 3148 48824 3188 48833
rect 3148 48581 3188 48784
rect 3244 48824 3284 50035
rect 3340 49496 3380 49505
rect 3436 49496 3476 52060
rect 3724 52016 3764 52480
rect 3532 51976 3764 52016
rect 3820 52520 3860 52529
rect 3532 51092 3572 51976
rect 3723 51848 3765 51857
rect 3723 51808 3724 51848
rect 3764 51808 3765 51848
rect 3723 51799 3765 51808
rect 3724 51714 3764 51799
rect 3820 51596 3860 52480
rect 3916 51773 3956 52648
rect 3915 51764 3957 51773
rect 3915 51724 3916 51764
rect 3956 51724 3957 51764
rect 3915 51715 3957 51724
rect 4108 51680 4148 53731
rect 4300 53528 4340 53815
rect 4396 53789 4436 60880
rect 4684 60866 4724 60875
rect 4780 60509 4820 65995
rect 5356 65960 5396 65969
rect 4928 65792 5296 65801
rect 4968 65752 5010 65792
rect 5050 65752 5092 65792
rect 5132 65752 5174 65792
rect 5214 65752 5256 65792
rect 4928 65743 5296 65752
rect 5356 65549 5396 65920
rect 5452 65633 5492 70699
rect 5548 70421 5588 71632
rect 5740 71513 5780 71968
rect 5644 71504 5684 71513
rect 5644 70832 5684 71464
rect 5739 71504 5781 71513
rect 5739 71464 5740 71504
rect 5780 71464 5781 71504
rect 5739 71455 5781 71464
rect 5644 70792 5972 70832
rect 5643 70664 5685 70673
rect 5643 70624 5644 70664
rect 5684 70624 5685 70664
rect 5643 70615 5685 70624
rect 5644 70530 5684 70615
rect 5835 70580 5877 70589
rect 5835 70540 5836 70580
rect 5876 70540 5877 70580
rect 5835 70531 5877 70540
rect 5547 70412 5589 70421
rect 5547 70372 5548 70412
rect 5588 70372 5589 70412
rect 5547 70363 5589 70372
rect 5836 69992 5876 70531
rect 5643 69320 5685 69329
rect 5643 69280 5644 69320
rect 5684 69280 5685 69320
rect 5643 69271 5685 69280
rect 5547 68648 5589 68657
rect 5547 68608 5548 68648
rect 5588 68608 5589 68648
rect 5547 68599 5589 68608
rect 5451 65624 5493 65633
rect 5451 65584 5452 65624
rect 5492 65584 5493 65624
rect 5451 65575 5493 65584
rect 5355 65540 5397 65549
rect 5355 65500 5356 65540
rect 5396 65500 5397 65540
rect 5355 65491 5397 65500
rect 5451 65456 5493 65465
rect 5451 65416 5452 65456
rect 5492 65416 5493 65456
rect 5451 65407 5493 65416
rect 5452 64616 5492 65407
rect 5452 64567 5492 64576
rect 4928 64280 5296 64289
rect 4968 64240 5010 64280
rect 5050 64240 5092 64280
rect 5132 64240 5174 64280
rect 5214 64240 5256 64280
rect 4928 64231 5296 64240
rect 4971 64112 5013 64121
rect 4971 64072 4972 64112
rect 5012 64072 5013 64112
rect 4971 64063 5013 64072
rect 4972 63939 5012 64063
rect 5163 64028 5205 64037
rect 5163 63988 5164 64028
rect 5204 63988 5205 64028
rect 5163 63979 5205 63988
rect 4972 63890 5012 63899
rect 5164 63894 5204 63979
rect 5355 63356 5397 63365
rect 5355 63316 5356 63356
rect 5396 63316 5397 63356
rect 5355 63307 5397 63316
rect 4928 62768 5296 62777
rect 4968 62728 5010 62768
rect 5050 62728 5092 62768
rect 5132 62728 5174 62768
rect 5214 62728 5256 62768
rect 4928 62719 5296 62728
rect 5356 61601 5396 63307
rect 5451 62936 5493 62945
rect 5451 62896 5452 62936
rect 5492 62896 5493 62936
rect 5451 62887 5493 62896
rect 5355 61592 5397 61601
rect 5355 61552 5356 61592
rect 5396 61552 5397 61592
rect 5355 61543 5397 61552
rect 5356 61458 5396 61543
rect 5452 61340 5492 62887
rect 5356 61300 5492 61340
rect 4928 61256 5296 61265
rect 4968 61216 5010 61256
rect 5050 61216 5092 61256
rect 5132 61216 5174 61256
rect 5214 61216 5256 61256
rect 4928 61207 5296 61216
rect 4876 61004 4916 61013
rect 4779 60500 4821 60509
rect 4779 60460 4780 60500
rect 4820 60460 4821 60500
rect 4779 60451 4821 60460
rect 4876 60173 4916 60964
rect 4875 60164 4917 60173
rect 4875 60124 4876 60164
rect 4916 60124 4917 60164
rect 4875 60115 4917 60124
rect 4492 59912 4532 59921
rect 4532 59872 4724 59912
rect 4492 59863 4532 59872
rect 4684 59403 4724 59872
rect 4928 59744 5296 59753
rect 4968 59704 5010 59744
rect 5050 59704 5092 59744
rect 5132 59704 5174 59744
rect 5214 59704 5256 59744
rect 4928 59695 5296 59704
rect 4875 59492 4917 59501
rect 4875 59452 4876 59492
rect 4916 59452 4917 59492
rect 4875 59443 4917 59452
rect 4684 59354 4724 59363
rect 4876 59358 4916 59443
rect 5356 58997 5396 61300
rect 5451 61088 5493 61097
rect 5451 61048 5452 61088
rect 5492 61048 5493 61088
rect 5451 61039 5493 61048
rect 5452 60920 5492 61039
rect 5452 60845 5492 60880
rect 5451 60836 5493 60845
rect 5451 60796 5452 60836
rect 5492 60796 5493 60836
rect 5451 60787 5493 60796
rect 5452 60756 5492 60787
rect 5451 59408 5493 59417
rect 5451 59368 5452 59408
rect 5492 59368 5493 59408
rect 5451 59359 5493 59368
rect 5355 58988 5397 58997
rect 5355 58948 5356 58988
rect 5396 58948 5397 58988
rect 5355 58939 5397 58948
rect 4779 58820 4821 58829
rect 4779 58780 4780 58820
rect 4820 58780 4821 58820
rect 4779 58771 4821 58780
rect 4491 58736 4533 58745
rect 4491 58696 4492 58736
rect 4532 58696 4533 58736
rect 4491 58687 4533 58696
rect 4492 56216 4532 58687
rect 4780 58568 4820 58771
rect 4684 58528 4780 58568
rect 4684 57989 4724 58528
rect 4780 58519 4820 58528
rect 5260 58568 5300 58577
rect 4972 58484 5012 58493
rect 5260 58484 5300 58528
rect 5356 58568 5396 58579
rect 5356 58493 5396 58528
rect 5012 58444 5300 58484
rect 5355 58484 5397 58493
rect 5355 58444 5356 58484
rect 5396 58444 5397 58484
rect 4972 58435 5012 58444
rect 5355 58435 5397 58444
rect 4779 58316 4821 58325
rect 4779 58276 4780 58316
rect 4820 58276 4821 58316
rect 4779 58267 4821 58276
rect 4683 57980 4725 57989
rect 4683 57940 4684 57980
rect 4724 57940 4725 57980
rect 4683 57931 4725 57940
rect 4636 57065 4676 57074
rect 4676 57025 4724 57056
rect 4636 57016 4724 57025
rect 4587 56720 4629 56729
rect 4587 56680 4588 56720
rect 4628 56680 4629 56720
rect 4587 56671 4629 56680
rect 4588 56384 4628 56671
rect 4684 56636 4724 57016
rect 4780 56972 4820 58267
rect 4928 58232 5296 58241
rect 4968 58192 5010 58232
rect 5050 58192 5092 58232
rect 5132 58192 5174 58232
rect 5214 58192 5256 58232
rect 4928 58183 5296 58192
rect 5452 58064 5492 59359
rect 5068 58024 5492 58064
rect 4971 57728 5013 57737
rect 4971 57688 4972 57728
rect 5012 57688 5013 57728
rect 4971 57679 5013 57688
rect 4972 57056 5012 57679
rect 4972 57007 5012 57016
rect 5068 57056 5108 58024
rect 5259 57896 5301 57905
rect 5259 57856 5260 57896
rect 5300 57856 5301 57896
rect 5259 57847 5301 57856
rect 5356 57896 5396 57907
rect 5068 57007 5108 57016
rect 4780 56923 4820 56932
rect 5260 56888 5300 57847
rect 5356 57821 5396 57856
rect 5355 57812 5397 57821
rect 5355 57772 5356 57812
rect 5396 57772 5397 57812
rect 5355 57763 5397 57772
rect 5355 57644 5397 57653
rect 5355 57604 5356 57644
rect 5396 57604 5397 57644
rect 5355 57595 5397 57604
rect 5260 56839 5300 56848
rect 4928 56720 5296 56729
rect 4968 56680 5010 56720
rect 5050 56680 5092 56720
rect 5132 56680 5174 56720
rect 5214 56680 5256 56720
rect 4928 56671 5296 56680
rect 4684 56596 4820 56636
rect 4780 56552 4820 56596
rect 4876 56552 4916 56561
rect 4780 56512 4876 56552
rect 4876 56503 4916 56512
rect 5068 56552 5108 56561
rect 5356 56552 5396 57595
rect 5108 56512 5396 56552
rect 5068 56503 5108 56512
rect 4684 56384 4724 56393
rect 4588 56344 4684 56384
rect 4492 56176 4628 56216
rect 4491 56048 4533 56057
rect 4491 56008 4492 56048
rect 4532 56008 4533 56048
rect 4491 55999 4533 56008
rect 4492 55544 4532 55999
rect 4588 55721 4628 56176
rect 4587 55712 4629 55721
rect 4587 55672 4588 55712
rect 4628 55672 4629 55712
rect 4587 55663 4629 55672
rect 4492 55495 4532 55504
rect 4588 54872 4628 54881
rect 4588 54713 4628 54832
rect 4587 54704 4629 54713
rect 4587 54664 4588 54704
rect 4628 54664 4629 54704
rect 4587 54655 4629 54664
rect 4684 54536 4724 56344
rect 5164 56384 5204 56393
rect 5164 55973 5204 56344
rect 5163 55964 5205 55973
rect 5163 55924 5164 55964
rect 5204 55924 5205 55964
rect 5163 55915 5205 55924
rect 5355 55964 5397 55973
rect 5355 55924 5356 55964
rect 5396 55924 5397 55964
rect 5355 55915 5397 55924
rect 4928 55208 5296 55217
rect 4968 55168 5010 55208
rect 5050 55168 5092 55208
rect 5132 55168 5174 55208
rect 5214 55168 5256 55208
rect 4928 55159 5296 55168
rect 5356 54704 5396 55915
rect 5548 55376 5588 68599
rect 5644 66884 5684 69271
rect 5836 69152 5876 69952
rect 5932 69329 5972 70792
rect 6028 70001 6068 72136
rect 6316 71588 6356 71597
rect 6124 71490 6164 71499
rect 6124 71009 6164 71450
rect 6316 71429 6356 71548
rect 6315 71420 6357 71429
rect 6315 71380 6316 71420
rect 6356 71380 6357 71420
rect 6315 71371 6357 71380
rect 6123 71000 6165 71009
rect 6123 70960 6124 71000
rect 6164 70960 6165 71000
rect 6123 70951 6165 70960
rect 6027 69992 6069 70001
rect 6027 69952 6028 69992
rect 6068 69952 6069 69992
rect 6027 69943 6069 69952
rect 6219 69992 6261 70001
rect 6219 69952 6220 69992
rect 6260 69952 6261 69992
rect 6219 69943 6261 69952
rect 6220 69858 6260 69943
rect 6027 69740 6069 69749
rect 6027 69700 6028 69740
rect 6068 69700 6069 69740
rect 6027 69691 6069 69700
rect 6028 69606 6068 69691
rect 5931 69320 5973 69329
rect 5931 69280 5932 69320
rect 5972 69280 5973 69320
rect 5931 69271 5973 69280
rect 6028 69173 6068 69182
rect 5836 69133 6028 69152
rect 5836 69112 6068 69133
rect 5836 67649 5876 69112
rect 6220 68984 6260 68993
rect 6220 68480 6260 68944
rect 6316 68480 6356 68489
rect 6220 68440 6316 68480
rect 6316 68431 6356 68440
rect 6411 68480 6453 68489
rect 6411 68440 6412 68480
rect 6452 68440 6453 68480
rect 6411 68431 6453 68440
rect 6412 68346 6452 68431
rect 6219 67808 6261 67817
rect 6508 67808 6548 73060
rect 6603 71504 6645 71513
rect 6603 71464 6604 71504
rect 6644 71464 6645 71504
rect 6603 71455 6645 71464
rect 6700 71504 6740 71513
rect 6604 71370 6644 71455
rect 6603 71252 6645 71261
rect 6603 71212 6604 71252
rect 6644 71212 6645 71252
rect 6603 71203 6645 71212
rect 6604 69824 6644 71203
rect 6700 69908 6740 71464
rect 6892 71009 6932 76000
rect 6987 74276 7029 74285
rect 6987 74236 6988 74276
rect 7028 74236 7029 74276
rect 6987 74227 7029 74236
rect 6988 73702 7028 74227
rect 6988 73653 7028 73662
rect 7084 73604 7124 83644
rect 7371 83516 7413 83525
rect 7371 83476 7372 83516
rect 7412 83476 7413 83516
rect 7371 83467 7413 83476
rect 7372 83382 7412 83467
rect 7659 82844 7701 82853
rect 7659 82804 7660 82844
rect 7700 82804 7701 82844
rect 7659 82795 7701 82804
rect 7660 74537 7700 82795
rect 7755 75452 7797 75461
rect 7755 75412 7756 75452
rect 7796 75412 7797 75452
rect 7755 75403 7797 75412
rect 7659 74528 7701 74537
rect 7659 74488 7660 74528
rect 7700 74488 7701 74528
rect 7659 74479 7701 74488
rect 7659 74360 7701 74369
rect 7659 74320 7660 74360
rect 7700 74320 7701 74360
rect 7659 74311 7701 74320
rect 6988 73564 7124 73604
rect 6891 71000 6933 71009
rect 6891 70960 6892 71000
rect 6932 70960 6933 71000
rect 6891 70951 6933 70960
rect 6892 70664 6932 70675
rect 6892 70589 6932 70624
rect 6891 70580 6933 70589
rect 6891 70540 6892 70580
rect 6932 70540 6933 70580
rect 6891 70531 6933 70540
rect 6700 69868 6932 69908
rect 6604 69784 6740 69824
rect 6603 69152 6645 69161
rect 6603 69112 6604 69152
rect 6644 69112 6645 69152
rect 6603 69103 6645 69112
rect 6219 67768 6220 67808
rect 6260 67768 6261 67808
rect 6219 67759 6261 67768
rect 6316 67768 6548 67808
rect 5835 67640 5877 67649
rect 5835 67600 5836 67640
rect 5876 67600 5877 67640
rect 5835 67591 5877 67600
rect 6220 67640 6260 67759
rect 5836 66977 5876 67591
rect 6027 67472 6069 67481
rect 6027 67432 6028 67472
rect 6068 67432 6069 67472
rect 6027 67423 6069 67432
rect 6028 67338 6068 67423
rect 6220 67145 6260 67600
rect 6219 67136 6261 67145
rect 6219 67096 6220 67136
rect 6260 67096 6261 67136
rect 6219 67087 6261 67096
rect 5835 66968 5877 66977
rect 6220 66968 6260 66977
rect 5835 66928 5836 66968
rect 5876 66928 5877 66968
rect 5835 66919 5877 66928
rect 6124 66928 6220 66968
rect 5644 66844 5780 66884
rect 5740 66641 5780 66844
rect 5835 66800 5877 66809
rect 6124 66800 6164 66928
rect 6220 66919 6260 66928
rect 5835 66760 5836 66800
rect 5876 66760 5877 66800
rect 5835 66751 5877 66760
rect 6028 66760 6164 66800
rect 5739 66632 5781 66641
rect 5739 66592 5740 66632
rect 5780 66592 5781 66632
rect 5739 66583 5781 66592
rect 5643 66464 5685 66473
rect 5643 66424 5644 66464
rect 5684 66424 5685 66464
rect 5643 66415 5685 66424
rect 5644 65372 5684 66415
rect 5739 66296 5781 66305
rect 5739 66256 5740 66296
rect 5780 66256 5781 66296
rect 5739 66247 5781 66256
rect 5740 65456 5780 66247
rect 5836 66128 5876 66751
rect 5836 66079 5876 66088
rect 5932 66128 5972 66137
rect 5932 65792 5972 66088
rect 6028 65876 6068 66760
rect 6219 66632 6261 66641
rect 6219 66592 6220 66632
rect 6260 66592 6261 66632
rect 6219 66583 6261 66592
rect 6028 65836 6164 65876
rect 5932 65752 6068 65792
rect 5931 65624 5973 65633
rect 5931 65584 5932 65624
rect 5972 65584 5973 65624
rect 5931 65575 5973 65584
rect 5836 65456 5876 65465
rect 5740 65416 5836 65456
rect 5836 65407 5876 65416
rect 5644 65332 5780 65372
rect 5643 64532 5685 64541
rect 5643 64492 5644 64532
rect 5684 64492 5685 64532
rect 5643 64483 5685 64492
rect 5644 64398 5684 64483
rect 5740 64037 5780 65332
rect 5836 64616 5876 64625
rect 5932 64616 5972 65575
rect 5876 64576 5972 64616
rect 5836 64567 5876 64576
rect 5739 64028 5781 64037
rect 5739 63988 5740 64028
rect 5780 63988 5781 64028
rect 5739 63979 5781 63988
rect 5643 63104 5685 63113
rect 5643 63064 5644 63104
rect 5684 63064 5685 63104
rect 5643 63055 5685 63064
rect 5644 62970 5684 63055
rect 5643 61592 5685 61601
rect 5643 61552 5644 61592
rect 5684 61552 5685 61592
rect 5643 61543 5685 61552
rect 5644 56393 5684 61543
rect 5740 59240 5780 63979
rect 5932 62945 5972 64576
rect 6028 63785 6068 65752
rect 6124 65465 6164 65836
rect 6123 65456 6165 65465
rect 6123 65416 6124 65456
rect 6164 65416 6165 65456
rect 6123 65407 6165 65416
rect 6123 65204 6165 65213
rect 6123 65164 6124 65204
rect 6164 65164 6165 65204
rect 6123 65155 6165 65164
rect 6027 63776 6069 63785
rect 6027 63736 6028 63776
rect 6068 63736 6069 63776
rect 6027 63727 6069 63736
rect 5931 62936 5973 62945
rect 5931 62896 5932 62936
rect 5972 62896 5973 62936
rect 5931 62887 5973 62896
rect 5836 62432 5876 62441
rect 6124 62432 6164 65155
rect 6220 63869 6260 66583
rect 6316 66212 6356 67768
rect 6412 66800 6452 66809
rect 6452 66760 6548 66800
rect 6412 66751 6452 66760
rect 6411 66548 6453 66557
rect 6411 66508 6412 66548
rect 6452 66508 6453 66548
rect 6411 66499 6453 66508
rect 6316 66137 6356 66172
rect 6412 66212 6452 66499
rect 6315 66128 6357 66137
rect 6315 66088 6316 66128
rect 6356 66088 6357 66128
rect 6315 66079 6357 66088
rect 6316 66048 6356 66079
rect 6412 65960 6452 66172
rect 6316 65920 6452 65960
rect 6219 63860 6261 63869
rect 6219 63820 6220 63860
rect 6260 63820 6261 63860
rect 6219 63811 6261 63820
rect 6220 63029 6260 63811
rect 6219 63020 6261 63029
rect 6219 62980 6220 63020
rect 6260 62980 6261 63020
rect 6219 62971 6261 62980
rect 5876 62392 6164 62432
rect 5836 60761 5876 62392
rect 6028 62180 6068 62189
rect 5931 61592 5973 61601
rect 5931 61552 5932 61592
rect 5972 61552 5973 61592
rect 5931 61543 5973 61552
rect 5835 60752 5877 60761
rect 5835 60712 5836 60752
rect 5876 60712 5877 60752
rect 5835 60703 5877 60712
rect 5932 59912 5972 61543
rect 6028 60080 6068 62140
rect 6219 62012 6261 62021
rect 6219 61972 6220 62012
rect 6260 61972 6261 62012
rect 6219 61963 6261 61972
rect 6220 60929 6260 61963
rect 6219 60920 6261 60929
rect 6219 60880 6220 60920
rect 6260 60880 6261 60920
rect 6219 60871 6261 60880
rect 6220 60089 6260 60871
rect 6124 60080 6164 60089
rect 6028 60040 6124 60080
rect 6124 60031 6164 60040
rect 6219 60080 6261 60089
rect 6219 60040 6220 60080
rect 6260 60040 6261 60080
rect 6219 60031 6261 60040
rect 6220 59946 6260 60031
rect 5932 59872 6164 59912
rect 6028 59417 6068 59502
rect 6027 59408 6069 59417
rect 6027 59368 6028 59408
rect 6068 59368 6069 59408
rect 6027 59359 6069 59368
rect 5740 59200 6068 59240
rect 5931 58988 5973 58997
rect 5931 58948 5932 58988
rect 5972 58948 5973 58988
rect 5931 58939 5973 58948
rect 5739 58820 5781 58829
rect 5739 58780 5740 58820
rect 5780 58780 5781 58820
rect 5739 58771 5781 58780
rect 5740 58652 5780 58771
rect 5835 58736 5877 58745
rect 5835 58696 5836 58736
rect 5876 58696 5877 58736
rect 5835 58687 5877 58696
rect 5740 58603 5780 58612
rect 5836 58652 5876 58687
rect 5836 58601 5876 58612
rect 5932 56645 5972 58939
rect 5931 56636 5973 56645
rect 5931 56596 5932 56636
rect 5972 56596 5973 56636
rect 5931 56587 5973 56596
rect 5643 56384 5685 56393
rect 5643 56344 5644 56384
rect 5684 56344 5685 56384
rect 5643 56335 5685 56344
rect 5835 56384 5877 56393
rect 5835 56344 5836 56384
rect 5876 56344 5877 56384
rect 5835 56335 5877 56344
rect 5836 56250 5876 56335
rect 5932 56132 5972 56587
rect 5836 56092 5972 56132
rect 5068 54664 5396 54704
rect 5452 55336 5588 55376
rect 5740 55544 5780 55553
rect 4588 54496 4724 54536
rect 4780 54620 4820 54629
rect 4588 53948 4628 54496
rect 4780 54116 4820 54580
rect 4684 54076 4820 54116
rect 4684 54046 4724 54076
rect 4684 53997 4724 54006
rect 5068 54032 5108 54664
rect 5452 54209 5492 55336
rect 5548 54872 5588 54881
rect 5548 54629 5588 54832
rect 5740 54713 5780 55504
rect 5739 54704 5781 54713
rect 5739 54664 5740 54704
rect 5780 54664 5781 54704
rect 5739 54655 5781 54664
rect 5547 54620 5589 54629
rect 5547 54580 5548 54620
rect 5588 54580 5589 54620
rect 5547 54571 5589 54580
rect 5739 54368 5781 54377
rect 5739 54328 5740 54368
rect 5780 54328 5781 54368
rect 5739 54319 5781 54328
rect 5451 54200 5493 54209
rect 5451 54160 5452 54200
rect 5492 54160 5493 54200
rect 5451 54151 5493 54160
rect 5068 53983 5108 53992
rect 5164 54032 5204 54041
rect 4588 53908 4820 53948
rect 4395 53780 4437 53789
rect 4395 53740 4396 53780
rect 4436 53740 4437 53780
rect 4395 53731 4437 53740
rect 4683 53612 4725 53621
rect 4683 53572 4684 53612
rect 4724 53572 4725 53612
rect 4683 53563 4725 53572
rect 4300 53488 4532 53528
rect 4396 53360 4436 53369
rect 4396 53201 4436 53320
rect 4395 53192 4437 53201
rect 4395 53152 4396 53192
rect 4436 53152 4437 53192
rect 4395 53143 4437 53152
rect 4203 52772 4245 52781
rect 4203 52732 4204 52772
rect 4244 52732 4245 52772
rect 4203 52723 4245 52732
rect 4204 52520 4244 52723
rect 4299 52688 4341 52697
rect 4299 52648 4300 52688
rect 4340 52648 4341 52688
rect 4299 52639 4341 52648
rect 4204 52193 4244 52480
rect 4203 52184 4245 52193
rect 4203 52144 4204 52184
rect 4244 52144 4245 52184
rect 4203 52135 4245 52144
rect 4300 52016 4340 52639
rect 4204 51976 4340 52016
rect 4204 51848 4244 51976
rect 4204 51799 4244 51808
rect 4299 51848 4341 51857
rect 4299 51808 4300 51848
rect 4340 51808 4341 51848
rect 4299 51799 4341 51808
rect 4300 51714 4340 51799
rect 4108 51640 4244 51680
rect 3820 51556 4148 51596
rect 3688 51428 4056 51437
rect 3728 51388 3770 51428
rect 3810 51388 3852 51428
rect 3892 51388 3934 51428
rect 3974 51388 4016 51428
rect 3688 51379 4056 51388
rect 3627 51260 3669 51269
rect 4108 51260 4148 51556
rect 3627 51220 3628 51260
rect 3668 51220 3669 51260
rect 3627 51211 3669 51220
rect 3820 51220 4148 51260
rect 3532 51043 3572 51052
rect 3628 51008 3668 51211
rect 3628 50959 3668 50968
rect 3820 51008 3860 51220
rect 4011 51092 4053 51101
rect 4011 51052 4012 51092
rect 4052 51052 4053 51092
rect 4011 51043 4053 51052
rect 3820 50959 3860 50968
rect 3915 51008 3957 51017
rect 3915 50968 3916 51008
rect 3956 50968 3957 51008
rect 3915 50959 3957 50968
rect 4012 51008 4052 51043
rect 3916 50874 3956 50959
rect 4012 50957 4052 50968
rect 4107 51008 4149 51017
rect 4107 50968 4108 51008
rect 4148 50968 4149 51008
rect 4107 50959 4149 50968
rect 4108 50874 4148 50959
rect 3819 50336 3861 50345
rect 3819 50296 3820 50336
rect 3860 50296 3861 50336
rect 3819 50287 3861 50296
rect 4108 50336 4148 50345
rect 3820 50202 3860 50287
rect 4012 50093 4052 50178
rect 4011 50084 4053 50093
rect 4011 50044 4012 50084
rect 4052 50044 4053 50084
rect 4011 50035 4053 50044
rect 3688 49916 4056 49925
rect 3728 49876 3770 49916
rect 3810 49876 3852 49916
rect 3892 49876 3934 49916
rect 3974 49876 4016 49916
rect 3688 49867 4056 49876
rect 3819 49664 3861 49673
rect 3819 49624 3820 49664
rect 3860 49624 3861 49664
rect 3819 49615 3861 49624
rect 3820 49580 3860 49615
rect 3820 49529 3860 49540
rect 3915 49580 3957 49589
rect 3915 49540 3916 49580
rect 3956 49540 3957 49580
rect 3915 49531 3957 49540
rect 3380 49456 3764 49496
rect 3340 49447 3380 49456
rect 3339 48992 3381 49001
rect 3628 48992 3668 49001
rect 3339 48952 3340 48992
rect 3380 48952 3628 48992
rect 3339 48943 3381 48952
rect 3628 48943 3668 48952
rect 3724 48908 3764 49456
rect 3916 49446 3956 49531
rect 3724 48868 3956 48908
rect 3436 48824 3476 48833
rect 3244 48775 3284 48784
rect 3340 48784 3436 48824
rect 3476 48814 3572 48824
rect 3772 48814 3812 48823
rect 3476 48784 3772 48814
rect 3147 48572 3189 48581
rect 3147 48532 3148 48572
rect 3188 48532 3189 48572
rect 3147 48523 3189 48532
rect 3147 48404 3189 48413
rect 3147 48364 3148 48404
rect 3188 48364 3189 48404
rect 3147 48355 3189 48364
rect 3052 47935 3092 47944
rect 2955 47816 2997 47825
rect 2955 47776 2956 47816
rect 2996 47776 2997 47816
rect 2955 47767 2997 47776
rect 2956 47682 2996 47767
rect 2668 47104 2900 47144
rect 2956 47312 2996 47321
rect 2859 46976 2901 46985
rect 2956 46976 2996 47272
rect 2859 46936 2860 46976
rect 2900 46936 2996 46976
rect 2859 46927 2901 46936
rect 2860 46565 2900 46927
rect 2859 46556 2901 46565
rect 2859 46516 2860 46556
rect 2900 46516 2901 46556
rect 2859 46507 2901 46516
rect 2956 46472 2996 46481
rect 2668 46388 2708 46397
rect 2956 46388 2996 46432
rect 2708 46348 2996 46388
rect 3052 46472 3092 46481
rect 2668 46339 2708 46348
rect 2667 46052 2709 46061
rect 2667 46012 2668 46052
rect 2708 46012 2709 46052
rect 2667 46003 2709 46012
rect 2668 45800 2708 46003
rect 2859 45968 2901 45977
rect 2859 45928 2860 45968
rect 2900 45928 2901 45968
rect 2859 45919 2901 45928
rect 2860 45834 2900 45919
rect 2668 45751 2708 45760
rect 3052 45641 3092 46432
rect 3051 45632 3093 45641
rect 3051 45592 3052 45632
rect 3092 45592 3093 45632
rect 3051 45583 3093 45592
rect 2955 45464 2997 45473
rect 2955 45424 2956 45464
rect 2996 45424 2997 45464
rect 2955 45415 2997 45424
rect 2571 44120 2613 44129
rect 2763 44120 2805 44129
rect 2571 44080 2572 44120
rect 2612 44080 2613 44120
rect 2571 44071 2613 44080
rect 2668 44080 2764 44120
rect 2804 44080 2805 44120
rect 2668 42944 2708 44080
rect 2763 44071 2805 44080
rect 2572 42904 2708 42944
rect 2475 42440 2517 42449
rect 2475 42400 2476 42440
rect 2516 42400 2517 42440
rect 2475 42391 2517 42400
rect 2476 41945 2516 42391
rect 2475 41936 2517 41945
rect 2475 41896 2476 41936
rect 2516 41896 2517 41936
rect 2475 41887 2517 41896
rect 2476 41802 2516 41887
rect 2572 41684 2612 42904
rect 2667 42776 2709 42785
rect 2667 42736 2668 42776
rect 2708 42736 2709 42776
rect 2667 42727 2709 42736
rect 2668 42642 2708 42727
rect 2860 42524 2900 42533
rect 2572 41644 2708 41684
rect 2571 41516 2613 41525
rect 2571 41476 2572 41516
rect 2612 41476 2613 41516
rect 2571 41467 2613 41476
rect 2572 40517 2612 41467
rect 2571 40508 2613 40517
rect 2571 40468 2572 40508
rect 2612 40468 2613 40508
rect 2571 40459 2613 40468
rect 2475 40340 2517 40349
rect 2475 40300 2476 40340
rect 2516 40300 2517 40340
rect 2475 40291 2517 40300
rect 2476 39752 2516 40291
rect 2668 40097 2708 41644
rect 2763 41432 2805 41441
rect 2763 41392 2764 41432
rect 2804 41392 2805 41432
rect 2763 41383 2805 41392
rect 2667 40088 2709 40097
rect 2667 40048 2668 40088
rect 2708 40048 2709 40088
rect 2667 40039 2709 40048
rect 2668 39920 2708 39929
rect 2764 39920 2804 41383
rect 2860 41273 2900 42484
rect 2859 41264 2901 41273
rect 2859 41224 2860 41264
rect 2900 41224 2901 41264
rect 2859 41215 2901 41224
rect 2956 40340 2996 45415
rect 3148 44456 3188 48355
rect 3244 48236 3284 48245
rect 3340 48236 3380 48784
rect 3436 48775 3476 48784
rect 3532 48774 3772 48784
rect 3772 48765 3812 48774
rect 3435 48656 3477 48665
rect 3627 48656 3669 48665
rect 3435 48616 3436 48656
rect 3476 48616 3477 48656
rect 3435 48607 3477 48616
rect 3532 48616 3628 48656
rect 3668 48616 3669 48656
rect 3436 48522 3476 48607
rect 3284 48196 3380 48236
rect 3244 48187 3284 48196
rect 3339 48068 3381 48077
rect 3339 48028 3340 48068
rect 3380 48028 3381 48068
rect 3339 48019 3381 48028
rect 3340 47900 3380 48019
rect 3436 47984 3476 47993
rect 3436 47900 3476 47944
rect 3340 47860 3476 47900
rect 3243 47732 3285 47741
rect 3243 47692 3244 47732
rect 3284 47692 3285 47732
rect 3243 47683 3285 47692
rect 3244 44960 3284 47683
rect 3340 46061 3380 47860
rect 3532 47816 3572 48616
rect 3627 48607 3669 48616
rect 3916 48572 3956 48868
rect 4108 48749 4148 50296
rect 4204 49673 4244 51640
rect 4396 51596 4436 53143
rect 4300 51556 4436 51596
rect 4300 50933 4340 51556
rect 4299 50924 4341 50933
rect 4299 50884 4300 50924
rect 4340 50884 4341 50924
rect 4299 50875 4341 50884
rect 4395 50840 4437 50849
rect 4395 50800 4396 50840
rect 4436 50800 4437 50840
rect 4395 50791 4437 50800
rect 4203 49664 4245 49673
rect 4203 49624 4204 49664
rect 4244 49624 4245 49664
rect 4203 49615 4245 49624
rect 4107 48740 4149 48749
rect 4107 48700 4108 48740
rect 4148 48700 4149 48740
rect 4107 48691 4149 48700
rect 3916 48532 4148 48572
rect 3688 48404 4056 48413
rect 3728 48364 3770 48404
rect 3810 48364 3852 48404
rect 3892 48364 3934 48404
rect 3974 48364 4016 48404
rect 3688 48355 4056 48364
rect 3819 48236 3861 48245
rect 3819 48196 3820 48236
rect 3860 48196 3861 48236
rect 3819 48187 3861 48196
rect 3436 47776 3572 47816
rect 3436 46556 3476 47776
rect 3820 47060 3860 48187
rect 3436 46507 3476 46516
rect 3532 47020 3860 47060
rect 3532 46472 3572 47020
rect 3688 46892 4056 46901
rect 3728 46852 3770 46892
rect 3810 46852 3852 46892
rect 3892 46852 3934 46892
rect 3974 46852 4016 46892
rect 3688 46843 4056 46852
rect 4108 46640 4148 48532
rect 4204 48245 4244 49615
rect 4299 49496 4341 49505
rect 4299 49456 4300 49496
rect 4340 49456 4341 49496
rect 4299 49447 4341 49456
rect 4396 49496 4436 50791
rect 4396 49447 4436 49456
rect 4300 49362 4340 49447
rect 4299 49244 4341 49253
rect 4299 49204 4300 49244
rect 4340 49204 4341 49244
rect 4299 49195 4341 49204
rect 4300 48824 4340 49195
rect 4300 48775 4340 48784
rect 4492 48488 4532 53488
rect 4587 52856 4629 52865
rect 4587 52816 4588 52856
rect 4628 52816 4629 52856
rect 4587 52807 4629 52816
rect 4588 51008 4628 52807
rect 4684 51848 4724 53563
rect 4780 52016 4820 53908
rect 4876 53873 4916 53958
rect 4875 53864 4917 53873
rect 4875 53824 4876 53864
rect 4916 53824 4917 53864
rect 4875 53815 4917 53824
rect 5067 53864 5109 53873
rect 5164 53864 5204 53992
rect 5260 54032 5300 54041
rect 5740 54032 5780 54319
rect 5836 54293 5876 56092
rect 5931 55796 5973 55805
rect 5931 55756 5932 55796
rect 5972 55756 5973 55796
rect 5931 55747 5973 55756
rect 5932 55662 5972 55747
rect 6028 55460 6068 59200
rect 5932 55420 6068 55460
rect 5835 54284 5877 54293
rect 5835 54244 5836 54284
rect 5876 54244 5877 54284
rect 5835 54235 5877 54244
rect 5260 53873 5300 53992
rect 5644 53992 5740 54032
rect 5067 53824 5068 53864
rect 5108 53824 5204 53864
rect 5259 53864 5301 53873
rect 5259 53824 5260 53864
rect 5300 53824 5301 53864
rect 5067 53815 5109 53824
rect 5259 53815 5301 53824
rect 5356 53864 5396 53873
rect 4928 53696 5296 53705
rect 4968 53656 5010 53696
rect 5050 53656 5092 53696
rect 5132 53656 5174 53696
rect 5214 53656 5256 53696
rect 4928 53647 5296 53656
rect 5356 52193 5396 53824
rect 5548 53864 5588 53873
rect 5451 53696 5493 53705
rect 5451 53656 5452 53696
rect 5492 53656 5493 53696
rect 5451 53647 5493 53656
rect 5452 52865 5492 53647
rect 5548 53537 5588 53824
rect 5547 53528 5589 53537
rect 5547 53488 5548 53528
rect 5588 53488 5589 53528
rect 5547 53479 5589 53488
rect 5644 53360 5684 53992
rect 5740 53983 5780 53992
rect 5835 53696 5877 53705
rect 5835 53656 5836 53696
rect 5876 53656 5877 53696
rect 5835 53647 5877 53656
rect 5836 53528 5876 53647
rect 5836 53479 5876 53488
rect 5548 53320 5644 53360
rect 5451 52856 5493 52865
rect 5451 52816 5452 52856
rect 5492 52816 5493 52856
rect 5451 52807 5493 52816
rect 5452 52520 5492 52529
rect 5548 52520 5588 53320
rect 5644 53311 5684 53320
rect 5932 52865 5972 55420
rect 6124 54377 6164 59872
rect 6316 58736 6356 65920
rect 6508 64280 6548 66760
rect 6412 64240 6548 64280
rect 6412 63944 6452 64240
rect 6412 63895 6452 63904
rect 6508 63944 6548 63953
rect 6508 62021 6548 63904
rect 6604 63281 6644 69103
rect 6700 68228 6740 69784
rect 6795 69740 6837 69749
rect 6795 69700 6796 69740
rect 6836 69700 6837 69740
rect 6795 69691 6837 69700
rect 6796 69152 6836 69691
rect 6796 69103 6836 69112
rect 6892 69152 6932 69868
rect 6892 68573 6932 69112
rect 6988 68732 7028 73564
rect 7180 73520 7220 73529
rect 7180 73100 7220 73480
rect 7660 73109 7700 74311
rect 7659 73100 7701 73109
rect 7180 73060 7316 73100
rect 7084 73016 7124 73025
rect 7084 71765 7124 72976
rect 7179 72176 7221 72185
rect 7179 72136 7180 72176
rect 7220 72136 7221 72176
rect 7179 72127 7221 72136
rect 7083 71756 7125 71765
rect 7083 71716 7084 71756
rect 7124 71716 7125 71756
rect 7083 71707 7125 71716
rect 7180 71597 7220 72127
rect 7179 71588 7221 71597
rect 7179 71548 7180 71588
rect 7220 71548 7221 71588
rect 7179 71539 7221 71548
rect 7276 71513 7316 73060
rect 7659 73060 7660 73100
rect 7700 73060 7701 73100
rect 7659 73051 7701 73060
rect 7659 72764 7701 72773
rect 7659 72724 7660 72764
rect 7700 72724 7701 72764
rect 7659 72715 7701 72724
rect 7563 72176 7605 72185
rect 7563 72136 7564 72176
rect 7604 72136 7605 72176
rect 7563 72127 7605 72136
rect 7564 72042 7604 72127
rect 7371 72008 7413 72017
rect 7371 71968 7372 72008
rect 7412 71968 7413 72008
rect 7371 71959 7413 71968
rect 7372 71874 7412 71959
rect 7371 71756 7413 71765
rect 7371 71716 7372 71756
rect 7412 71716 7413 71756
rect 7371 71707 7413 71716
rect 7275 71504 7317 71513
rect 7275 71464 7276 71504
rect 7316 71464 7317 71504
rect 7275 71455 7317 71464
rect 7084 71420 7124 71429
rect 7084 70664 7124 71380
rect 7180 71420 7220 71429
rect 7180 71261 7220 71380
rect 7179 71252 7221 71261
rect 7179 71212 7180 71252
rect 7220 71212 7221 71252
rect 7179 71203 7221 71212
rect 7275 70832 7317 70841
rect 7275 70792 7276 70832
rect 7316 70792 7317 70832
rect 7275 70783 7317 70792
rect 7276 70673 7316 70783
rect 7275 70664 7317 70673
rect 7084 70624 7220 70664
rect 7084 70496 7124 70505
rect 7084 69245 7124 70456
rect 7083 69236 7125 69245
rect 7083 69196 7084 69236
rect 7124 69196 7125 69236
rect 7083 69187 7125 69196
rect 7180 69161 7220 70624
rect 7275 70624 7276 70664
rect 7316 70624 7317 70664
rect 7275 70615 7317 70624
rect 7276 70530 7316 70615
rect 7372 69824 7412 71707
rect 7660 71672 7700 72715
rect 7564 71632 7700 71672
rect 7467 70580 7509 70589
rect 7467 70540 7468 70580
rect 7508 70540 7509 70580
rect 7467 70531 7509 70540
rect 7468 69992 7508 70531
rect 7468 69943 7508 69952
rect 7372 69784 7508 69824
rect 7179 69152 7221 69161
rect 7179 69112 7180 69152
rect 7220 69112 7221 69152
rect 7179 69103 7221 69112
rect 7276 69152 7316 69161
rect 6988 68692 7220 68732
rect 6891 68564 6933 68573
rect 6891 68524 6892 68564
rect 6932 68524 6933 68564
rect 6891 68515 6933 68524
rect 6796 68405 6836 68490
rect 6795 68396 6837 68405
rect 6795 68356 6796 68396
rect 6836 68356 6837 68396
rect 6795 68347 6837 68356
rect 6892 68396 6932 68405
rect 6892 68228 6932 68356
rect 6700 68188 6932 68228
rect 6699 68060 6741 68069
rect 6699 68020 6700 68060
rect 6740 68020 6741 68060
rect 6699 68011 6741 68020
rect 6603 63272 6645 63281
rect 6603 63232 6604 63272
rect 6644 63232 6645 63272
rect 6603 63223 6645 63232
rect 6507 62012 6549 62021
rect 6507 61972 6508 62012
rect 6548 61972 6549 62012
rect 6507 61963 6549 61972
rect 6411 61760 6453 61769
rect 6604 61760 6644 63223
rect 6700 61769 6740 68011
rect 6795 67892 6837 67901
rect 6795 67852 6796 67892
rect 6836 67852 6837 67892
rect 6795 67843 6837 67852
rect 6796 64205 6836 67843
rect 6892 66473 6932 68188
rect 6891 66464 6933 66473
rect 6891 66424 6892 66464
rect 6932 66424 6933 66464
rect 6891 66415 6933 66424
rect 6892 66128 6932 66137
rect 6892 65297 6932 66088
rect 7083 65456 7125 65465
rect 7083 65416 7084 65456
rect 7124 65416 7125 65456
rect 7083 65407 7125 65416
rect 6891 65288 6933 65297
rect 6891 65248 6892 65288
rect 6932 65248 6933 65288
rect 6891 65239 6933 65248
rect 7084 64709 7124 65407
rect 7083 64700 7125 64709
rect 7083 64660 7084 64700
rect 7124 64660 7125 64700
rect 7083 64651 7125 64660
rect 7084 64616 7124 64651
rect 6891 64364 6933 64373
rect 6891 64324 6892 64364
rect 6932 64324 6933 64364
rect 6891 64315 6933 64324
rect 6795 64196 6837 64205
rect 6795 64156 6796 64196
rect 6836 64156 6837 64196
rect 6795 64147 6837 64156
rect 6892 63860 6932 64315
rect 6988 63869 7028 63954
rect 6796 63820 6892 63860
rect 6796 62357 6836 63820
rect 6892 63811 6932 63820
rect 6987 63860 7029 63869
rect 6987 63820 6988 63860
rect 7028 63820 7029 63860
rect 6987 63811 7029 63820
rect 7084 63692 7124 64576
rect 6892 63652 7124 63692
rect 6892 63104 6932 63652
rect 6795 62348 6837 62357
rect 6795 62308 6796 62348
rect 6836 62308 6837 62348
rect 6795 62299 6837 62308
rect 6411 61720 6412 61760
rect 6452 61720 6453 61760
rect 6411 61711 6453 61720
rect 6508 61720 6644 61760
rect 6699 61760 6741 61769
rect 6699 61720 6700 61760
rect 6740 61720 6741 61760
rect 6412 59333 6452 61711
rect 6508 60845 6548 61720
rect 6699 61711 6741 61720
rect 6603 61592 6645 61601
rect 6603 61552 6604 61592
rect 6644 61552 6645 61592
rect 6603 61543 6645 61552
rect 6604 61458 6644 61543
rect 6795 61424 6837 61433
rect 6795 61384 6796 61424
rect 6836 61384 6837 61424
rect 6795 61375 6837 61384
rect 6796 61290 6836 61375
rect 6892 61172 6932 63064
rect 7083 63020 7125 63029
rect 7083 62980 7084 63020
rect 7124 62980 7125 63020
rect 7083 62971 7125 62980
rect 7084 62886 7124 62971
rect 7180 61769 7220 68692
rect 7276 68405 7316 69112
rect 7371 69152 7413 69161
rect 7371 69112 7372 69152
rect 7412 69112 7413 69152
rect 7371 69103 7413 69112
rect 7372 69018 7412 69103
rect 7372 68480 7412 68489
rect 7275 68396 7317 68405
rect 7275 68356 7276 68396
rect 7316 68356 7317 68396
rect 7275 68347 7317 68356
rect 7372 67985 7412 68440
rect 7468 68069 7508 69784
rect 7564 69572 7604 71632
rect 7659 71504 7701 71513
rect 7659 71464 7660 71504
rect 7700 71464 7701 71504
rect 7659 71455 7701 71464
rect 7660 70589 7700 71455
rect 7659 70580 7701 70589
rect 7659 70540 7660 70580
rect 7700 70540 7701 70580
rect 7659 70531 7701 70540
rect 7756 70001 7796 75403
rect 7852 73949 7892 83887
rect 7948 83777 7988 85936
rect 8140 84029 8180 85936
rect 8139 84020 8181 84029
rect 8139 83980 8140 84020
rect 8180 83980 8181 84020
rect 8139 83971 8181 83980
rect 7947 83768 7989 83777
rect 7947 83728 7948 83768
rect 7988 83728 7989 83768
rect 7947 83719 7989 83728
rect 8332 83768 8372 85936
rect 8524 85457 8564 85936
rect 8523 85448 8565 85457
rect 8523 85408 8524 85448
rect 8564 85408 8565 85448
rect 8523 85399 8565 85408
rect 8523 84692 8565 84701
rect 8523 84652 8524 84692
rect 8564 84652 8565 84692
rect 8523 84643 8565 84652
rect 8427 84440 8469 84449
rect 8427 84400 8428 84440
rect 8468 84400 8469 84440
rect 8427 84391 8469 84400
rect 8332 83719 8372 83728
rect 7948 83516 7988 83525
rect 7948 83189 7988 83476
rect 8139 83516 8181 83525
rect 8139 83476 8140 83516
rect 8180 83476 8181 83516
rect 8139 83467 8181 83476
rect 8140 83382 8180 83467
rect 7947 83180 7989 83189
rect 7947 83140 7948 83180
rect 7988 83140 7989 83180
rect 7947 83131 7989 83140
rect 8428 78392 8468 84391
rect 8524 83768 8564 84643
rect 8716 83945 8756 85936
rect 8715 83936 8757 83945
rect 8715 83896 8716 83936
rect 8756 83896 8757 83936
rect 8715 83887 8757 83896
rect 8524 83719 8564 83728
rect 8715 83516 8757 83525
rect 8715 83476 8716 83516
rect 8756 83476 8757 83516
rect 8715 83467 8757 83476
rect 8716 83382 8756 83467
rect 8619 83348 8661 83357
rect 8619 83308 8620 83348
rect 8660 83308 8661 83348
rect 8619 83299 8661 83308
rect 8523 83264 8565 83273
rect 8523 83224 8524 83264
rect 8564 83224 8565 83264
rect 8523 83215 8565 83224
rect 8428 77720 8468 78352
rect 8428 76889 8468 77680
rect 8427 76880 8469 76889
rect 8427 76840 8428 76880
rect 8468 76840 8469 76880
rect 8427 76831 8469 76840
rect 8524 76721 8564 83215
rect 7948 76712 7988 76721
rect 7948 76049 7988 76672
rect 8428 76712 8468 76721
rect 8140 76628 8180 76637
rect 8428 76628 8468 76672
rect 8523 76712 8565 76721
rect 8523 76672 8524 76712
rect 8564 76672 8565 76712
rect 8523 76663 8565 76672
rect 8180 76588 8468 76628
rect 8140 76579 8180 76588
rect 8524 76578 8564 76663
rect 8427 76208 8469 76217
rect 8427 76168 8428 76208
rect 8468 76168 8469 76208
rect 8427 76159 8469 76168
rect 7947 76040 7989 76049
rect 7947 76000 7948 76040
rect 7988 76000 7989 76040
rect 7947 75991 7989 76000
rect 7948 75200 7988 75991
rect 8140 75788 8180 75797
rect 8180 75748 8372 75788
rect 8140 75739 8180 75748
rect 8332 75200 8372 75748
rect 8428 75368 8468 76159
rect 8428 75319 8468 75328
rect 8620 75200 8660 83299
rect 8812 77552 8852 77563
rect 8812 77477 8852 77512
rect 8811 77468 8853 77477
rect 8811 77428 8812 77468
rect 8852 77428 8853 77468
rect 8811 77419 8853 77428
rect 8908 77048 8948 85936
rect 9003 80492 9045 80501
rect 9003 80452 9004 80492
rect 9044 80452 9045 80492
rect 9003 80443 9045 80452
rect 8812 77008 8948 77048
rect 8715 76628 8757 76637
rect 8715 76588 8716 76628
rect 8756 76588 8757 76628
rect 8715 76579 8757 76588
rect 8716 76040 8756 76579
rect 8716 75991 8756 76000
rect 7988 75160 8084 75200
rect 8332 75160 8564 75200
rect 8620 75160 8756 75200
rect 7948 75151 7988 75160
rect 7947 74948 7989 74957
rect 7947 74908 7948 74948
rect 7988 74908 7989 74948
rect 7947 74899 7989 74908
rect 7851 73940 7893 73949
rect 7851 73900 7852 73940
rect 7892 73900 7893 73940
rect 7851 73891 7893 73900
rect 7851 73100 7893 73109
rect 7851 73060 7852 73100
rect 7892 73060 7893 73100
rect 7851 73051 7893 73060
rect 7852 72941 7892 73051
rect 7851 72932 7893 72941
rect 7851 72892 7852 72932
rect 7892 72892 7893 72932
rect 7851 72883 7893 72892
rect 7755 69992 7797 70001
rect 7755 69952 7756 69992
rect 7796 69952 7797 69992
rect 7755 69943 7797 69952
rect 7660 69740 7700 69749
rect 7700 69700 7796 69740
rect 7660 69691 7700 69700
rect 7564 69532 7700 69572
rect 7563 68480 7605 68489
rect 7563 68440 7564 68480
rect 7604 68440 7605 68480
rect 7563 68431 7605 68440
rect 7467 68060 7509 68069
rect 7467 68020 7468 68060
rect 7508 68020 7509 68060
rect 7467 68011 7509 68020
rect 7371 67976 7413 67985
rect 7371 67936 7372 67976
rect 7412 67936 7413 67976
rect 7371 67927 7413 67936
rect 7467 67640 7509 67649
rect 7467 67600 7468 67640
rect 7508 67600 7509 67640
rect 7467 67591 7509 67600
rect 7468 67506 7508 67591
rect 7371 67472 7413 67481
rect 7371 67432 7372 67472
rect 7412 67432 7413 67472
rect 7371 67423 7413 67432
rect 7372 66142 7412 67423
rect 7467 67388 7509 67397
rect 7467 67348 7468 67388
rect 7508 67348 7509 67388
rect 7467 67339 7509 67348
rect 7468 67220 7508 67339
rect 7564 67304 7604 68431
rect 7660 67649 7700 69532
rect 7756 68984 7796 69700
rect 7851 69320 7893 69329
rect 7851 69280 7852 69320
rect 7892 69280 7893 69320
rect 7851 69271 7893 69280
rect 7852 69152 7892 69271
rect 7852 69103 7892 69112
rect 7756 68944 7892 68984
rect 7852 68475 7892 68944
rect 7852 68426 7892 68435
rect 7851 68228 7893 68237
rect 7851 68188 7852 68228
rect 7892 68188 7893 68228
rect 7851 68179 7893 68188
rect 7659 67640 7701 67649
rect 7659 67600 7660 67640
rect 7700 67600 7701 67640
rect 7659 67591 7701 67600
rect 7852 67640 7892 68179
rect 7948 67901 7988 74899
rect 8044 74528 8084 75160
rect 8139 75032 8181 75041
rect 8139 74992 8140 75032
rect 8180 74992 8181 75032
rect 8139 74983 8181 74992
rect 8332 75032 8372 75041
rect 8140 74898 8180 74983
rect 8332 74612 8372 74992
rect 8044 74369 8084 74488
rect 8140 74572 8372 74612
rect 8043 74360 8085 74369
rect 8043 74320 8044 74360
rect 8084 74320 8085 74360
rect 8043 74311 8085 74320
rect 8140 73100 8180 74572
rect 8524 74528 8564 75160
rect 8524 74479 8564 74488
rect 8619 74528 8661 74537
rect 8619 74488 8620 74528
rect 8660 74488 8661 74528
rect 8619 74479 8661 74488
rect 8620 74394 8660 74479
rect 8236 74276 8276 74285
rect 8276 74236 8564 74276
rect 8236 74227 8276 74236
rect 8524 73688 8564 74236
rect 8716 73697 8756 75160
rect 8812 74957 8852 77008
rect 8907 76880 8949 76889
rect 8907 76840 8908 76880
rect 8948 76840 8949 76880
rect 9004 76880 9044 80443
rect 9100 79241 9140 85936
rect 9292 83945 9332 85936
rect 9291 83936 9333 83945
rect 9291 83896 9292 83936
rect 9332 83896 9333 83936
rect 9291 83887 9333 83896
rect 9291 83516 9333 83525
rect 9291 83476 9292 83516
rect 9332 83476 9333 83516
rect 9291 83467 9333 83476
rect 9195 83264 9237 83273
rect 9195 83224 9196 83264
rect 9236 83224 9237 83264
rect 9195 83215 9237 83224
rect 9099 79232 9141 79241
rect 9099 79192 9100 79232
rect 9140 79192 9141 79232
rect 9099 79183 9141 79192
rect 9100 79064 9140 79073
rect 9100 78905 9140 79024
rect 9099 78896 9141 78905
rect 9099 78856 9100 78896
rect 9140 78856 9141 78896
rect 9099 78847 9141 78856
rect 9196 77561 9236 83215
rect 9195 77552 9237 77561
rect 9195 77512 9196 77552
rect 9236 77512 9237 77552
rect 9195 77503 9237 77512
rect 9195 76880 9237 76889
rect 9004 76840 9140 76880
rect 8907 76831 8949 76840
rect 8908 76796 8948 76831
rect 8908 76217 8948 76756
rect 9003 76712 9045 76721
rect 9003 76672 9004 76712
rect 9044 76672 9045 76712
rect 9003 76663 9045 76672
rect 9004 76578 9044 76663
rect 8907 76208 8949 76217
rect 8907 76168 8908 76208
rect 8948 76168 8949 76208
rect 8907 76159 8949 76168
rect 8907 75368 8949 75377
rect 8907 75328 8908 75368
rect 8948 75328 8949 75368
rect 8907 75319 8949 75328
rect 8811 74948 8853 74957
rect 8811 74908 8812 74948
rect 8852 74908 8853 74948
rect 8811 74899 8853 74908
rect 8908 73865 8948 75319
rect 9100 74780 9140 76840
rect 9195 76840 9196 76880
rect 9236 76840 9237 76880
rect 9195 76831 9237 76840
rect 9196 75377 9236 76831
rect 9195 75368 9237 75377
rect 9195 75328 9196 75368
rect 9236 75328 9237 75368
rect 9195 75319 9237 75328
rect 9196 75200 9236 75209
rect 9196 74957 9236 75160
rect 9195 74948 9237 74957
rect 9195 74908 9196 74948
rect 9236 74908 9237 74948
rect 9195 74899 9237 74908
rect 9100 74740 9236 74780
rect 9003 74528 9045 74537
rect 9003 74488 9004 74528
rect 9044 74488 9045 74528
rect 9003 74479 9045 74488
rect 9004 74394 9044 74479
rect 9099 74444 9141 74453
rect 9099 74404 9100 74444
rect 9140 74404 9141 74444
rect 9099 74395 9141 74404
rect 9100 74310 9140 74395
rect 8907 73856 8949 73865
rect 8907 73816 8908 73856
rect 8948 73816 8949 73856
rect 8907 73807 8949 73816
rect 9003 73772 9045 73781
rect 9003 73732 9004 73772
rect 9044 73732 9045 73772
rect 9003 73723 9045 73732
rect 8524 73639 8564 73648
rect 8620 73688 8660 73697
rect 8715 73688 8757 73697
rect 8660 73648 8716 73688
rect 8756 73648 8757 73688
rect 8620 73639 8660 73648
rect 8715 73639 8757 73648
rect 8235 73604 8277 73613
rect 8235 73564 8236 73604
rect 8276 73564 8277 73604
rect 8235 73555 8277 73564
rect 8044 73060 8180 73100
rect 8044 68732 8084 73060
rect 8139 72008 8181 72017
rect 8139 71968 8140 72008
rect 8180 71968 8181 72008
rect 8139 71959 8181 71968
rect 8140 71499 8180 71959
rect 8140 71450 8180 71459
rect 8236 70757 8276 73555
rect 8716 73554 8756 73639
rect 8524 73100 8564 73140
rect 9004 73100 9044 73723
rect 9099 73688 9141 73697
rect 9099 73648 9100 73688
rect 9140 73648 9141 73688
rect 9099 73639 9141 73648
rect 9100 73554 9140 73639
rect 8524 73025 8564 73060
rect 8908 73060 9044 73100
rect 8523 73016 8565 73025
rect 8332 72974 8372 72983
rect 8331 72934 8332 72941
rect 8523 72976 8524 73016
rect 8564 72976 8565 73016
rect 8523 72967 8565 72976
rect 8716 73016 8756 73025
rect 8524 72965 8564 72967
rect 8372 72934 8373 72941
rect 8331 72932 8373 72934
rect 8331 72892 8332 72932
rect 8372 72892 8373 72932
rect 8716 72932 8756 72976
rect 8811 72932 8853 72941
rect 8716 72892 8812 72932
rect 8852 72892 8853 72932
rect 8331 72883 8373 72892
rect 8811 72883 8853 72892
rect 8332 72764 8372 72883
rect 8332 72724 8468 72764
rect 8331 72596 8373 72605
rect 8331 72556 8332 72596
rect 8372 72556 8373 72596
rect 8331 72547 8373 72556
rect 8332 71672 8372 72547
rect 8428 72092 8468 72724
rect 8812 72176 8852 72185
rect 8812 72092 8852 72136
rect 8428 72052 8852 72092
rect 8427 71756 8469 71765
rect 8427 71716 8428 71756
rect 8468 71716 8469 71756
rect 8427 71707 8469 71716
rect 8332 71623 8372 71632
rect 8235 70748 8277 70757
rect 8235 70708 8236 70748
rect 8276 70708 8277 70748
rect 8235 70699 8277 70708
rect 8428 70328 8468 71707
rect 8523 71420 8565 71429
rect 8523 71380 8524 71420
rect 8564 71380 8565 71420
rect 8523 71371 8565 71380
rect 8524 71286 8564 71371
rect 8524 70664 8564 70673
rect 8620 70664 8660 72052
rect 8715 71252 8757 71261
rect 8715 71212 8716 71252
rect 8756 71212 8757 71252
rect 8715 71203 8757 71212
rect 8716 71118 8756 71203
rect 8715 70916 8757 70925
rect 8715 70876 8716 70916
rect 8756 70876 8757 70916
rect 8715 70867 8757 70876
rect 8716 70782 8756 70867
rect 8908 70664 8948 73060
rect 9004 72008 9044 72017
rect 9004 71504 9044 71968
rect 9004 71455 9044 71464
rect 9099 71504 9141 71513
rect 9099 71464 9100 71504
rect 9140 71464 9141 71504
rect 9099 71455 9141 71464
rect 9100 71370 9140 71455
rect 9003 70748 9045 70757
rect 9003 70708 9004 70748
rect 9044 70708 9045 70748
rect 9003 70699 9045 70708
rect 8564 70624 8660 70664
rect 8812 70624 8948 70664
rect 8524 70615 8564 70624
rect 8428 70288 8564 70328
rect 8235 70076 8277 70085
rect 8235 70036 8236 70076
rect 8276 70036 8277 70076
rect 8235 70027 8277 70036
rect 8044 68692 8180 68732
rect 8043 68564 8085 68573
rect 8043 68524 8044 68564
rect 8084 68524 8085 68564
rect 8043 68515 8085 68524
rect 8044 68430 8084 68515
rect 7947 67892 7989 67901
rect 7947 67852 7948 67892
rect 7988 67852 7989 67892
rect 7947 67843 7989 67852
rect 7852 67591 7892 67600
rect 8043 67640 8085 67649
rect 8043 67600 8044 67640
rect 8084 67600 8085 67640
rect 8043 67591 8085 67600
rect 7660 67472 7700 67481
rect 7660 67388 7700 67432
rect 7660 67348 7988 67388
rect 7564 67264 7700 67304
rect 7468 67180 7604 67220
rect 7372 66093 7412 66102
rect 7564 66044 7604 67180
rect 7564 65995 7604 66004
rect 7468 65456 7508 65465
rect 7276 65204 7316 65213
rect 7276 64625 7316 65164
rect 7275 64616 7317 64625
rect 7275 64576 7276 64616
rect 7316 64576 7317 64616
rect 7275 64567 7317 64576
rect 7275 64448 7317 64457
rect 7275 64408 7276 64448
rect 7316 64408 7317 64448
rect 7275 64399 7317 64408
rect 7276 64314 7316 64399
rect 7468 64121 7508 65416
rect 7564 64616 7604 64627
rect 7564 64541 7604 64576
rect 7660 64616 7700 67264
rect 7948 66968 7988 67348
rect 7948 66919 7988 66928
rect 8044 66968 8084 67591
rect 8044 66919 8084 66928
rect 8140 66800 8180 68692
rect 8236 68489 8276 70027
rect 8427 69992 8469 70001
rect 8427 69952 8428 69992
rect 8468 69952 8469 69992
rect 8427 69943 8469 69952
rect 8428 69858 8468 69943
rect 8331 69236 8373 69245
rect 8331 69196 8332 69236
rect 8372 69196 8373 69236
rect 8331 69187 8373 69196
rect 8332 69166 8372 69187
rect 8332 69101 8372 69126
rect 8524 69068 8564 70288
rect 8524 69019 8564 69028
rect 8235 68480 8277 68489
rect 8235 68440 8236 68480
rect 8276 68440 8277 68480
rect 8235 68431 8277 68440
rect 8619 68396 8661 68405
rect 8619 68356 8620 68396
rect 8660 68356 8661 68396
rect 8619 68347 8661 68356
rect 8523 66968 8565 66977
rect 8523 66928 8524 66968
rect 8564 66928 8565 66968
rect 8523 66919 8565 66928
rect 8427 66884 8469 66893
rect 8427 66844 8428 66884
rect 8468 66844 8469 66884
rect 8427 66835 8469 66844
rect 7563 64532 7605 64541
rect 7563 64492 7564 64532
rect 7604 64492 7605 64532
rect 7563 64483 7605 64492
rect 7660 64289 7700 64576
rect 7852 66760 8180 66800
rect 7659 64280 7701 64289
rect 7659 64240 7660 64280
rect 7700 64240 7701 64280
rect 7659 64231 7701 64240
rect 7275 64112 7317 64121
rect 7275 64072 7276 64112
rect 7316 64072 7317 64112
rect 7275 64063 7317 64072
rect 7467 64112 7509 64121
rect 7467 64072 7468 64112
rect 7508 64072 7509 64112
rect 7467 64063 7509 64072
rect 7179 61760 7221 61769
rect 7179 61720 7180 61760
rect 7220 61720 7221 61760
rect 7179 61711 7221 61720
rect 7180 61592 7220 61601
rect 7083 61508 7125 61517
rect 7180 61508 7220 61552
rect 7083 61468 7084 61508
rect 7124 61468 7220 61508
rect 7083 61459 7125 61468
rect 7179 61340 7221 61349
rect 7179 61300 7180 61340
rect 7220 61300 7221 61340
rect 7179 61291 7221 61300
rect 6796 61132 6932 61172
rect 6700 60920 6740 60929
rect 6507 60836 6549 60845
rect 6507 60796 6508 60836
rect 6548 60796 6549 60836
rect 6507 60787 6549 60796
rect 6700 60761 6740 60880
rect 6699 60752 6741 60761
rect 6699 60712 6700 60752
rect 6740 60712 6741 60752
rect 6699 60703 6741 60712
rect 6699 60164 6741 60173
rect 6699 60124 6700 60164
rect 6740 60124 6741 60164
rect 6699 60115 6741 60124
rect 6603 60080 6645 60089
rect 6603 60040 6604 60080
rect 6644 60040 6645 60080
rect 6603 60031 6645 60040
rect 6604 59946 6644 60031
rect 6700 60030 6740 60115
rect 6699 59912 6741 59921
rect 6699 59872 6700 59912
rect 6740 59872 6741 59912
rect 6699 59863 6741 59872
rect 6411 59324 6453 59333
rect 6411 59284 6412 59324
rect 6452 59284 6453 59324
rect 6411 59275 6453 59284
rect 6316 58696 6452 58736
rect 6315 58568 6357 58577
rect 6315 58528 6316 58568
rect 6356 58528 6357 58568
rect 6315 58519 6357 58528
rect 6316 58434 6356 58519
rect 6219 58400 6261 58409
rect 6219 58360 6220 58400
rect 6260 58360 6261 58400
rect 6219 58351 6261 58360
rect 6220 57485 6260 58351
rect 6219 57476 6261 57485
rect 6219 57436 6220 57476
rect 6260 57436 6261 57476
rect 6219 57427 6261 57436
rect 6219 55796 6261 55805
rect 6219 55756 6220 55796
rect 6260 55756 6261 55796
rect 6219 55747 6261 55756
rect 6220 55544 6260 55747
rect 6220 55495 6260 55504
rect 6316 55544 6356 55553
rect 6316 54377 6356 55504
rect 6412 55460 6452 58696
rect 6700 58493 6740 59863
rect 6796 59249 6836 61132
rect 7180 60920 7220 61291
rect 7276 61097 7316 64063
rect 7467 63944 7509 63953
rect 7467 63904 7468 63944
rect 7508 63904 7509 63944
rect 7467 63895 7509 63904
rect 7468 63810 7508 63895
rect 7371 63104 7413 63113
rect 7371 63064 7372 63104
rect 7412 63064 7413 63104
rect 7371 63055 7413 63064
rect 7275 61088 7317 61097
rect 7275 61048 7276 61088
rect 7316 61048 7317 61088
rect 7275 61039 7317 61048
rect 7180 60871 7220 60880
rect 7275 60920 7317 60929
rect 7275 60880 7276 60920
rect 7316 60880 7317 60920
rect 7275 60871 7317 60880
rect 6987 60836 7029 60845
rect 6987 60796 6988 60836
rect 7028 60796 7029 60836
rect 6987 60787 7029 60796
rect 6891 60668 6933 60677
rect 6891 60628 6892 60668
rect 6932 60628 6933 60668
rect 6891 60619 6933 60628
rect 6892 60534 6932 60619
rect 6988 60416 7028 60787
rect 7276 60786 7316 60871
rect 6892 60376 7028 60416
rect 6795 59240 6837 59249
rect 6795 59200 6796 59240
rect 6836 59200 6837 59240
rect 6795 59191 6837 59200
rect 6796 58573 6836 58582
rect 6699 58484 6741 58493
rect 6699 58444 6700 58484
rect 6740 58444 6741 58484
rect 6699 58435 6741 58444
rect 6796 58064 6836 58533
rect 6796 58015 6836 58024
rect 6603 57980 6645 57989
rect 6603 57940 6604 57980
rect 6644 57940 6645 57980
rect 6603 57931 6645 57940
rect 6604 57896 6644 57931
rect 6604 57845 6644 57856
rect 6795 56216 6837 56225
rect 6795 56176 6796 56216
rect 6836 56176 6837 56216
rect 6795 56167 6837 56176
rect 6796 55721 6836 56167
rect 6795 55712 6837 55721
rect 6795 55672 6796 55712
rect 6836 55672 6837 55712
rect 6795 55663 6837 55672
rect 6603 55628 6645 55637
rect 6603 55588 6604 55628
rect 6644 55588 6645 55628
rect 6603 55579 6645 55588
rect 6604 55460 6644 55579
rect 6700 55553 6740 55638
rect 6699 55544 6741 55553
rect 6699 55504 6700 55544
rect 6740 55504 6741 55544
rect 6699 55495 6741 55504
rect 6796 55544 6836 55553
rect 6412 55420 6644 55460
rect 6507 55208 6549 55217
rect 6507 55168 6508 55208
rect 6548 55168 6549 55208
rect 6507 55159 6549 55168
rect 6411 55040 6453 55049
rect 6411 55000 6412 55040
rect 6452 55000 6453 55040
rect 6411 54991 6453 55000
rect 6123 54368 6165 54377
rect 6123 54328 6124 54368
rect 6164 54328 6165 54368
rect 6123 54319 6165 54328
rect 6315 54368 6357 54377
rect 6315 54328 6316 54368
rect 6356 54328 6357 54368
rect 6315 54319 6357 54328
rect 6316 54032 6356 54319
rect 6220 53992 6356 54032
rect 6220 53621 6260 53992
rect 6315 53864 6357 53873
rect 6315 53824 6316 53864
rect 6356 53824 6357 53864
rect 6315 53815 6357 53824
rect 6219 53612 6261 53621
rect 6219 53572 6220 53612
rect 6260 53572 6261 53612
rect 6219 53563 6261 53572
rect 6028 53444 6068 53453
rect 5931 52856 5973 52865
rect 5931 52816 5932 52856
rect 5972 52816 5973 52856
rect 5931 52807 5973 52816
rect 6028 52533 6068 53404
rect 6219 53444 6261 53453
rect 6219 53404 6220 53444
rect 6260 53404 6261 53444
rect 6219 53395 6261 53404
rect 5492 52480 5588 52520
rect 5452 52471 5492 52480
rect 4928 52184 5296 52193
rect 4968 52144 5010 52184
rect 5050 52144 5092 52184
rect 5132 52144 5174 52184
rect 5214 52144 5256 52184
rect 4928 52135 5296 52144
rect 5355 52184 5397 52193
rect 5355 52144 5356 52184
rect 5396 52144 5397 52184
rect 5355 52135 5397 52144
rect 5451 52016 5493 52025
rect 4780 51976 4916 52016
rect 4684 51799 4724 51808
rect 4780 51848 4820 51857
rect 4780 51101 4820 51808
rect 4876 51353 4916 51976
rect 5451 51976 5452 52016
rect 5492 51976 5493 52016
rect 5451 51967 5493 51976
rect 5355 51932 5397 51941
rect 5355 51892 5356 51932
rect 5396 51892 5397 51932
rect 5355 51883 5397 51892
rect 5356 51848 5396 51883
rect 5452 51882 5492 51967
rect 5356 51797 5396 51808
rect 4875 51344 4917 51353
rect 4875 51304 4876 51344
rect 4916 51304 4917 51344
rect 4875 51295 4917 51304
rect 4779 51092 4821 51101
rect 4779 51052 4780 51092
rect 4820 51052 4821 51092
rect 4779 51043 4821 51052
rect 4684 51008 4724 51017
rect 4588 50968 4684 51008
rect 4684 50765 4724 50968
rect 4683 50756 4725 50765
rect 4683 50716 4684 50756
rect 4724 50716 4725 50756
rect 4683 50707 4725 50716
rect 4928 50672 5296 50681
rect 4968 50632 5010 50672
rect 5050 50632 5092 50672
rect 5132 50632 5174 50672
rect 5214 50632 5256 50672
rect 4928 50623 5296 50632
rect 4588 50336 4628 50345
rect 4588 50009 4628 50296
rect 4587 50000 4629 50009
rect 4587 49960 4588 50000
rect 4628 49960 4629 50000
rect 4587 49951 4629 49960
rect 5451 49664 5493 49673
rect 4588 49624 4916 49664
rect 4588 48581 4628 49624
rect 4780 49496 4820 49505
rect 4683 49328 4725 49337
rect 4683 49288 4684 49328
rect 4724 49288 4725 49328
rect 4683 49279 4725 49288
rect 4684 49194 4724 49279
rect 4780 49169 4820 49456
rect 4876 49496 4916 49624
rect 5451 49624 5452 49664
rect 5492 49624 5493 49664
rect 5451 49615 5493 49624
rect 4876 49447 4916 49456
rect 4972 49496 5012 49507
rect 4972 49421 5012 49456
rect 4971 49412 5013 49421
rect 4971 49372 4972 49412
rect 5012 49372 5013 49412
rect 4971 49363 5013 49372
rect 4779 49160 4821 49169
rect 4779 49120 4780 49160
rect 4820 49120 4821 49160
rect 4779 49111 4821 49120
rect 4928 49160 5296 49169
rect 4968 49120 5010 49160
rect 5050 49120 5092 49160
rect 5132 49120 5174 49160
rect 5214 49120 5256 49160
rect 4928 49111 5296 49120
rect 4875 48992 4917 49001
rect 4875 48952 4876 48992
rect 4916 48952 4917 48992
rect 4875 48943 4917 48952
rect 4779 48908 4821 48917
rect 4779 48868 4780 48908
rect 4820 48868 4821 48908
rect 4779 48859 4821 48868
rect 4780 48824 4820 48859
rect 4780 48773 4820 48784
rect 4876 48824 4916 48943
rect 5452 48917 5492 49615
rect 5451 48908 5493 48917
rect 5451 48868 5452 48908
rect 5492 48868 5493 48908
rect 5451 48859 5493 48868
rect 4876 48775 4916 48784
rect 5259 48824 5301 48833
rect 5259 48784 5260 48824
rect 5300 48784 5301 48824
rect 5259 48775 5301 48784
rect 5356 48824 5396 48833
rect 5260 48690 5300 48775
rect 5356 48581 5396 48784
rect 4587 48572 4629 48581
rect 4587 48532 4588 48572
rect 4628 48532 4629 48572
rect 4587 48523 4629 48532
rect 5355 48572 5397 48581
rect 5355 48532 5356 48572
rect 5396 48532 5397 48572
rect 5355 48523 5397 48532
rect 4300 48448 4532 48488
rect 4203 48236 4245 48245
rect 4203 48196 4204 48236
rect 4244 48196 4245 48236
rect 4203 48187 4245 48196
rect 4203 47900 4245 47909
rect 4203 47860 4204 47900
rect 4244 47860 4245 47900
rect 4203 47851 4245 47860
rect 4204 47312 4244 47851
rect 4204 47263 4244 47272
rect 4300 46640 4340 48448
rect 5355 48404 5397 48413
rect 5355 48364 5356 48404
rect 5396 48364 5397 48404
rect 5355 48355 5397 48364
rect 4683 47984 4725 47993
rect 4683 47944 4684 47984
rect 4724 47944 4725 47984
rect 4683 47935 4725 47944
rect 5356 47984 5396 48355
rect 5548 48077 5588 52480
rect 5836 52520 5876 52529
rect 6028 52484 6068 52493
rect 6220 53355 6260 53395
rect 6220 52520 6260 53315
rect 5644 52436 5684 52445
rect 5836 52436 5876 52480
rect 6220 52471 6260 52480
rect 5684 52396 5876 52436
rect 6316 52436 6356 53815
rect 6412 53789 6452 54991
rect 6508 54200 6548 55159
rect 6604 54284 6644 55420
rect 6796 55049 6836 55504
rect 6795 55040 6837 55049
rect 6795 55000 6796 55040
rect 6836 55000 6837 55040
rect 6795 54991 6837 55000
rect 6796 54872 6836 54881
rect 6796 54713 6836 54832
rect 6795 54704 6837 54713
rect 6795 54664 6796 54704
rect 6836 54664 6837 54704
rect 6795 54655 6837 54664
rect 6604 54244 6740 54284
rect 6508 54160 6644 54200
rect 6604 53957 6644 54160
rect 6603 53948 6645 53957
rect 6603 53908 6604 53948
rect 6644 53908 6645 53948
rect 6603 53899 6645 53908
rect 6411 53780 6453 53789
rect 6411 53740 6412 53780
rect 6452 53740 6453 53780
rect 6411 53731 6453 53740
rect 6412 52697 6452 53731
rect 6507 53696 6549 53705
rect 6507 53656 6508 53696
rect 6548 53656 6549 53696
rect 6507 53647 6549 53656
rect 6508 53369 6548 53647
rect 6507 53360 6549 53369
rect 6507 53320 6508 53360
rect 6548 53320 6549 53360
rect 6507 53311 6549 53320
rect 6411 52688 6453 52697
rect 6411 52648 6412 52688
rect 6452 52648 6453 52688
rect 6411 52639 6453 52648
rect 5644 52387 5684 52396
rect 5643 52184 5685 52193
rect 5643 52144 5644 52184
rect 5684 52144 5685 52184
rect 5643 52135 5685 52144
rect 5644 51848 5684 52135
rect 5644 51799 5684 51808
rect 5740 51848 5780 52396
rect 6316 52387 6356 52396
rect 6412 52520 6452 52529
rect 5740 51799 5780 51808
rect 5932 52352 5972 52361
rect 5932 51848 5972 52312
rect 6412 52025 6452 52480
rect 6508 52520 6548 53311
rect 6604 52697 6644 53899
rect 6700 53873 6740 54244
rect 6795 54200 6837 54209
rect 6795 54160 6796 54200
rect 6836 54160 6837 54200
rect 6795 54151 6837 54160
rect 6699 53864 6741 53873
rect 6699 53824 6700 53864
rect 6740 53824 6741 53864
rect 6699 53815 6741 53824
rect 6700 53360 6740 53815
rect 6700 53311 6740 53320
rect 6603 52688 6645 52697
rect 6603 52648 6604 52688
rect 6644 52648 6645 52688
rect 6603 52639 6645 52648
rect 6508 52471 6548 52480
rect 6603 52436 6645 52445
rect 6603 52396 6604 52436
rect 6644 52396 6645 52436
rect 6603 52387 6645 52396
rect 6411 52016 6453 52025
rect 5932 51799 5972 51808
rect 6028 51976 6260 52016
rect 5931 51680 5973 51689
rect 5931 51640 5932 51680
rect 5972 51640 5973 51680
rect 5931 51631 5973 51640
rect 5643 51596 5685 51605
rect 5643 51556 5644 51596
rect 5684 51556 5685 51596
rect 5643 51547 5685 51556
rect 5644 49496 5684 51547
rect 5932 51546 5972 51631
rect 5931 51344 5973 51353
rect 5931 51304 5932 51344
rect 5972 51304 5973 51344
rect 5931 51295 5973 51304
rect 5932 51008 5972 51295
rect 5932 50959 5972 50968
rect 6028 50345 6068 51976
rect 6123 51848 6165 51857
rect 6123 51808 6124 51848
rect 6164 51808 6165 51848
rect 6123 51799 6165 51808
rect 6220 51848 6260 51976
rect 6411 51976 6412 52016
rect 6452 51976 6453 52016
rect 6411 51967 6453 51976
rect 6604 52016 6644 52387
rect 6604 51967 6644 51976
rect 6700 52352 6740 52361
rect 6796 52352 6836 54151
rect 6892 52940 6932 60376
rect 7180 60080 7220 60089
rect 7180 59921 7220 60040
rect 7179 59912 7221 59921
rect 7179 59872 7180 59912
rect 7220 59872 7221 59912
rect 7179 59863 7221 59872
rect 6987 59408 7029 59417
rect 7276 59408 7316 59417
rect 6987 59368 6988 59408
rect 7028 59368 7029 59408
rect 6987 59359 7029 59368
rect 7180 59368 7276 59408
rect 6988 58484 7028 59359
rect 7180 59249 7220 59368
rect 7276 59359 7316 59368
rect 7179 59240 7221 59249
rect 7372 59240 7412 63055
rect 7563 63020 7605 63029
rect 7563 62980 7564 63020
rect 7604 62980 7605 63020
rect 7563 62971 7605 62980
rect 7564 62432 7604 62971
rect 7564 62383 7604 62392
rect 7659 62432 7701 62441
rect 7659 62392 7660 62432
rect 7700 62392 7701 62432
rect 7659 62383 7701 62392
rect 7467 62348 7509 62357
rect 7467 62308 7468 62348
rect 7508 62308 7509 62348
rect 7467 62299 7509 62308
rect 7468 60089 7508 62299
rect 7660 62298 7700 62383
rect 7563 62096 7605 62105
rect 7563 62056 7564 62096
rect 7604 62056 7605 62096
rect 7563 62047 7605 62056
rect 7467 60080 7509 60089
rect 7467 60040 7468 60080
rect 7508 60040 7509 60080
rect 7467 60031 7509 60040
rect 7564 59921 7604 62047
rect 7659 61676 7701 61685
rect 7659 61636 7660 61676
rect 7700 61636 7701 61676
rect 7659 61627 7701 61636
rect 7660 61517 7700 61627
rect 7659 61508 7701 61517
rect 7659 61468 7660 61508
rect 7700 61468 7701 61508
rect 7659 61459 7701 61468
rect 7660 60845 7700 60930
rect 7659 60836 7701 60845
rect 7659 60796 7660 60836
rect 7700 60796 7701 60836
rect 7659 60787 7701 60796
rect 7756 60836 7796 60845
rect 7659 60668 7701 60677
rect 7659 60628 7660 60668
rect 7700 60628 7701 60668
rect 7659 60619 7701 60628
rect 7660 60094 7700 60619
rect 7756 60173 7796 60796
rect 7755 60164 7797 60173
rect 7755 60124 7756 60164
rect 7796 60124 7797 60164
rect 7755 60115 7797 60124
rect 7660 60045 7700 60054
rect 7563 59912 7605 59921
rect 7563 59872 7564 59912
rect 7604 59872 7605 59912
rect 7563 59863 7605 59872
rect 7179 59200 7180 59240
rect 7220 59200 7221 59240
rect 7179 59191 7221 59200
rect 7276 59200 7412 59240
rect 7468 59240 7508 59249
rect 7508 59200 7604 59240
rect 6988 58435 7028 58444
rect 7179 58484 7221 58493
rect 7179 58444 7180 58484
rect 7220 58444 7221 58484
rect 7179 58435 7221 58444
rect 7180 57812 7220 58435
rect 7084 57772 7220 57812
rect 6988 57056 7028 57065
rect 6988 56729 7028 57016
rect 6987 56720 7029 56729
rect 6987 56680 6988 56720
rect 7028 56680 7029 56720
rect 6987 56671 7029 56680
rect 7084 56645 7124 57772
rect 7180 57317 7220 57402
rect 7179 57308 7221 57317
rect 7179 57268 7180 57308
rect 7220 57268 7221 57308
rect 7179 57259 7221 57268
rect 7179 57056 7221 57065
rect 7179 57016 7180 57056
rect 7220 57016 7221 57056
rect 7179 57007 7221 57016
rect 7180 56922 7220 57007
rect 7276 56804 7316 59200
rect 7468 59191 7508 59200
rect 7564 58568 7604 59200
rect 7659 58736 7701 58745
rect 7659 58696 7660 58736
rect 7700 58696 7701 58736
rect 7659 58687 7701 58696
rect 7564 58519 7604 58528
rect 7660 58568 7700 58687
rect 7660 58519 7700 58528
rect 7371 58400 7413 58409
rect 7371 58360 7372 58400
rect 7412 58360 7413 58400
rect 7371 58351 7413 58360
rect 7180 56764 7316 56804
rect 7372 57056 7412 58351
rect 7564 57989 7604 58020
rect 7563 57980 7605 57989
rect 7563 57940 7564 57980
rect 7604 57940 7605 57980
rect 7563 57931 7605 57940
rect 7564 57896 7604 57931
rect 7564 57401 7604 57856
rect 7563 57392 7605 57401
rect 7563 57352 7564 57392
rect 7604 57352 7605 57392
rect 7563 57343 7605 57352
rect 7083 56636 7125 56645
rect 7083 56596 7084 56636
rect 7124 56596 7125 56636
rect 7083 56587 7125 56596
rect 6987 56552 7029 56561
rect 6987 56512 6988 56552
rect 7028 56512 7029 56552
rect 6987 56503 7029 56512
rect 6988 55217 7028 56503
rect 7084 56384 7124 56393
rect 6987 55208 7029 55217
rect 6987 55168 6988 55208
rect 7028 55168 7029 55208
rect 6987 55159 7029 55168
rect 6987 55040 7029 55049
rect 6987 55000 6988 55040
rect 7028 55000 7029 55040
rect 6987 54991 7029 55000
rect 6988 54906 7028 54991
rect 7084 54713 7124 56344
rect 7180 55217 7220 56764
rect 7275 56636 7317 56645
rect 7275 56596 7276 56636
rect 7316 56596 7317 56636
rect 7275 56587 7317 56596
rect 7276 56384 7316 56587
rect 7372 56561 7412 57016
rect 7468 57056 7508 57065
rect 7371 56552 7413 56561
rect 7371 56512 7372 56552
rect 7412 56512 7413 56552
rect 7371 56503 7413 56512
rect 7468 56384 7508 57016
rect 7564 57056 7604 57065
rect 7564 56552 7604 57016
rect 7659 56888 7701 56897
rect 7659 56848 7660 56888
rect 7700 56848 7701 56888
rect 7659 56839 7701 56848
rect 7660 56754 7700 56839
rect 7564 56512 7700 56552
rect 7564 56384 7604 56393
rect 7276 56344 7412 56384
rect 7275 56216 7317 56225
rect 7275 56176 7276 56216
rect 7316 56176 7317 56216
rect 7275 56167 7317 56176
rect 7276 56082 7316 56167
rect 7276 55553 7316 55638
rect 7275 55544 7317 55553
rect 7275 55504 7276 55544
rect 7316 55504 7317 55544
rect 7275 55495 7317 55504
rect 7179 55208 7221 55217
rect 7179 55168 7180 55208
rect 7220 55168 7221 55208
rect 7179 55159 7221 55168
rect 7372 55124 7412 56344
rect 7468 56344 7564 56384
rect 7468 55553 7508 56344
rect 7564 56335 7604 56344
rect 7563 56216 7605 56225
rect 7563 56176 7564 56216
rect 7604 56176 7605 56216
rect 7563 56167 7605 56176
rect 7467 55544 7509 55553
rect 7467 55504 7468 55544
rect 7508 55504 7509 55544
rect 7467 55495 7509 55504
rect 7276 55084 7412 55124
rect 7083 54704 7125 54713
rect 7083 54664 7084 54704
rect 7124 54664 7125 54704
rect 7083 54655 7125 54664
rect 7179 54200 7221 54209
rect 7179 54160 7180 54200
rect 7220 54160 7221 54200
rect 7276 54200 7316 55084
rect 7468 55049 7508 55495
rect 7467 55040 7509 55049
rect 7467 55000 7468 55040
rect 7508 55000 7509 55040
rect 7467 54991 7509 55000
rect 7372 54872 7412 54881
rect 7372 54461 7412 54832
rect 7468 54872 7508 54991
rect 7564 54965 7604 56167
rect 7660 55040 7700 56512
rect 7756 56132 7796 60115
rect 7852 60089 7892 66760
rect 8428 66750 8468 66835
rect 8524 66834 8564 66919
rect 8139 66632 8181 66641
rect 8620 66632 8660 68347
rect 8715 67976 8757 67985
rect 8715 67936 8716 67976
rect 8756 67936 8757 67976
rect 8715 67927 8757 67936
rect 8716 66809 8756 67927
rect 8715 66800 8757 66809
rect 8715 66760 8716 66800
rect 8756 66760 8757 66800
rect 8715 66751 8757 66760
rect 8139 66592 8140 66632
rect 8180 66592 8181 66632
rect 8139 66583 8181 66592
rect 8428 66592 8660 66632
rect 8140 64700 8180 66583
rect 8044 64616 8084 64625
rect 7947 64448 7989 64457
rect 7947 64408 7948 64448
rect 7988 64408 7989 64448
rect 7947 64399 7989 64408
rect 7948 63939 7988 64399
rect 8044 64373 8084 64576
rect 8043 64364 8085 64373
rect 8043 64324 8044 64364
rect 8084 64324 8085 64364
rect 8043 64315 8085 64324
rect 8140 64196 8180 64660
rect 7948 63890 7988 63899
rect 8044 64156 8180 64196
rect 8044 63692 8084 64156
rect 8140 64028 8180 64037
rect 8140 63869 8180 63988
rect 8331 64028 8373 64037
rect 8331 63988 8332 64028
rect 8372 63988 8373 64028
rect 8331 63979 8373 63988
rect 8139 63860 8181 63869
rect 8139 63820 8140 63860
rect 8180 63820 8181 63860
rect 8139 63811 8181 63820
rect 8044 63652 8180 63692
rect 7947 62516 7989 62525
rect 7947 62476 7948 62516
rect 7988 62476 7989 62516
rect 7947 62467 7989 62476
rect 7851 60080 7893 60089
rect 7851 60040 7852 60080
rect 7892 60040 7893 60080
rect 7851 60031 7893 60040
rect 7851 59912 7893 59921
rect 7851 59872 7852 59912
rect 7892 59872 7893 59912
rect 7851 59863 7893 59872
rect 7852 59778 7892 59863
rect 7851 59576 7893 59585
rect 7851 59536 7852 59576
rect 7892 59536 7893 59576
rect 7851 59527 7893 59536
rect 7852 59408 7892 59527
rect 7852 59333 7892 59368
rect 7851 59324 7893 59333
rect 7851 59284 7852 59324
rect 7892 59284 7893 59324
rect 7851 59275 7893 59284
rect 7948 57989 7988 62467
rect 8043 62348 8085 62357
rect 8043 62308 8044 62348
rect 8084 62308 8085 62348
rect 8043 62299 8085 62308
rect 8140 62348 8180 63652
rect 8235 62432 8277 62441
rect 8235 62392 8236 62432
rect 8276 62392 8277 62432
rect 8235 62383 8277 62392
rect 8044 62214 8084 62299
rect 8043 61928 8085 61937
rect 8043 61888 8044 61928
rect 8084 61888 8085 61928
rect 8043 61879 8085 61888
rect 8044 61433 8084 61879
rect 8043 61424 8085 61433
rect 8043 61384 8044 61424
rect 8084 61384 8085 61424
rect 8043 61375 8085 61384
rect 8044 58577 8084 58662
rect 8043 58568 8085 58577
rect 8043 58528 8044 58568
rect 8084 58528 8085 58568
rect 8043 58519 8085 58528
rect 8140 58568 8180 62308
rect 8236 60920 8276 62383
rect 8236 59165 8276 60880
rect 8235 59156 8277 59165
rect 8235 59116 8236 59156
rect 8276 59116 8277 59156
rect 8235 59107 8277 59116
rect 8140 58493 8180 58528
rect 8139 58484 8181 58493
rect 8139 58444 8140 58484
rect 8180 58444 8181 58484
rect 8139 58435 8181 58444
rect 7947 57980 7989 57989
rect 7947 57940 7948 57980
rect 7988 57940 7989 57980
rect 7947 57931 7989 57940
rect 7852 57056 7892 57065
rect 7852 56561 7892 57016
rect 8139 56888 8181 56897
rect 8139 56848 8140 56888
rect 8180 56848 8181 56888
rect 8139 56839 8181 56848
rect 7947 56804 7989 56813
rect 7947 56764 7948 56804
rect 7988 56764 7989 56804
rect 7947 56755 7989 56764
rect 7851 56552 7893 56561
rect 7851 56512 7852 56552
rect 7892 56512 7893 56552
rect 7851 56503 7893 56512
rect 7948 56468 7988 56755
rect 7948 56419 7988 56428
rect 7851 56384 7893 56393
rect 7851 56344 7852 56384
rect 7892 56344 7893 56384
rect 7851 56335 7893 56344
rect 7852 56250 7892 56335
rect 7947 56132 7989 56141
rect 7756 56092 7892 56132
rect 7756 55553 7796 55639
rect 7755 55549 7797 55553
rect 7755 55504 7756 55549
rect 7796 55504 7797 55549
rect 7755 55495 7797 55504
rect 7755 55376 7797 55385
rect 7755 55336 7756 55376
rect 7796 55336 7797 55376
rect 7755 55327 7797 55336
rect 7660 54991 7700 55000
rect 7563 54956 7605 54965
rect 7563 54916 7564 54956
rect 7604 54916 7605 54956
rect 7563 54907 7605 54916
rect 7468 54823 7508 54832
rect 7371 54452 7413 54461
rect 7371 54412 7372 54452
rect 7412 54412 7508 54452
rect 7371 54403 7413 54412
rect 7276 54160 7412 54200
rect 7179 54151 7221 54160
rect 6988 54032 7028 54041
rect 7028 53992 7124 54032
rect 6988 53983 7028 53992
rect 6892 52900 7028 52940
rect 6892 52529 6932 52614
rect 6891 52520 6933 52529
rect 6891 52480 6892 52520
rect 6932 52480 6933 52520
rect 6891 52471 6933 52480
rect 6796 52312 6932 52352
rect 6220 51799 6260 51808
rect 6412 51848 6452 51857
rect 6700 51848 6740 52312
rect 6452 51808 6548 51848
rect 6700 51838 6788 51848
rect 6700 51808 6748 51838
rect 6412 51799 6452 51808
rect 6124 51714 6164 51799
rect 6219 51680 6261 51689
rect 6219 51640 6220 51680
rect 6260 51640 6261 51680
rect 6219 51631 6261 51640
rect 6124 51260 6164 51269
rect 6220 51260 6260 51631
rect 6164 51220 6260 51260
rect 6412 51596 6452 51605
rect 6124 51211 6164 51220
rect 6316 51008 6356 51019
rect 6316 50933 6356 50968
rect 6315 50924 6357 50933
rect 6315 50884 6316 50924
rect 6356 50884 6357 50924
rect 6315 50875 6357 50884
rect 6412 50504 6452 51556
rect 6316 50464 6452 50504
rect 5836 50336 5876 50345
rect 5739 50084 5781 50093
rect 5739 50044 5740 50084
rect 5780 50044 5781 50084
rect 5739 50035 5781 50044
rect 5547 48068 5589 48077
rect 5547 48028 5548 48068
rect 5588 48028 5589 48068
rect 5644 48068 5684 49456
rect 5740 48824 5780 50035
rect 5836 49925 5876 50296
rect 6027 50336 6069 50345
rect 6027 50296 6028 50336
rect 6068 50296 6069 50336
rect 6027 50287 6069 50296
rect 6028 50093 6068 50287
rect 6027 50084 6069 50093
rect 6027 50044 6028 50084
rect 6068 50044 6069 50084
rect 6027 50035 6069 50044
rect 6028 49950 6068 50035
rect 5835 49916 5877 49925
rect 5835 49876 5836 49916
rect 5876 49876 5877 49916
rect 5835 49867 5877 49876
rect 6123 49916 6165 49925
rect 6123 49876 6124 49916
rect 6164 49876 6165 49916
rect 6123 49867 6165 49876
rect 5835 49496 5877 49505
rect 5835 49456 5836 49496
rect 5876 49456 5877 49496
rect 5835 49447 5877 49456
rect 5740 48775 5780 48784
rect 5836 48824 5876 49447
rect 6124 49421 6164 49867
rect 6316 49505 6356 50464
rect 6508 50429 6548 51808
rect 6748 51789 6788 51798
rect 6892 51680 6932 52312
rect 6700 51640 6932 51680
rect 6507 50420 6549 50429
rect 6507 50380 6508 50420
rect 6548 50380 6549 50420
rect 6507 50371 6549 50380
rect 6412 50336 6452 50345
rect 6315 49496 6357 49505
rect 6315 49456 6316 49496
rect 6356 49456 6357 49496
rect 6315 49447 6357 49456
rect 6123 49412 6165 49421
rect 6123 49372 6124 49412
rect 6164 49372 6165 49412
rect 6123 49363 6165 49372
rect 5876 48784 5972 48824
rect 5836 48775 5876 48784
rect 5644 48028 5780 48068
rect 5547 48019 5589 48028
rect 5356 47935 5396 47944
rect 4684 47850 4724 47935
rect 5740 47732 5780 48028
rect 5452 47692 5780 47732
rect 4928 47648 5296 47657
rect 4968 47608 5010 47648
rect 5050 47608 5092 47648
rect 5132 47608 5174 47648
rect 5214 47608 5256 47648
rect 4928 47599 5296 47608
rect 4588 47321 4628 47406
rect 4587 47312 4629 47321
rect 4587 47272 4588 47312
rect 4628 47272 4629 47312
rect 4587 47263 4629 47272
rect 4876 47312 4916 47321
rect 3532 46313 3572 46432
rect 4012 46600 4148 46640
rect 4204 46600 4340 46640
rect 4396 47060 4436 47069
rect 4396 46640 4436 47020
rect 4588 47060 4628 47069
rect 4396 46600 4532 46640
rect 4012 46472 4052 46600
rect 4012 46423 4052 46432
rect 3531 46304 3573 46313
rect 3531 46264 3532 46304
rect 3572 46264 3573 46304
rect 3531 46255 3573 46264
rect 4011 46304 4053 46313
rect 4011 46264 4012 46304
rect 4052 46264 4053 46304
rect 4011 46255 4053 46264
rect 3339 46052 3381 46061
rect 3339 46012 3340 46052
rect 3380 46012 3381 46052
rect 3339 46003 3381 46012
rect 3339 45884 3381 45893
rect 3339 45844 3340 45884
rect 3380 45844 3381 45884
rect 3339 45835 3381 45844
rect 3340 45750 3380 45835
rect 4012 45800 4052 46255
rect 3532 45786 3572 45795
rect 4012 45751 4052 45760
rect 3436 45212 3476 45221
rect 3532 45212 3572 45746
rect 4204 45473 4244 46600
rect 4492 46486 4532 46600
rect 4492 46437 4532 46446
rect 4588 45884 4628 47020
rect 4876 46640 4916 47272
rect 5452 46649 5492 47692
rect 5643 47564 5685 47573
rect 5643 47524 5644 47564
rect 5684 47524 5685 47564
rect 5643 47515 5685 47524
rect 5547 47228 5589 47237
rect 5547 47188 5548 47228
rect 5588 47188 5589 47228
rect 5547 47179 5589 47188
rect 5451 46640 5493 46649
rect 4876 46600 5108 46640
rect 4971 46472 5013 46481
rect 4971 46432 4972 46472
rect 5012 46432 5013 46472
rect 4971 46423 5013 46432
rect 5068 46472 5108 46600
rect 5451 46600 5452 46640
rect 5492 46600 5493 46640
rect 5451 46591 5493 46600
rect 4972 46338 5012 46423
rect 5068 46397 5108 46432
rect 5164 46472 5204 46481
rect 5067 46388 5109 46397
rect 5067 46348 5068 46388
rect 5108 46348 5109 46388
rect 5067 46339 5109 46348
rect 4683 46304 4725 46313
rect 4876 46304 4916 46313
rect 4683 46264 4684 46304
rect 4724 46264 4725 46304
rect 4683 46255 4725 46264
rect 4780 46264 4876 46304
rect 5164 46304 5204 46432
rect 5164 46264 5396 46304
rect 4684 46170 4724 46255
rect 4396 45844 4628 45884
rect 4683 45884 4725 45893
rect 4683 45844 4684 45884
rect 4724 45844 4725 45884
rect 4203 45464 4245 45473
rect 4203 45424 4204 45464
rect 4244 45424 4245 45464
rect 4203 45415 4245 45424
rect 3688 45380 4056 45389
rect 3728 45340 3770 45380
rect 3810 45340 3852 45380
rect 3892 45340 3934 45380
rect 3974 45340 4016 45380
rect 3688 45331 4056 45340
rect 4396 45305 4436 45844
rect 4683 45835 4725 45844
rect 4492 45716 4532 45725
rect 4492 45557 4532 45676
rect 4587 45716 4629 45725
rect 4587 45676 4588 45716
rect 4628 45676 4629 45716
rect 4587 45667 4629 45676
rect 4588 45582 4628 45667
rect 4491 45548 4533 45557
rect 4491 45508 4492 45548
rect 4532 45508 4533 45548
rect 4491 45499 4533 45508
rect 4395 45296 4437 45305
rect 4395 45256 4396 45296
rect 4436 45256 4437 45296
rect 4395 45247 4437 45256
rect 3915 45212 3957 45221
rect 3476 45172 3764 45212
rect 3436 45163 3476 45172
rect 3244 44633 3284 44920
rect 3724 44960 3764 45172
rect 3915 45172 3916 45212
rect 3956 45172 3957 45212
rect 3915 45163 3957 45172
rect 3724 44911 3764 44920
rect 3916 44960 3956 45163
rect 4012 45128 4052 45137
rect 4396 45128 4436 45137
rect 4052 45088 4396 45128
rect 4012 45079 4052 45088
rect 4396 45079 4436 45088
rect 3916 44911 3956 44920
rect 4011 44960 4053 44969
rect 4011 44920 4012 44960
rect 4052 44920 4053 44960
rect 4011 44911 4053 44920
rect 4396 44952 4436 44961
rect 4012 44826 4052 44911
rect 4299 44876 4341 44885
rect 4299 44836 4300 44876
rect 4340 44836 4341 44876
rect 4299 44827 4341 44836
rect 4203 44792 4245 44801
rect 4203 44752 4204 44792
rect 4244 44752 4245 44792
rect 4203 44743 4245 44752
rect 4204 44658 4244 44743
rect 3243 44624 3285 44633
rect 3243 44584 3244 44624
rect 3284 44584 3285 44624
rect 3243 44575 3285 44584
rect 3052 44416 3188 44456
rect 3339 44456 3381 44465
rect 3339 44416 3340 44456
rect 3380 44416 3381 44456
rect 3052 43457 3092 44416
rect 3339 44407 3381 44416
rect 3148 44288 3188 44297
rect 3148 44129 3188 44248
rect 3147 44120 3189 44129
rect 3147 44080 3148 44120
rect 3188 44080 3189 44120
rect 3147 44071 3189 44080
rect 3051 43448 3093 43457
rect 3051 43408 3052 43448
rect 3092 43408 3093 43448
rect 3051 43399 3093 43408
rect 3340 43448 3380 44407
rect 4107 44288 4149 44297
rect 4107 44248 4108 44288
rect 4148 44248 4149 44288
rect 4107 44239 4149 44248
rect 3688 43868 4056 43877
rect 3728 43828 3770 43868
rect 3810 43828 3852 43868
rect 3892 43828 3934 43868
rect 3974 43828 4016 43868
rect 3688 43819 4056 43828
rect 3628 43448 3668 43457
rect 3340 43408 3628 43448
rect 3052 42953 3092 43399
rect 3051 42944 3093 42953
rect 3051 42904 3052 42944
rect 3092 42904 3093 42944
rect 3051 42895 3093 42904
rect 3148 42776 3188 42785
rect 3051 42104 3093 42113
rect 3051 42064 3052 42104
rect 3092 42064 3093 42104
rect 3051 42055 3093 42064
rect 3052 41264 3092 42055
rect 3148 41441 3188 42736
rect 3243 42776 3285 42785
rect 3243 42736 3244 42776
rect 3284 42736 3285 42776
rect 3243 42727 3285 42736
rect 3244 42642 3284 42727
rect 3243 41936 3285 41945
rect 3243 41896 3244 41936
rect 3284 41896 3285 41936
rect 3243 41887 3285 41896
rect 3147 41432 3189 41441
rect 3147 41392 3148 41432
rect 3188 41392 3189 41432
rect 3147 41383 3189 41392
rect 3244 41432 3284 41887
rect 3244 41383 3284 41392
rect 3340 41264 3380 43408
rect 3628 43399 3668 43408
rect 3628 42692 3668 42703
rect 3628 42617 3668 42652
rect 3723 42692 3765 42701
rect 3723 42652 3724 42692
rect 3764 42652 3765 42692
rect 3723 42643 3765 42652
rect 3627 42608 3669 42617
rect 3627 42568 3628 42608
rect 3668 42568 3669 42608
rect 3627 42559 3669 42568
rect 3724 42558 3764 42643
rect 3688 42356 4056 42365
rect 3728 42316 3770 42356
rect 3810 42316 3852 42356
rect 3892 42316 3934 42356
rect 3974 42316 4016 42356
rect 3688 42307 4056 42316
rect 3915 42188 3957 42197
rect 4108 42188 4148 44239
rect 4300 42944 4340 44827
rect 4396 44792 4436 44912
rect 4684 44960 4724 45835
rect 4780 44969 4820 46264
rect 4876 46255 4916 46264
rect 4928 46136 5296 46145
rect 4968 46096 5010 46136
rect 5050 46096 5092 46136
rect 5132 46096 5174 46136
rect 5214 46096 5256 46136
rect 4928 46087 5296 46096
rect 5356 46061 5396 46264
rect 5355 46052 5397 46061
rect 5355 46012 5356 46052
rect 5396 46012 5397 46052
rect 5355 46003 5397 46012
rect 5067 45968 5109 45977
rect 5067 45928 5068 45968
rect 5108 45928 5109 45968
rect 5067 45919 5109 45928
rect 4972 45800 5012 45809
rect 4972 45641 5012 45760
rect 5068 45800 5108 45919
rect 5068 45751 5108 45760
rect 4971 45632 5013 45641
rect 4971 45592 4972 45632
rect 5012 45592 5013 45632
rect 4971 45583 5013 45592
rect 4972 45389 5012 45583
rect 4971 45380 5013 45389
rect 4971 45340 4972 45380
rect 5012 45340 5013 45380
rect 4971 45331 5013 45340
rect 4971 45128 5013 45137
rect 4971 45088 4972 45128
rect 5012 45088 5013 45128
rect 4971 45079 5013 45088
rect 4684 44911 4724 44920
rect 4779 44960 4821 44969
rect 4779 44920 4780 44960
rect 4820 44920 4821 44960
rect 4779 44911 4821 44920
rect 4972 44960 5012 45079
rect 4972 44911 5012 44920
rect 5548 44960 5588 47179
rect 4876 44792 4916 44801
rect 4396 44752 4876 44792
rect 4876 44743 4916 44752
rect 4395 44624 4437 44633
rect 4395 44584 4396 44624
rect 4436 44584 4437 44624
rect 4395 44575 4437 44584
rect 4928 44624 5296 44633
rect 4968 44584 5010 44624
rect 5050 44584 5092 44624
rect 5132 44584 5174 44624
rect 5214 44584 5256 44624
rect 4928 44575 5296 44584
rect 4396 44288 4436 44575
rect 4587 44456 4629 44465
rect 4587 44416 4588 44456
rect 4628 44416 4629 44456
rect 4587 44407 4629 44416
rect 4588 44322 4628 44407
rect 4875 44288 4917 44297
rect 4436 44248 4532 44288
rect 4396 44239 4436 44248
rect 4300 42904 4436 42944
rect 4203 42860 4245 42869
rect 4203 42820 4204 42860
rect 4244 42820 4245 42860
rect 4203 42811 4245 42820
rect 4204 42776 4244 42811
rect 4204 42725 4244 42736
rect 4299 42776 4341 42785
rect 4299 42736 4300 42776
rect 4340 42736 4341 42776
rect 4299 42727 4341 42736
rect 3915 42148 3916 42188
rect 3956 42148 3957 42188
rect 3915 42139 3957 42148
rect 4012 42148 4148 42188
rect 3723 42104 3765 42113
rect 3723 42064 3724 42104
rect 3764 42064 3765 42104
rect 3723 42055 3765 42064
rect 3724 41936 3764 42055
rect 3916 42054 3956 42139
rect 3724 41887 3764 41896
rect 3819 41600 3861 41609
rect 3819 41560 3820 41600
rect 3860 41560 3861 41600
rect 3819 41551 3861 41560
rect 3092 41224 3188 41264
rect 3052 41215 3092 41224
rect 3148 40424 3188 41224
rect 3148 40349 3188 40384
rect 3244 41224 3380 41264
rect 3723 41264 3765 41273
rect 3723 41224 3724 41264
rect 3764 41224 3765 41264
rect 3147 40340 3189 40349
rect 2956 40300 3092 40340
rect 2708 39880 2804 39920
rect 2668 39871 2708 39880
rect 2380 39712 2476 39752
rect 2283 39668 2325 39677
rect 2283 39628 2284 39668
rect 2324 39628 2325 39668
rect 2283 39619 2325 39628
rect 2187 32192 2229 32201
rect 2187 32152 2188 32192
rect 2228 32152 2229 32192
rect 2187 32143 2229 32152
rect 2092 31564 2228 31604
rect 2091 31352 2133 31361
rect 2091 31312 2092 31352
rect 2132 31312 2133 31352
rect 2091 31303 2133 31312
rect 1995 30092 2037 30101
rect 1995 30052 1996 30092
rect 2036 30052 2037 30092
rect 1995 30043 2037 30052
rect 1995 29924 2037 29933
rect 1995 29884 1996 29924
rect 2036 29884 2037 29924
rect 1995 29875 2037 29884
rect 1996 29840 2036 29875
rect 1996 29789 2036 29800
rect 1708 26984 1748 27616
rect 1708 26935 1748 26944
rect 1804 27952 1940 27992
rect 1996 29336 2036 29345
rect 1516 26767 1556 26776
rect 1228 26682 1268 26767
rect 1708 26648 1748 26657
rect 1419 26312 1461 26321
rect 1419 26272 1420 26312
rect 1460 26272 1461 26312
rect 1419 26263 1461 26272
rect 1708 26312 1748 26608
rect 1227 26228 1269 26237
rect 1227 26188 1228 26228
rect 1268 26188 1269 26228
rect 1227 26179 1269 26188
rect 1228 26094 1268 26179
rect 1323 26144 1365 26153
rect 1323 26104 1324 26144
rect 1364 26104 1365 26144
rect 1323 26095 1365 26104
rect 1420 26144 1460 26263
rect 1420 26095 1460 26104
rect 1516 26144 1556 26153
rect 1324 26010 1364 26095
rect 1516 25901 1556 26104
rect 1515 25892 1557 25901
rect 1515 25852 1516 25892
rect 1556 25852 1557 25892
rect 1515 25843 1557 25852
rect 1708 25472 1748 26272
rect 1228 25304 1268 25313
rect 1131 24716 1173 24725
rect 1131 24676 1132 24716
rect 1172 24676 1173 24716
rect 1131 24667 1173 24676
rect 1132 20768 1172 24667
rect 1228 24641 1268 25264
rect 1420 25304 1460 25313
rect 1323 25136 1365 25145
rect 1323 25096 1324 25136
rect 1364 25096 1365 25136
rect 1323 25087 1365 25096
rect 1324 25002 1364 25087
rect 1420 24977 1460 25264
rect 1516 25304 1556 25313
rect 1419 24968 1461 24977
rect 1419 24928 1420 24968
rect 1460 24928 1461 24968
rect 1419 24919 1461 24928
rect 1420 24800 1460 24809
rect 1516 24800 1556 25264
rect 1611 25304 1653 25313
rect 1611 25264 1612 25304
rect 1652 25264 1653 25304
rect 1611 25255 1653 25264
rect 1460 24760 1556 24800
rect 1420 24751 1460 24760
rect 1227 24632 1269 24641
rect 1227 24592 1228 24632
rect 1268 24592 1269 24632
rect 1227 24583 1269 24592
rect 1324 24632 1364 24641
rect 1324 23213 1364 24592
rect 1516 24632 1556 24641
rect 1612 24632 1652 25255
rect 1556 24592 1652 24632
rect 1708 24800 1748 25432
rect 1516 24583 1556 24592
rect 1708 24464 1748 24760
rect 1516 24424 1748 24464
rect 1516 23960 1556 24424
rect 1804 24296 1844 27952
rect 1996 27917 2036 29296
rect 1995 27908 2037 27917
rect 1995 27868 1996 27908
rect 2036 27868 2037 27908
rect 1995 27859 2037 27868
rect 1995 26816 2037 26825
rect 1995 26776 1996 26816
rect 2036 26776 2037 26816
rect 1995 26767 2037 26776
rect 1996 26682 2036 26767
rect 1995 26396 2037 26405
rect 1995 26356 1996 26396
rect 2036 26356 2037 26396
rect 1995 26347 2037 26356
rect 1899 26228 1941 26237
rect 1899 26188 1900 26228
rect 1940 26188 1941 26228
rect 1899 26179 1941 26188
rect 1900 25304 1940 26179
rect 1996 26144 2036 26347
rect 1996 26095 2036 26104
rect 1996 25556 2036 25565
rect 2092 25556 2132 31303
rect 2188 29849 2228 31564
rect 2187 29840 2229 29849
rect 2187 29800 2188 29840
rect 2228 29800 2229 29840
rect 2187 29791 2229 29800
rect 2284 29345 2324 39619
rect 2380 38240 2420 39712
rect 2476 39703 2516 39712
rect 2667 39752 2709 39761
rect 2667 39712 2668 39752
rect 2708 39712 2709 39752
rect 2667 39703 2709 39712
rect 2476 38912 2516 38921
rect 2476 38408 2516 38872
rect 2572 38912 2612 38921
rect 2572 38585 2612 38872
rect 2571 38576 2613 38585
rect 2571 38536 2572 38576
rect 2612 38536 2613 38576
rect 2571 38527 2613 38536
rect 2668 38408 2708 39703
rect 3052 38996 3092 40300
rect 3147 40300 3148 40340
rect 3188 40300 3189 40340
rect 3147 40291 3189 40300
rect 3148 40260 3188 40291
rect 3147 40088 3189 40097
rect 3147 40048 3148 40088
rect 3188 40048 3189 40088
rect 3147 40039 3189 40048
rect 2955 38912 2997 38921
rect 2955 38872 2956 38912
rect 2996 38872 2997 38912
rect 2955 38863 2997 38872
rect 2956 38778 2996 38863
rect 3052 38753 3092 38956
rect 3051 38744 3093 38753
rect 3051 38704 3052 38744
rect 3092 38704 3093 38744
rect 3051 38695 3093 38704
rect 3051 38576 3093 38585
rect 3051 38536 3052 38576
rect 3092 38536 3093 38576
rect 3051 38527 3093 38536
rect 2476 38368 2612 38408
rect 2476 38240 2516 38249
rect 2380 38200 2476 38240
rect 2380 37409 2420 38200
rect 2476 38191 2516 38200
rect 2379 37400 2421 37409
rect 2379 37360 2380 37400
rect 2420 37360 2421 37400
rect 2379 37351 2421 37360
rect 2476 37400 2516 37409
rect 2380 34376 2420 37351
rect 2476 36989 2516 37360
rect 2475 36980 2517 36989
rect 2475 36940 2476 36980
rect 2516 36940 2517 36980
rect 2475 36931 2517 36940
rect 2476 36728 2516 36737
rect 2476 35981 2516 36688
rect 2572 36140 2612 38368
rect 2668 38359 2708 38368
rect 2956 38240 2996 38249
rect 2956 37820 2996 38200
rect 2764 37780 2996 37820
rect 3052 38240 3092 38527
rect 2667 36896 2709 36905
rect 2667 36856 2668 36896
rect 2708 36856 2709 36896
rect 2667 36847 2709 36856
rect 2668 36762 2708 36847
rect 2668 36140 2708 36149
rect 2572 36100 2668 36140
rect 2668 36091 2708 36100
rect 2475 35972 2517 35981
rect 2475 35932 2476 35972
rect 2516 35932 2517 35972
rect 2475 35923 2517 35932
rect 2476 35888 2516 35923
rect 2476 35838 2516 35848
rect 2572 35216 2612 35225
rect 2476 34376 2516 34385
rect 2380 34336 2476 34376
rect 2476 33704 2516 34336
rect 2476 32864 2516 33664
rect 2476 32192 2516 32824
rect 2572 32360 2612 35176
rect 2667 35216 2709 35225
rect 2667 35176 2668 35216
rect 2708 35176 2709 35216
rect 2667 35167 2709 35176
rect 2668 35082 2708 35167
rect 2668 34628 2708 34637
rect 2764 34628 2804 37780
rect 2956 35888 2996 35897
rect 2708 34588 2804 34628
rect 2860 35848 2956 35888
rect 2668 34579 2708 34588
rect 2860 34376 2900 35848
rect 2956 35839 2996 35848
rect 3052 35888 3092 38200
rect 3148 36233 3188 40039
rect 3147 36224 3189 36233
rect 3147 36184 3148 36224
rect 3188 36184 3189 36224
rect 3147 36175 3189 36184
rect 3052 35309 3092 35848
rect 3051 35300 3093 35309
rect 3051 35260 3052 35300
rect 3092 35260 3093 35300
rect 3051 35251 3093 35260
rect 3051 35132 3093 35141
rect 3051 35092 3052 35132
rect 3092 35092 3093 35132
rect 3051 35083 3093 35092
rect 3148 35132 3188 35143
rect 3052 34998 3092 35083
rect 3148 35057 3188 35092
rect 3147 35048 3189 35057
rect 3147 35008 3148 35048
rect 3188 35008 3189 35048
rect 3147 34999 3189 35008
rect 3052 34385 3092 34470
rect 2668 34336 2900 34376
rect 3051 34376 3093 34385
rect 3051 34336 3052 34376
rect 3092 34336 3093 34376
rect 2668 33620 2708 34336
rect 3051 34327 3093 34336
rect 2763 34208 2805 34217
rect 2763 34168 2764 34208
rect 2804 34168 2805 34208
rect 2763 34159 2805 34168
rect 2860 34208 2900 34217
rect 2764 33872 2804 34159
rect 2860 34040 2900 34168
rect 3244 34133 3284 41224
rect 3723 41215 3765 41224
rect 3820 41264 3860 41551
rect 3820 41215 3860 41224
rect 3724 41130 3764 41215
rect 4012 41021 4052 42148
rect 4203 41936 4245 41945
rect 4203 41896 4204 41936
rect 4244 41896 4245 41936
rect 4203 41887 4245 41896
rect 4300 41936 4340 42727
rect 4396 42701 4436 42904
rect 4492 42785 4532 44248
rect 4875 44248 4876 44288
rect 4916 44248 4917 44288
rect 4875 44239 4917 44248
rect 4876 44154 4916 44239
rect 5068 43616 5108 43625
rect 5108 43576 5492 43616
rect 5068 43567 5108 43576
rect 4875 43448 4917 43457
rect 4875 43408 4876 43448
rect 4916 43408 4917 43448
rect 4875 43399 4917 43408
rect 5260 43448 5300 43457
rect 5300 43408 5396 43448
rect 5260 43399 5300 43408
rect 4876 43314 4916 43399
rect 4928 43112 5296 43121
rect 4968 43072 5010 43112
rect 5050 43072 5092 43112
rect 5132 43072 5174 43112
rect 5214 43072 5256 43112
rect 4928 43063 5296 43072
rect 5356 42953 5396 43408
rect 5355 42944 5397 42953
rect 5355 42904 5356 42944
rect 5396 42904 5397 42944
rect 5355 42895 5397 42904
rect 4876 42860 4916 42869
rect 4491 42776 4533 42785
rect 4491 42736 4492 42776
rect 4532 42736 4533 42776
rect 4491 42727 4533 42736
rect 4684 42762 4724 42771
rect 4395 42692 4437 42701
rect 4395 42652 4396 42692
rect 4436 42652 4437 42692
rect 4395 42643 4437 42652
rect 4396 42029 4436 42643
rect 4491 42608 4533 42617
rect 4491 42568 4492 42608
rect 4532 42568 4533 42608
rect 4491 42559 4533 42568
rect 4395 42020 4437 42029
rect 4395 41980 4396 42020
rect 4436 41980 4437 42020
rect 4395 41971 4437 41980
rect 4204 41802 4244 41887
rect 4300 41609 4340 41896
rect 4107 41600 4149 41609
rect 4107 41560 4108 41600
rect 4148 41560 4149 41600
rect 4107 41551 4149 41560
rect 4299 41600 4341 41609
rect 4299 41560 4300 41600
rect 4340 41560 4341 41600
rect 4299 41551 4341 41560
rect 4011 41012 4053 41021
rect 4011 40972 4012 41012
rect 4052 40972 4053 41012
rect 4011 40963 4053 40972
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 3339 40592 3381 40601
rect 3339 40552 3340 40592
rect 3380 40552 3381 40592
rect 3339 40543 3381 40552
rect 3340 40458 3380 40543
rect 3531 40508 3573 40517
rect 3531 40468 3532 40508
rect 3572 40468 3573 40508
rect 3531 40459 3573 40468
rect 3532 40424 3572 40459
rect 3532 40373 3572 40384
rect 3819 39752 3861 39761
rect 3819 39712 3820 39752
rect 3860 39712 3861 39752
rect 3819 39703 3861 39712
rect 3916 39752 3956 39761
rect 4108 39752 4148 41551
rect 4300 41264 4340 41273
rect 4396 41264 4436 41971
rect 4340 41224 4436 41264
rect 4300 41215 4340 41224
rect 4204 41180 4244 41189
rect 4204 41105 4244 41140
rect 4203 41096 4245 41105
rect 4203 41056 4204 41096
rect 4244 41056 4245 41096
rect 4203 41047 4245 41056
rect 3956 39712 4148 39752
rect 3916 39703 3956 39712
rect 3820 39618 3860 39703
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 4108 39089 4148 39712
rect 4204 39668 4244 41047
rect 4396 39752 4436 41224
rect 4492 41852 4532 42559
rect 4684 42197 4724 42722
rect 4683 42188 4725 42197
rect 4683 42148 4684 42188
rect 4724 42148 4725 42188
rect 4683 42139 4725 42148
rect 4779 42020 4821 42029
rect 4779 41980 4780 42020
rect 4820 41980 4821 42020
rect 4779 41971 4821 41980
rect 4684 41936 4724 41945
rect 4684 41852 4724 41896
rect 4780 41886 4820 41971
rect 4492 41812 4724 41852
rect 4492 41105 4532 41812
rect 4876 41768 4916 42820
rect 5259 42860 5301 42869
rect 5259 42820 5260 42860
rect 5300 42820 5301 42860
rect 5259 42811 5301 42820
rect 5067 42776 5109 42785
rect 5067 42736 5068 42776
rect 5108 42736 5109 42776
rect 5067 42727 5109 42736
rect 5068 41777 5108 42727
rect 5163 42524 5205 42533
rect 5163 42484 5164 42524
rect 5204 42484 5205 42524
rect 5163 42475 5205 42484
rect 5164 42390 5204 42475
rect 5260 41936 5300 42811
rect 5356 42776 5396 42785
rect 5356 42701 5396 42736
rect 5355 42692 5397 42701
rect 5355 42652 5356 42692
rect 5396 42652 5397 42692
rect 5355 42643 5397 42652
rect 5356 42449 5396 42643
rect 5355 42440 5397 42449
rect 5355 42400 5356 42440
rect 5396 42400 5397 42440
rect 5355 42391 5397 42400
rect 5356 42113 5396 42391
rect 5355 42104 5397 42113
rect 5355 42064 5356 42104
rect 5396 42064 5397 42104
rect 5355 42055 5397 42064
rect 5260 41777 5300 41896
rect 4588 41728 4916 41768
rect 5067 41768 5109 41777
rect 5067 41728 5068 41768
rect 5108 41728 5109 41768
rect 4491 41096 4533 41105
rect 4491 41056 4492 41096
rect 4532 41056 4533 41096
rect 4491 41047 4533 41056
rect 4299 39668 4341 39677
rect 4204 39628 4300 39668
rect 4340 39628 4341 39668
rect 4299 39619 4341 39628
rect 4300 39534 4340 39619
rect 4396 39416 4436 39712
rect 4300 39376 4436 39416
rect 4203 39248 4245 39257
rect 4203 39208 4204 39248
rect 4244 39208 4245 39248
rect 4203 39199 4245 39208
rect 4107 39080 4149 39089
rect 4107 39040 4108 39080
rect 4148 39040 4149 39080
rect 4107 39031 4149 39040
rect 3339 38912 3381 38921
rect 3339 38872 3340 38912
rect 3380 38872 3381 38912
rect 3339 38863 3381 38872
rect 3532 38912 3572 38921
rect 4012 38917 4052 38926
rect 3572 38872 3668 38912
rect 3532 38863 3572 38872
rect 3340 38249 3380 38863
rect 3531 38744 3573 38753
rect 3531 38704 3532 38744
rect 3572 38704 3573 38744
rect 3531 38695 3573 38704
rect 3339 38240 3381 38249
rect 3436 38240 3476 38268
rect 3339 38200 3340 38240
rect 3380 38200 3436 38240
rect 3339 38191 3381 38200
rect 3436 38191 3476 38200
rect 3532 38240 3572 38695
rect 3340 36896 3380 38191
rect 3532 38072 3572 38200
rect 3628 38165 3668 38872
rect 4012 38408 4052 38877
rect 4204 38828 4244 39199
rect 4204 38779 4244 38788
rect 3916 38368 4052 38408
rect 3627 38156 3669 38165
rect 3627 38116 3628 38156
rect 3668 38116 3669 38156
rect 3627 38107 3669 38116
rect 3436 38032 3572 38072
rect 3436 37073 3476 38032
rect 3916 37988 3956 38368
rect 4012 38240 4052 38249
rect 4012 38081 4052 38200
rect 4011 38072 4053 38081
rect 4011 38032 4012 38072
rect 4052 38032 4053 38072
rect 4011 38023 4053 38032
rect 3532 37948 3956 37988
rect 4107 37988 4149 37997
rect 4107 37948 4108 37988
rect 4148 37948 4149 37988
rect 3435 37064 3477 37073
rect 3435 37024 3436 37064
rect 3476 37024 3477 37064
rect 3435 37015 3477 37024
rect 3532 36905 3572 37948
rect 4107 37939 4149 37948
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 3916 37652 3956 37661
rect 4108 37652 4148 37939
rect 3956 37612 4148 37652
rect 3916 37603 3956 37612
rect 3723 37400 3765 37409
rect 3723 37360 3724 37400
rect 3764 37360 3765 37400
rect 3723 37351 3765 37360
rect 4108 37400 4148 37409
rect 3724 37266 3764 37351
rect 4108 37241 4148 37360
rect 4107 37232 4149 37241
rect 4107 37192 4108 37232
rect 4148 37192 4149 37232
rect 4107 37183 4149 37192
rect 3627 37064 3669 37073
rect 3627 37024 3628 37064
rect 3668 37024 3669 37064
rect 3627 37015 3669 37024
rect 3531 36896 3573 36905
rect 3340 36856 3476 36896
rect 3340 36728 3380 36737
rect 3340 36653 3380 36688
rect 3339 36644 3381 36653
rect 3339 36604 3340 36644
rect 3380 36604 3381 36644
rect 3339 36595 3381 36604
rect 3340 36401 3380 36595
rect 3339 36392 3381 36401
rect 3339 36352 3340 36392
rect 3380 36352 3381 36392
rect 3339 36343 3381 36352
rect 3339 35972 3381 35981
rect 3339 35932 3340 35972
rect 3380 35932 3381 35972
rect 3339 35923 3381 35932
rect 3243 34124 3285 34133
rect 3243 34084 3244 34124
rect 3284 34084 3285 34124
rect 3243 34075 3285 34084
rect 2860 34000 2996 34040
rect 2956 33881 2996 34000
rect 3051 33956 3093 33965
rect 3051 33916 3052 33956
rect 3092 33916 3093 33956
rect 3051 33907 3093 33916
rect 2860 33872 2900 33881
rect 2764 33832 2860 33872
rect 2860 33823 2900 33832
rect 2955 33872 2997 33881
rect 2955 33832 2956 33872
rect 2996 33832 2997 33872
rect 2955 33823 2997 33832
rect 2955 33704 2997 33713
rect 2955 33664 2956 33704
rect 2996 33664 2997 33704
rect 2955 33655 2997 33664
rect 2668 33580 2804 33620
rect 2667 33452 2709 33461
rect 2667 33412 2668 33452
rect 2708 33412 2709 33452
rect 2667 33403 2709 33412
rect 2668 33318 2708 33403
rect 2668 33116 2708 33125
rect 2764 33116 2804 33580
rect 2956 33570 2996 33655
rect 2708 33076 2804 33116
rect 2668 33067 2708 33076
rect 2859 32864 2901 32873
rect 2859 32824 2860 32864
rect 2900 32824 2901 32864
rect 2859 32815 2901 32824
rect 3052 32864 3092 33907
rect 3243 33872 3285 33881
rect 3243 33832 3244 33872
rect 3284 33832 3285 33872
rect 3243 33823 3285 33832
rect 3244 33738 3284 33823
rect 3340 33041 3380 35923
rect 3436 35888 3476 36856
rect 3531 36856 3532 36896
rect 3572 36856 3573 36896
rect 3531 36847 3573 36856
rect 3628 36728 3668 37015
rect 3436 35141 3476 35848
rect 3532 36688 3668 36728
rect 3532 35888 3572 36688
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 3723 36140 3765 36149
rect 3723 36100 3724 36140
rect 3764 36100 3765 36140
rect 3723 36091 3765 36100
rect 4011 36140 4053 36149
rect 4011 36100 4012 36140
rect 4052 36100 4053 36140
rect 4011 36091 4053 36100
rect 3435 35132 3477 35141
rect 3435 35092 3436 35132
rect 3476 35092 3477 35132
rect 3435 35083 3477 35092
rect 3532 35057 3572 35848
rect 3627 35216 3669 35225
rect 3627 35176 3628 35216
rect 3668 35176 3669 35216
rect 3627 35167 3669 35176
rect 3628 35082 3668 35167
rect 3531 35048 3573 35057
rect 3531 35008 3532 35048
rect 3572 35008 3573 35048
rect 3531 34999 3573 35008
rect 3724 34973 3764 36091
rect 4012 35888 4052 36091
rect 4012 35225 4052 35848
rect 4300 35468 4340 39376
rect 4492 38226 4532 38235
rect 4492 37997 4532 38186
rect 4491 37988 4533 37997
rect 4491 37948 4492 37988
rect 4532 37948 4533 37988
rect 4491 37939 4533 37948
rect 4588 37820 4628 41728
rect 5067 41719 5109 41728
rect 5259 41768 5301 41777
rect 5259 41728 5260 41768
rect 5300 41728 5301 41768
rect 5259 41719 5301 41728
rect 4779 41600 4821 41609
rect 4779 41560 4780 41600
rect 4820 41560 4821 41600
rect 4779 41551 4821 41560
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 4780 41264 4820 41551
rect 5452 41516 5492 43576
rect 5548 42281 5588 44920
rect 5547 42272 5589 42281
rect 5547 42232 5548 42272
rect 5588 42232 5589 42272
rect 5547 42223 5589 42232
rect 5644 41609 5684 47515
rect 5739 47396 5781 47405
rect 5739 47356 5740 47396
rect 5780 47356 5781 47396
rect 5739 47347 5781 47356
rect 5740 42869 5780 47347
rect 5835 46220 5877 46229
rect 5835 46180 5836 46220
rect 5876 46180 5877 46220
rect 5835 46171 5877 46180
rect 5836 45800 5876 46171
rect 5836 45641 5876 45760
rect 5932 45800 5972 48784
rect 6124 47825 6164 49363
rect 6219 49076 6261 49085
rect 6219 49036 6220 49076
rect 6260 49036 6261 49076
rect 6219 49027 6261 49036
rect 6220 48833 6260 49027
rect 6315 48908 6357 48917
rect 6315 48868 6316 48908
rect 6356 48868 6357 48908
rect 6315 48859 6357 48868
rect 6219 48824 6261 48833
rect 6219 48784 6220 48824
rect 6260 48784 6261 48824
rect 6219 48775 6261 48784
rect 6316 48824 6356 48859
rect 6220 48690 6260 48775
rect 6123 47816 6165 47825
rect 6123 47776 6124 47816
rect 6164 47776 6165 47816
rect 6123 47767 6165 47776
rect 6123 47312 6165 47321
rect 6123 47272 6124 47312
rect 6164 47272 6165 47312
rect 6123 47263 6165 47272
rect 6124 46556 6164 47263
rect 6316 46901 6356 48784
rect 6412 47657 6452 50296
rect 6507 49244 6549 49253
rect 6507 49204 6508 49244
rect 6548 49204 6549 49244
rect 6507 49195 6549 49204
rect 6508 48833 6548 49195
rect 6507 48824 6549 48833
rect 6507 48784 6508 48824
rect 6548 48784 6549 48824
rect 6507 48775 6549 48784
rect 6411 47648 6453 47657
rect 6411 47608 6412 47648
rect 6452 47608 6453 47648
rect 6411 47599 6453 47608
rect 6412 47480 6452 47489
rect 6315 46892 6357 46901
rect 6315 46852 6316 46892
rect 6356 46852 6357 46892
rect 6315 46843 6357 46852
rect 6412 46640 6452 47440
rect 6220 46565 6260 46609
rect 6316 46600 6452 46640
rect 6219 46556 6261 46565
rect 6124 46514 6165 46556
rect 6164 46474 6165 46514
rect 6219 46516 6220 46556
rect 6260 46516 6261 46556
rect 6219 46514 6261 46516
rect 6219 46507 6220 46514
rect 6260 46507 6261 46514
rect 6124 46465 6164 46474
rect 6220 46465 6260 46474
rect 6316 46472 6356 46600
rect 6316 46423 6356 46432
rect 6411 46472 6453 46481
rect 6411 46432 6412 46472
rect 6452 46432 6453 46472
rect 6411 46423 6453 46432
rect 6412 46338 6452 46423
rect 6315 46052 6357 46061
rect 6315 46012 6316 46052
rect 6356 46012 6357 46052
rect 6315 46003 6357 46012
rect 6219 45884 6261 45893
rect 6219 45844 6220 45884
rect 6260 45844 6261 45884
rect 6219 45835 6261 45844
rect 5835 45632 5877 45641
rect 5835 45592 5836 45632
rect 5876 45592 5877 45632
rect 5835 45583 5877 45592
rect 5932 45389 5972 45760
rect 6027 45716 6069 45725
rect 6027 45676 6028 45716
rect 6068 45676 6069 45716
rect 6027 45667 6069 45676
rect 5931 45380 5973 45389
rect 5931 45340 5932 45380
rect 5972 45340 5973 45380
rect 5931 45331 5973 45340
rect 5739 42860 5781 42869
rect 5739 42820 5740 42860
rect 5780 42820 5781 42860
rect 5739 42811 5781 42820
rect 5835 42776 5877 42785
rect 5835 42736 5836 42776
rect 5876 42736 5877 42776
rect 5835 42727 5877 42736
rect 5739 42524 5781 42533
rect 5739 42484 5740 42524
rect 5780 42484 5781 42524
rect 5739 42475 5781 42484
rect 5740 41950 5780 42475
rect 5740 41901 5780 41910
rect 5643 41600 5685 41609
rect 5643 41560 5644 41600
rect 5684 41560 5685 41600
rect 5643 41551 5685 41560
rect 5356 41476 5492 41516
rect 5356 41264 5396 41476
rect 5739 41432 5781 41441
rect 5739 41392 5740 41432
rect 5780 41392 5781 41432
rect 5739 41383 5781 41392
rect 4684 41224 4780 41264
rect 4684 39752 4724 41224
rect 4780 41215 4820 41224
rect 5308 41254 5396 41264
rect 5348 41224 5396 41254
rect 5452 41348 5492 41357
rect 5308 41205 5348 41214
rect 5163 41012 5205 41021
rect 5163 40972 5164 41012
rect 5204 40972 5205 41012
rect 5163 40963 5205 40972
rect 4779 40760 4821 40769
rect 4779 40720 4780 40760
rect 4820 40720 4821 40760
rect 4779 40711 4821 40720
rect 4780 40424 4820 40711
rect 4780 40375 4820 40384
rect 4972 40349 5012 40434
rect 5164 40433 5204 40963
rect 5355 40592 5397 40601
rect 5355 40552 5356 40592
rect 5396 40552 5397 40592
rect 5355 40543 5397 40552
rect 5163 40424 5205 40433
rect 5163 40384 5164 40424
rect 5204 40384 5205 40424
rect 5163 40375 5205 40384
rect 4971 40340 5013 40349
rect 4971 40300 4972 40340
rect 5012 40300 5013 40340
rect 4971 40291 5013 40300
rect 5164 40290 5204 40375
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 4876 39752 4916 39761
rect 4684 39712 4876 39752
rect 4876 39703 4916 39712
rect 5163 39752 5205 39761
rect 5163 39712 5164 39752
rect 5204 39712 5205 39752
rect 5163 39703 5205 39712
rect 5356 39747 5396 40543
rect 4683 38996 4725 39005
rect 4683 38956 4684 38996
rect 4724 38956 4725 38996
rect 4683 38947 4725 38956
rect 4684 38408 4724 38947
rect 5164 38921 5204 39703
rect 5356 39698 5396 39707
rect 5163 38912 5205 38921
rect 5163 38872 5164 38912
rect 5204 38872 5205 38912
rect 5163 38863 5205 38872
rect 5355 38912 5397 38921
rect 5355 38872 5356 38912
rect 5396 38872 5397 38912
rect 5355 38863 5397 38872
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 4684 38359 4724 38368
rect 5356 37820 5396 38863
rect 5452 38417 5492 41308
rect 5643 40424 5685 40433
rect 5643 40384 5644 40424
rect 5684 40384 5685 40424
rect 5643 40375 5685 40384
rect 5548 39836 5588 39845
rect 5451 38408 5493 38417
rect 5451 38368 5452 38408
rect 5492 38368 5493 38408
rect 5451 38359 5493 38368
rect 5451 38156 5493 38165
rect 5451 38116 5452 38156
rect 5492 38116 5493 38156
rect 5451 38107 5493 38116
rect 4204 35428 4340 35468
rect 4396 37780 4628 37820
rect 5260 37780 5396 37820
rect 4011 35216 4053 35225
rect 4011 35176 4012 35216
rect 4052 35176 4053 35216
rect 4011 35167 4053 35176
rect 4108 35202 4148 35211
rect 3723 34964 3765 34973
rect 3723 34924 3724 34964
rect 3764 34924 3765 34964
rect 3723 34915 3765 34924
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 3435 33788 3477 33797
rect 3435 33748 3436 33788
rect 3476 33748 3477 33788
rect 3435 33739 3477 33748
rect 3436 33699 3476 33739
rect 3436 33650 3476 33659
rect 3915 33704 3957 33713
rect 3915 33664 3916 33704
rect 3956 33664 3957 33704
rect 3915 33655 3957 33664
rect 3916 33570 3956 33655
rect 4108 33461 4148 35162
rect 4204 33965 4244 35428
rect 4396 35384 4436 37780
rect 4587 37400 4629 37409
rect 4587 37360 4588 37400
rect 4628 37360 4629 37400
rect 4587 37351 4629 37360
rect 4588 36728 4628 37351
rect 5260 37241 5300 37780
rect 5355 37400 5397 37409
rect 5355 37360 5356 37400
rect 5396 37360 5397 37400
rect 5355 37351 5397 37360
rect 5356 37266 5396 37351
rect 5259 37232 5301 37241
rect 5259 37192 5260 37232
rect 5300 37192 5301 37232
rect 5259 37183 5301 37192
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 4588 36679 4628 36688
rect 4875 36560 4917 36569
rect 4875 36520 4876 36560
rect 4916 36520 4917 36560
rect 4875 36511 4917 36520
rect 4780 36476 4820 36485
rect 4684 36436 4780 36476
rect 4684 35972 4724 36436
rect 4780 36427 4820 36436
rect 4876 36308 4916 36511
rect 4540 35932 4724 35972
rect 4780 36268 4916 36308
rect 4540 35930 4580 35932
rect 4540 35881 4580 35890
rect 4684 35720 4724 35729
rect 4396 35344 4532 35384
rect 4300 35300 4340 35309
rect 4340 35260 4436 35300
rect 4300 35251 4340 35260
rect 4300 34469 4340 34500
rect 4299 34460 4341 34469
rect 4299 34420 4300 34460
rect 4340 34420 4341 34460
rect 4299 34411 4341 34420
rect 4300 34376 4340 34411
rect 4300 34133 4340 34336
rect 4299 34124 4341 34133
rect 4299 34084 4300 34124
rect 4340 34084 4341 34124
rect 4299 34075 4341 34084
rect 4203 33956 4245 33965
rect 4203 33916 4204 33956
rect 4244 33916 4245 33956
rect 4203 33907 4245 33916
rect 4396 33881 4436 35260
rect 4492 35057 4532 35344
rect 4491 35048 4533 35057
rect 4491 35008 4492 35048
rect 4532 35008 4533 35048
rect 4491 34999 4533 35008
rect 4492 34376 4532 34387
rect 4492 34301 4532 34336
rect 4587 34376 4629 34385
rect 4587 34336 4588 34376
rect 4628 34336 4629 34376
rect 4587 34327 4629 34336
rect 4491 34292 4533 34301
rect 4491 34252 4492 34292
rect 4532 34252 4533 34292
rect 4491 34243 4533 34252
rect 4492 34049 4532 34243
rect 4491 34040 4533 34049
rect 4491 34000 4492 34040
rect 4532 34000 4533 34040
rect 4491 33991 4533 34000
rect 4395 33872 4437 33881
rect 4395 33832 4396 33872
rect 4436 33832 4437 33872
rect 4395 33823 4437 33832
rect 4203 33704 4245 33713
rect 4203 33664 4204 33704
rect 4244 33664 4245 33704
rect 4203 33655 4245 33664
rect 4107 33452 4149 33461
rect 4107 33412 4108 33452
rect 4148 33412 4149 33452
rect 4107 33403 4149 33412
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 3916 33116 3956 33125
rect 4204 33116 4244 33655
rect 4395 33620 4437 33629
rect 4395 33580 4396 33620
rect 4436 33580 4437 33620
rect 4395 33571 4437 33580
rect 4492 33620 4532 33629
rect 4396 33486 4436 33571
rect 4492 33461 4532 33580
rect 4491 33452 4533 33461
rect 4491 33412 4492 33452
rect 4532 33412 4533 33452
rect 4491 33403 4533 33412
rect 4395 33284 4437 33293
rect 4395 33244 4396 33284
rect 4436 33244 4437 33284
rect 4395 33235 4437 33244
rect 3956 33076 4244 33116
rect 3916 33067 3956 33076
rect 3339 33032 3381 33041
rect 3339 32992 3340 33032
rect 3380 32992 3381 33032
rect 3339 32983 3381 32992
rect 3374 32873 3414 32880
rect 2860 32696 2900 32815
rect 2860 32647 2900 32656
rect 2668 32360 2708 32369
rect 2572 32320 2668 32360
rect 2668 32311 2708 32320
rect 2476 32117 2516 32152
rect 2859 32192 2901 32201
rect 2859 32152 2860 32192
rect 2900 32152 2901 32192
rect 2859 32143 2901 32152
rect 2475 32108 2517 32117
rect 2475 32068 2476 32108
rect 2516 32068 2517 32108
rect 2475 32059 2517 32068
rect 2763 32108 2805 32117
rect 2763 32068 2764 32108
rect 2804 32068 2805 32108
rect 2763 32059 2805 32068
rect 2475 31940 2517 31949
rect 2475 31900 2476 31940
rect 2516 31900 2517 31940
rect 2475 31891 2517 31900
rect 2380 31361 2420 31446
rect 2379 31352 2421 31361
rect 2379 31312 2380 31352
rect 2420 31312 2421 31352
rect 2379 31303 2421 31312
rect 2476 31352 2516 31891
rect 2476 30689 2516 31312
rect 2475 30680 2517 30689
rect 2475 30640 2476 30680
rect 2516 30640 2517 30680
rect 2475 30631 2517 30640
rect 2667 30092 2709 30101
rect 2667 30052 2668 30092
rect 2708 30052 2709 30092
rect 2667 30043 2709 30052
rect 2668 29429 2708 30043
rect 2667 29420 2709 29429
rect 2667 29380 2668 29420
rect 2708 29380 2709 29420
rect 2667 29371 2709 29380
rect 2283 29336 2325 29345
rect 2283 29296 2284 29336
rect 2324 29296 2325 29336
rect 2283 29287 2325 29296
rect 2187 29168 2229 29177
rect 2187 29128 2188 29168
rect 2228 29128 2229 29168
rect 2476 29168 2516 29177
rect 2668 29168 2708 29371
rect 2187 29119 2229 29128
rect 2320 29158 2360 29167
rect 2188 29034 2228 29119
rect 2516 29128 2708 29168
rect 2476 29119 2516 29128
rect 2320 29093 2360 29118
rect 2283 29084 2360 29093
rect 2283 29044 2284 29084
rect 2324 29044 2360 29084
rect 2283 29035 2325 29044
rect 2379 28832 2421 28841
rect 2379 28792 2380 28832
rect 2420 28792 2421 28832
rect 2379 28783 2421 28792
rect 2283 26480 2325 26489
rect 2283 26440 2284 26480
rect 2324 26440 2325 26480
rect 2283 26431 2325 26440
rect 2036 25516 2132 25556
rect 1996 25507 2036 25516
rect 2187 25388 2229 25397
rect 2187 25348 2188 25388
rect 2228 25348 2229 25388
rect 2187 25339 2229 25348
rect 2188 25304 2228 25339
rect 1900 25264 2132 25304
rect 1899 25136 1941 25145
rect 1899 25096 1900 25136
rect 1940 25096 1941 25136
rect 1899 25087 1941 25096
rect 1516 23911 1556 23920
rect 1612 24256 1844 24296
rect 1323 23204 1365 23213
rect 1323 23164 1324 23204
rect 1364 23164 1365 23204
rect 1323 23155 1365 23164
rect 1228 22280 1268 22289
rect 1323 22280 1365 22289
rect 1268 22240 1324 22280
rect 1364 22240 1365 22280
rect 1228 22231 1268 22240
rect 1323 22231 1365 22240
rect 1515 21608 1557 21617
rect 1515 21568 1516 21608
rect 1556 21568 1557 21608
rect 1515 21559 1557 21568
rect 1516 21474 1556 21559
rect 1515 20936 1557 20945
rect 1515 20896 1516 20936
rect 1556 20896 1557 20936
rect 1515 20887 1557 20896
rect 1228 20768 1268 20777
rect 1132 20728 1228 20768
rect 1228 20719 1268 20728
rect 1228 20096 1268 20105
rect 1419 20096 1461 20105
rect 1268 20056 1420 20096
rect 1460 20056 1461 20096
rect 1228 20047 1268 20056
rect 1419 20047 1461 20056
rect 1228 19256 1268 19265
rect 1268 19216 1364 19256
rect 1228 19207 1268 19216
rect 1324 19097 1364 19216
rect 1323 19088 1365 19097
rect 1323 19048 1324 19088
rect 1364 19048 1365 19088
rect 1323 19039 1365 19048
rect 1228 18584 1268 18593
rect 1268 18544 1364 18584
rect 1228 18535 1268 18544
rect 1131 18332 1173 18341
rect 1131 18292 1132 18332
rect 1172 18292 1173 18332
rect 1131 18283 1173 18292
rect 1132 16904 1172 18283
rect 1324 17249 1364 18544
rect 1323 17240 1365 17249
rect 1323 17200 1324 17240
rect 1364 17200 1365 17240
rect 1323 17191 1365 17200
rect 1228 17072 1268 17081
rect 1420 17072 1460 20047
rect 1516 18164 1556 20887
rect 1612 18341 1652 24256
rect 1803 23876 1845 23885
rect 1803 23836 1804 23876
rect 1844 23836 1845 23876
rect 1803 23827 1845 23836
rect 1804 23742 1844 23827
rect 1900 23717 1940 25087
rect 1996 24632 2036 24641
rect 1996 24473 2036 24592
rect 1995 24464 2037 24473
rect 1995 24424 1996 24464
rect 2036 24424 2037 24464
rect 1995 24415 2037 24424
rect 1995 23876 2037 23885
rect 1995 23836 1996 23876
rect 2036 23836 2037 23876
rect 1995 23827 2037 23836
rect 1996 23792 2036 23827
rect 1996 23741 2036 23752
rect 1899 23708 1941 23717
rect 1899 23668 1900 23708
rect 1940 23668 1941 23708
rect 1899 23659 1941 23668
rect 2092 23633 2132 25264
rect 2188 25253 2228 25264
rect 2091 23624 2133 23633
rect 2091 23584 2092 23624
rect 2132 23584 2133 23624
rect 2091 23575 2133 23584
rect 1995 23540 2037 23549
rect 1995 23500 1996 23540
rect 2036 23500 2037 23540
rect 1995 23491 2037 23500
rect 1708 23120 1748 23129
rect 1708 20357 1748 23080
rect 1707 20348 1749 20357
rect 1707 20308 1708 20348
rect 1748 20308 1749 20348
rect 1707 20299 1749 20308
rect 1707 19760 1749 19769
rect 1707 19720 1708 19760
rect 1748 19720 1749 19760
rect 1707 19711 1749 19720
rect 1611 18332 1653 18341
rect 1611 18292 1612 18332
rect 1652 18292 1653 18332
rect 1611 18283 1653 18292
rect 1516 18124 1652 18164
rect 1515 17996 1557 18005
rect 1515 17956 1516 17996
rect 1556 17956 1557 17996
rect 1515 17947 1557 17956
rect 1268 17032 1460 17072
rect 1228 17023 1268 17032
rect 1132 16864 1364 16904
rect 1324 15308 1364 16864
rect 1516 15392 1556 17947
rect 1612 15821 1652 18124
rect 1708 17576 1748 19711
rect 1803 18332 1845 18341
rect 1803 18292 1804 18332
rect 1844 18292 1845 18332
rect 1803 18283 1845 18292
rect 1804 17744 1844 18283
rect 1900 17795 1940 17852
rect 1899 17786 1941 17795
rect 1899 17737 1900 17786
rect 1940 17737 1941 17786
rect 1900 17708 1940 17717
rect 1804 17695 1844 17704
rect 1708 17536 1940 17576
rect 1803 17408 1845 17417
rect 1803 17368 1804 17408
rect 1844 17368 1845 17408
rect 1803 17359 1845 17368
rect 1707 16232 1749 16241
rect 1707 16192 1708 16232
rect 1748 16192 1749 16232
rect 1707 16183 1749 16192
rect 1611 15812 1653 15821
rect 1611 15772 1612 15812
rect 1652 15772 1653 15812
rect 1611 15763 1653 15772
rect 1612 15560 1652 15569
rect 1708 15560 1748 16183
rect 1652 15520 1748 15560
rect 1612 15511 1652 15520
rect 1516 15352 1652 15392
rect 1324 15268 1556 15308
rect 1228 14720 1268 14729
rect 1323 14720 1365 14729
rect 1268 14680 1324 14720
rect 1364 14680 1365 14720
rect 1228 14671 1268 14680
rect 1323 14671 1365 14680
rect 1227 14552 1269 14561
rect 1227 14512 1228 14552
rect 1268 14512 1269 14552
rect 1227 14503 1269 14512
rect 1035 13712 1077 13721
rect 1035 13672 1036 13712
rect 1076 13672 1077 13712
rect 1035 13663 1077 13672
rect 1228 12536 1268 14503
rect 1516 13301 1556 15268
rect 1515 13292 1557 13301
rect 1515 13252 1516 13292
rect 1556 13252 1557 13292
rect 1515 13243 1557 13252
rect 1420 12545 1460 12630
rect 1228 12487 1268 12496
rect 1419 12536 1461 12545
rect 1419 12496 1420 12536
rect 1460 12496 1461 12536
rect 1419 12487 1461 12496
rect 1516 12536 1556 12545
rect 1420 12368 1460 12377
rect 1228 11696 1268 11705
rect 459 11360 501 11369
rect 459 11320 460 11360
rect 500 11320 501 11360
rect 459 11311 501 11320
rect 1228 11201 1268 11656
rect 1420 11696 1460 12328
rect 1516 11873 1556 12496
rect 1515 11864 1557 11873
rect 1515 11824 1516 11864
rect 1556 11824 1557 11864
rect 1515 11815 1557 11824
rect 1420 11647 1460 11656
rect 1516 11696 1556 11705
rect 1323 11528 1365 11537
rect 1323 11488 1324 11528
rect 1364 11488 1365 11528
rect 1323 11479 1365 11488
rect 1324 11394 1364 11479
rect 1516 11453 1556 11656
rect 1515 11444 1557 11453
rect 1515 11404 1516 11444
rect 1556 11404 1557 11444
rect 1515 11395 1557 11404
rect 1227 11192 1269 11201
rect 1227 11152 1228 11192
rect 1268 11152 1269 11192
rect 1227 11143 1269 11152
rect 1228 11024 1268 11033
rect 1323 11024 1365 11033
rect 1268 10984 1324 11024
rect 1364 10984 1365 11024
rect 1228 10975 1268 10984
rect 1323 10975 1365 10984
rect 1228 10184 1268 10193
rect 1612 10184 1652 15352
rect 1708 14048 1748 15520
rect 1804 14225 1844 17359
rect 1900 15821 1940 17536
rect 1996 15989 2036 23491
rect 2187 20768 2229 20777
rect 2187 20728 2188 20768
rect 2228 20728 2229 20768
rect 2187 20719 2229 20728
rect 2091 18500 2133 18509
rect 2091 18460 2092 18500
rect 2132 18460 2133 18500
rect 2091 18451 2133 18460
rect 2092 17996 2132 18451
rect 2188 18005 2228 20719
rect 2092 17947 2132 17956
rect 2187 17996 2229 18005
rect 2187 17956 2188 17996
rect 2228 17956 2229 17996
rect 2187 17947 2229 17956
rect 2187 17828 2229 17837
rect 2092 17788 2188 17828
rect 2228 17788 2229 17828
rect 2092 17744 2132 17788
rect 2187 17779 2229 17788
rect 2092 17695 2132 17704
rect 2187 17408 2229 17417
rect 2187 17368 2188 17408
rect 2228 17368 2229 17408
rect 2187 17359 2229 17368
rect 2091 17240 2133 17249
rect 2091 17200 2092 17240
rect 2132 17200 2133 17240
rect 2091 17191 2133 17200
rect 1995 15980 2037 15989
rect 1995 15940 1996 15980
rect 2036 15940 2037 15980
rect 1995 15931 2037 15940
rect 1899 15812 1941 15821
rect 1899 15772 1900 15812
rect 1940 15772 1941 15812
rect 1899 15763 1941 15772
rect 1995 15728 2037 15737
rect 1995 15688 1996 15728
rect 2036 15688 2037 15728
rect 1995 15679 2037 15688
rect 1899 15560 1941 15569
rect 1899 15520 1900 15560
rect 1940 15520 1941 15560
rect 1899 15511 1941 15520
rect 1803 14216 1845 14225
rect 1803 14176 1804 14216
rect 1844 14176 1845 14216
rect 1803 14167 1845 14176
rect 1708 13999 1748 14008
rect 1708 13217 1748 13302
rect 1707 13208 1749 13217
rect 1707 13168 1708 13208
rect 1748 13168 1749 13208
rect 1707 13159 1749 13168
rect 1707 12956 1749 12965
rect 1707 12916 1708 12956
rect 1748 12916 1749 12956
rect 1707 12907 1749 12916
rect 1708 12536 1748 12907
rect 1803 12788 1845 12797
rect 1803 12748 1804 12788
rect 1844 12748 1845 12788
rect 1803 12739 1845 12748
rect 1708 12487 1748 12496
rect 1708 11696 1748 11705
rect 1804 11696 1844 12739
rect 1748 11656 1844 11696
rect 1708 11647 1748 11656
rect 1900 10772 1940 15511
rect 1996 13217 2036 15679
rect 1995 13208 2037 13217
rect 1995 13168 1996 13208
rect 2036 13168 2037 13208
rect 1995 13159 2037 13168
rect 1995 12536 2037 12545
rect 1995 12496 1996 12536
rect 2036 12496 2037 12536
rect 1995 12487 2037 12496
rect 1996 10949 2036 12487
rect 2092 11285 2132 17191
rect 2188 14384 2228 17359
rect 2284 16400 2324 26431
rect 2380 23549 2420 28783
rect 2571 26732 2613 26741
rect 2571 26692 2572 26732
rect 2612 26692 2613 26732
rect 2571 26683 2613 26692
rect 2379 23540 2421 23549
rect 2379 23500 2380 23540
rect 2420 23500 2421 23540
rect 2379 23491 2421 23500
rect 2475 22364 2517 22373
rect 2475 22324 2476 22364
rect 2516 22324 2517 22364
rect 2475 22315 2517 22324
rect 2476 22280 2516 22315
rect 2476 20768 2516 22240
rect 2476 20096 2516 20728
rect 2572 20525 2612 26683
rect 2668 25313 2708 29128
rect 2667 25304 2709 25313
rect 2667 25264 2668 25304
rect 2708 25264 2709 25304
rect 2667 25255 2709 25264
rect 2764 23801 2804 32059
rect 2860 32058 2900 32143
rect 2956 31436 2996 31445
rect 3052 31436 3092 32824
rect 3148 32871 3414 32873
rect 3148 32864 3374 32871
rect 3188 32833 3374 32864
rect 3148 32815 3188 32824
rect 3532 32864 3572 32873
rect 3147 32696 3189 32705
rect 3147 32656 3148 32696
rect 3188 32656 3189 32696
rect 3147 32647 3189 32656
rect 2996 31396 3092 31436
rect 2956 31387 2996 31396
rect 2860 31352 2900 31361
rect 2860 31109 2900 31312
rect 2859 31100 2901 31109
rect 2859 31060 2860 31100
rect 2900 31060 2901 31100
rect 2859 31051 2901 31060
rect 3148 30428 3188 32647
rect 3374 32528 3414 32831
rect 3531 32824 3532 32864
rect 3531 32782 3572 32824
rect 3532 32537 3572 32782
rect 3628 32864 3668 32873
rect 3244 32488 3414 32528
rect 3531 32528 3573 32537
rect 3531 32488 3532 32528
rect 3572 32488 3573 32528
rect 3244 32117 3284 32488
rect 3531 32479 3573 32488
rect 3531 32192 3573 32201
rect 3628 32192 3668 32824
rect 3819 32864 3861 32873
rect 3819 32824 3820 32864
rect 3860 32824 3861 32864
rect 3819 32815 3861 32824
rect 3916 32864 3956 32873
rect 3820 32730 3860 32815
rect 3916 32360 3956 32824
rect 4107 32864 4149 32873
rect 4107 32824 4108 32864
rect 4148 32824 4149 32864
rect 4107 32815 4149 32824
rect 4108 32730 4148 32815
rect 4300 32360 4340 32369
rect 4396 32360 4436 33235
rect 4588 32780 4628 34327
rect 4684 32957 4724 35680
rect 4780 35216 4820 36268
rect 5260 35888 5300 35897
rect 5452 35888 5492 38107
rect 5548 37820 5588 39796
rect 5644 38921 5684 40375
rect 5740 39761 5780 41383
rect 5739 39752 5781 39761
rect 5739 39712 5740 39752
rect 5780 39712 5781 39752
rect 5739 39703 5781 39712
rect 5739 39080 5781 39089
rect 5739 39040 5740 39080
rect 5780 39040 5781 39080
rect 5739 39031 5781 39040
rect 5643 38912 5685 38921
rect 5643 38872 5644 38912
rect 5684 38872 5685 38912
rect 5643 38863 5685 38872
rect 5740 38912 5780 39031
rect 5740 38863 5780 38872
rect 5836 38165 5876 42727
rect 6028 41936 6068 45667
rect 6123 44288 6165 44297
rect 6123 44248 6124 44288
rect 6164 44248 6165 44288
rect 6123 44239 6165 44248
rect 6124 44154 6164 44239
rect 6220 43457 6260 45835
rect 6316 45800 6356 46003
rect 6411 45884 6453 45893
rect 6411 45844 6412 45884
rect 6452 45844 6453 45884
rect 6411 45835 6453 45844
rect 6316 45751 6356 45760
rect 6412 45800 6452 45835
rect 6508 45800 6548 48775
rect 6604 47984 6644 47995
rect 6604 47909 6644 47944
rect 6603 47900 6645 47909
rect 6603 47860 6604 47900
rect 6644 47860 6645 47900
rect 6700 47900 6740 51640
rect 6891 50672 6933 50681
rect 6891 50632 6892 50672
rect 6932 50632 6933 50672
rect 6891 50623 6933 50632
rect 6892 49496 6932 50623
rect 6892 49421 6932 49456
rect 6891 49412 6933 49421
rect 6891 49372 6892 49412
rect 6932 49372 6933 49412
rect 6891 49363 6933 49372
rect 6988 48917 7028 52900
rect 7084 52613 7124 53992
rect 7180 53360 7220 54151
rect 7275 54032 7317 54041
rect 7275 53992 7276 54032
rect 7316 53992 7317 54032
rect 7275 53983 7317 53992
rect 7276 53898 7316 53983
rect 7180 53311 7220 53320
rect 7275 53276 7317 53285
rect 7275 53236 7276 53276
rect 7316 53236 7317 53276
rect 7275 53227 7317 53236
rect 7276 53142 7316 53227
rect 7179 52688 7221 52697
rect 7179 52648 7180 52688
rect 7220 52648 7221 52688
rect 7179 52639 7221 52648
rect 7083 52604 7125 52613
rect 7083 52564 7084 52604
rect 7124 52564 7125 52604
rect 7083 52555 7125 52564
rect 7083 52436 7125 52445
rect 7083 52396 7084 52436
rect 7124 52396 7125 52436
rect 7083 52387 7125 52396
rect 7084 51353 7124 52387
rect 7180 52025 7220 52639
rect 7179 52016 7221 52025
rect 7179 51976 7180 52016
rect 7220 51976 7221 52016
rect 7179 51967 7221 51976
rect 7179 51848 7221 51857
rect 7179 51808 7180 51848
rect 7220 51808 7221 51848
rect 7179 51799 7221 51808
rect 7276 51848 7316 51857
rect 7372 51848 7412 54160
rect 7468 53537 7508 54412
rect 7564 54209 7604 54907
rect 7756 54872 7796 55327
rect 7660 54832 7796 54872
rect 7563 54200 7605 54209
rect 7563 54160 7564 54200
rect 7604 54160 7605 54200
rect 7563 54151 7605 54160
rect 7563 53612 7605 53621
rect 7563 53572 7564 53612
rect 7604 53572 7605 53612
rect 7563 53563 7605 53572
rect 7467 53528 7509 53537
rect 7467 53488 7468 53528
rect 7508 53488 7509 53528
rect 7467 53479 7509 53488
rect 7316 51808 7508 51848
rect 7276 51799 7316 51808
rect 7083 51344 7125 51353
rect 7083 51304 7084 51344
rect 7124 51304 7125 51344
rect 7083 51295 7125 51304
rect 7084 50597 7124 51295
rect 7083 50588 7125 50597
rect 7083 50548 7084 50588
rect 7124 50548 7125 50588
rect 7083 50539 7125 50548
rect 7083 49748 7125 49757
rect 7083 49708 7084 49748
rect 7124 49708 7125 49748
rect 7180 49748 7220 51799
rect 7371 51680 7413 51689
rect 7371 51640 7372 51680
rect 7412 51640 7413 51680
rect 7371 51631 7413 51640
rect 7372 50336 7412 51631
rect 7468 51017 7508 51808
rect 7564 51269 7604 53563
rect 7660 53453 7700 54832
rect 7852 54452 7892 56092
rect 7947 56092 7948 56132
rect 7988 56092 7989 56132
rect 7947 56083 7989 56092
rect 7948 55460 7988 56083
rect 8140 56048 8180 56839
rect 8332 56636 8372 63979
rect 8428 63533 8468 66592
rect 8523 66380 8565 66389
rect 8523 66340 8524 66380
rect 8564 66340 8565 66380
rect 8523 66331 8565 66340
rect 8524 65549 8564 66331
rect 8523 65540 8565 65549
rect 8523 65500 8524 65540
rect 8564 65500 8565 65540
rect 8523 65491 8565 65500
rect 8716 65456 8756 65465
rect 8716 64709 8756 65416
rect 8523 64700 8565 64709
rect 8523 64660 8524 64700
rect 8564 64660 8565 64700
rect 8523 64651 8565 64660
rect 8715 64700 8757 64709
rect 8715 64660 8716 64700
rect 8756 64660 8757 64700
rect 8715 64651 8757 64660
rect 8524 64280 8564 64651
rect 8620 64616 8660 64627
rect 8620 64541 8660 64576
rect 8619 64532 8661 64541
rect 8619 64492 8620 64532
rect 8660 64492 8756 64532
rect 8619 64483 8661 64492
rect 8524 64240 8660 64280
rect 8523 64112 8565 64121
rect 8523 64072 8524 64112
rect 8564 64072 8565 64112
rect 8523 64063 8565 64072
rect 8524 63869 8564 64063
rect 8523 63860 8565 63869
rect 8523 63820 8524 63860
rect 8564 63820 8565 63860
rect 8523 63811 8565 63820
rect 8427 63524 8469 63533
rect 8427 63484 8428 63524
rect 8468 63484 8469 63524
rect 8427 63475 8469 63484
rect 8428 62684 8468 63475
rect 8620 63113 8660 64240
rect 8619 63104 8661 63113
rect 8619 63064 8620 63104
rect 8660 63064 8661 63104
rect 8619 63055 8661 63064
rect 8620 62970 8660 63055
rect 8428 62644 8564 62684
rect 8428 61601 8468 61686
rect 8427 61592 8469 61601
rect 8427 61552 8428 61592
rect 8468 61552 8469 61592
rect 8427 61543 8469 61552
rect 8427 61424 8469 61433
rect 8427 61384 8428 61424
rect 8468 61384 8469 61424
rect 8427 61375 8469 61384
rect 8428 56897 8468 61375
rect 8524 60593 8564 62644
rect 8619 62432 8661 62441
rect 8716 62432 8756 64492
rect 8812 64280 8852 70624
rect 9004 70614 9044 70699
rect 9196 70673 9236 74740
rect 9292 71513 9332 83467
rect 9387 83180 9429 83189
rect 9387 83140 9388 83180
rect 9428 83140 9429 83180
rect 9387 83131 9429 83140
rect 9291 71504 9333 71513
rect 9291 71464 9292 71504
rect 9332 71464 9333 71504
rect 9291 71455 9333 71464
rect 9388 71420 9428 83131
rect 9484 76880 9524 85936
rect 9579 83936 9621 83945
rect 9579 83896 9580 83936
rect 9620 83896 9621 83936
rect 9579 83887 9621 83896
rect 9580 79577 9620 83887
rect 9579 79568 9621 79577
rect 9579 79528 9580 79568
rect 9620 79528 9621 79568
rect 9579 79519 9621 79528
rect 9484 76840 9620 76880
rect 9483 76712 9525 76721
rect 9483 76672 9484 76712
rect 9524 76672 9525 76712
rect 9483 76663 9525 76672
rect 9484 76578 9524 76663
rect 9580 75788 9620 76840
rect 9484 75748 9620 75788
rect 9484 74537 9524 75748
rect 9579 75620 9621 75629
rect 9579 75580 9580 75620
rect 9620 75580 9621 75620
rect 9579 75571 9621 75580
rect 9483 74528 9525 74537
rect 9483 74488 9484 74528
rect 9524 74488 9525 74528
rect 9483 74479 9525 74488
rect 9580 74528 9620 75571
rect 9580 74479 9620 74488
rect 9676 73781 9716 85936
rect 9868 81920 9908 85936
rect 10060 84449 10100 85936
rect 10059 84440 10101 84449
rect 10059 84400 10060 84440
rect 10100 84400 10101 84440
rect 10059 84391 10101 84400
rect 10155 82340 10197 82349
rect 10155 82300 10156 82340
rect 10196 82300 10197 82340
rect 10155 82291 10197 82300
rect 9868 81880 10004 81920
rect 9771 79232 9813 79241
rect 9771 79192 9772 79232
rect 9812 79192 9813 79232
rect 9771 79183 9813 79192
rect 9675 73772 9717 73781
rect 9675 73732 9676 73772
rect 9716 73732 9717 73772
rect 9675 73723 9717 73732
rect 9579 73688 9621 73697
rect 9579 73648 9580 73688
rect 9620 73648 9621 73688
rect 9579 73639 9621 73648
rect 9580 73554 9620 73639
rect 9675 71588 9717 71597
rect 9675 71548 9676 71588
rect 9716 71548 9717 71588
rect 9675 71539 9717 71548
rect 9484 71420 9524 71429
rect 9388 71380 9484 71420
rect 9195 70664 9237 70673
rect 9195 70624 9196 70664
rect 9236 70624 9237 70664
rect 9195 70615 9237 70624
rect 9003 70496 9045 70505
rect 9003 70456 9004 70496
rect 9044 70456 9045 70496
rect 9003 70447 9045 70456
rect 8907 70412 8949 70421
rect 8907 70372 8908 70412
rect 8948 70372 8949 70412
rect 8907 70363 8949 70372
rect 8908 69152 8948 70363
rect 8908 66128 8948 69112
rect 9004 68321 9044 70447
rect 9484 69572 9524 71380
rect 9580 71420 9620 71429
rect 9580 70757 9620 71380
rect 9579 70748 9621 70757
rect 9579 70708 9580 70748
rect 9620 70708 9621 70748
rect 9579 70699 9621 70708
rect 9676 70673 9716 71539
rect 9675 70664 9717 70673
rect 9675 70624 9676 70664
rect 9716 70624 9717 70664
rect 9675 70615 9717 70624
rect 9676 69992 9716 70615
rect 9484 69532 9620 69572
rect 9195 69152 9237 69161
rect 9195 69112 9196 69152
rect 9236 69112 9237 69152
rect 9195 69103 9237 69112
rect 9003 68312 9045 68321
rect 9003 68272 9004 68312
rect 9044 68272 9045 68312
rect 9003 68263 9045 68272
rect 9004 66968 9044 68263
rect 9099 67892 9141 67901
rect 9099 67852 9100 67892
rect 9140 67852 9141 67892
rect 9099 67843 9141 67852
rect 9100 67733 9140 67843
rect 9099 67724 9141 67733
rect 9099 67684 9100 67724
rect 9140 67684 9141 67724
rect 9099 67675 9141 67684
rect 9100 67640 9140 67675
rect 9100 67589 9140 67600
rect 9004 66919 9044 66928
rect 9099 66128 9141 66137
rect 8908 66088 9100 66128
rect 9140 66088 9141 66128
rect 9099 66079 9141 66088
rect 9100 65994 9140 66079
rect 9100 65456 9140 65467
rect 9100 65381 9140 65416
rect 9099 65372 9141 65381
rect 9099 65332 9100 65372
rect 9140 65332 9141 65372
rect 9099 65323 9141 65332
rect 8908 65204 8948 65213
rect 8948 65164 9140 65204
rect 8908 65155 8948 65164
rect 9100 64630 9140 65164
rect 9100 64581 9140 64590
rect 8812 64240 8948 64280
rect 8811 63272 8853 63281
rect 8811 63232 8812 63272
rect 8852 63232 8853 63272
rect 8811 63223 8853 63232
rect 8812 63138 8852 63223
rect 8908 62852 8948 64240
rect 9100 63944 9140 63953
rect 9100 63701 9140 63904
rect 9099 63692 9141 63701
rect 9099 63652 9100 63692
rect 9140 63652 9141 63692
rect 9099 63643 9141 63652
rect 9099 63272 9141 63281
rect 9099 63232 9100 63272
rect 9140 63232 9141 63272
rect 9099 63223 9141 63232
rect 9003 63188 9045 63197
rect 9003 63148 9004 63188
rect 9044 63148 9045 63188
rect 9003 63139 9045 63148
rect 9004 63104 9044 63139
rect 9004 63053 9044 63064
rect 8908 62812 9044 62852
rect 8811 62768 8853 62777
rect 8811 62728 8812 62768
rect 8852 62728 8853 62768
rect 8811 62719 8853 62728
rect 8619 62392 8620 62432
rect 8660 62392 8756 62432
rect 8619 62383 8661 62392
rect 8620 62298 8660 62383
rect 8812 61592 8852 62719
rect 8907 61760 8949 61769
rect 8907 61720 8908 61760
rect 8948 61720 8949 61760
rect 8907 61711 8949 61720
rect 8812 61543 8852 61552
rect 8620 61424 8660 61433
rect 8660 61384 8756 61424
rect 8620 61375 8660 61384
rect 8716 60915 8756 61384
rect 8908 61088 8948 61711
rect 8908 61039 8948 61048
rect 8716 60866 8756 60875
rect 9004 60845 9044 62812
rect 9100 62427 9140 63223
rect 9100 62378 9140 62387
rect 9100 60920 9140 60929
rect 9196 60920 9236 69103
rect 9483 68480 9525 68489
rect 9483 68440 9484 68480
rect 9524 68440 9525 68480
rect 9483 68431 9525 68440
rect 9484 67733 9524 68431
rect 9483 67724 9525 67733
rect 9483 67684 9484 67724
rect 9524 67684 9525 67724
rect 9483 67675 9525 67684
rect 9292 67472 9332 67481
rect 9332 67432 9524 67472
rect 9292 67423 9332 67432
rect 9484 66963 9524 67432
rect 9484 66914 9524 66923
rect 9387 66128 9429 66137
rect 9387 66088 9388 66128
rect 9428 66088 9429 66128
rect 9387 66079 9429 66088
rect 9291 64448 9333 64457
rect 9291 64408 9292 64448
rect 9332 64408 9333 64448
rect 9291 64399 9333 64408
rect 9292 64314 9332 64399
rect 9291 62684 9333 62693
rect 9291 62644 9292 62684
rect 9332 62644 9333 62684
rect 9291 62635 9333 62644
rect 9292 62600 9332 62635
rect 9292 62549 9332 62560
rect 9140 60880 9236 60920
rect 9003 60836 9045 60845
rect 9003 60796 9004 60836
rect 9044 60796 9045 60836
rect 9003 60787 9045 60796
rect 9003 60668 9045 60677
rect 9003 60628 9004 60668
rect 9044 60628 9045 60668
rect 9003 60619 9045 60628
rect 8523 60584 8565 60593
rect 8523 60544 8524 60584
rect 8564 60544 8565 60584
rect 8523 60535 8565 60544
rect 9004 59408 9044 60619
rect 9100 59912 9140 60880
rect 9195 60248 9237 60257
rect 9195 60208 9196 60248
rect 9236 60208 9237 60248
rect 9195 60199 9237 60208
rect 9196 60080 9236 60199
rect 9196 60031 9236 60040
rect 9100 59872 9236 59912
rect 9100 59408 9140 59417
rect 9004 59368 9100 59408
rect 8811 59240 8853 59249
rect 8811 59200 8812 59240
rect 8852 59200 8853 59240
rect 8811 59191 8853 59200
rect 8619 59156 8661 59165
rect 8619 59116 8620 59156
rect 8660 59116 8661 59156
rect 8619 59107 8661 59116
rect 8620 58568 8660 59107
rect 8620 57149 8660 58528
rect 8812 57896 8852 59191
rect 9100 58997 9140 59368
rect 9099 58988 9141 58997
rect 9099 58948 9100 58988
rect 9140 58948 9141 58988
rect 9099 58939 9141 58948
rect 9100 58573 9140 58582
rect 9004 58064 9044 58073
rect 9100 58064 9140 58533
rect 9044 58024 9140 58064
rect 9004 58015 9044 58024
rect 8812 57847 8852 57856
rect 9099 57896 9141 57905
rect 9099 57856 9100 57896
rect 9140 57856 9141 57896
rect 9099 57847 9141 57856
rect 8619 57140 8661 57149
rect 8619 57100 8620 57140
rect 8660 57100 8661 57140
rect 8619 57091 8661 57100
rect 8811 57056 8853 57065
rect 8811 57016 8812 57056
rect 8852 57016 8853 57056
rect 8811 57007 8853 57016
rect 9100 57056 9140 57847
rect 8427 56888 8469 56897
rect 8427 56848 8428 56888
rect 8468 56848 8469 56888
rect 8427 56839 8469 56848
rect 8236 56596 8372 56636
rect 8236 56393 8276 56596
rect 8332 56512 8756 56552
rect 8235 56384 8277 56393
rect 8235 56344 8236 56384
rect 8276 56344 8277 56384
rect 8235 56335 8277 56344
rect 8236 56216 8276 56225
rect 8332 56216 8372 56512
rect 8428 56384 8468 56393
rect 8620 56384 8660 56393
rect 8468 56344 8564 56384
rect 8428 56335 8468 56344
rect 8276 56176 8372 56216
rect 8427 56216 8469 56225
rect 8427 56176 8428 56216
rect 8468 56176 8469 56216
rect 8236 56167 8276 56176
rect 8427 56167 8469 56176
rect 8428 56082 8468 56167
rect 8140 56008 8276 56048
rect 8139 55796 8181 55805
rect 8139 55756 8140 55796
rect 8180 55756 8181 55796
rect 8139 55747 8181 55756
rect 8140 55544 8180 55747
rect 8140 55495 8180 55504
rect 8236 55544 8276 56008
rect 8331 55712 8373 55721
rect 8331 55672 8332 55712
rect 8372 55672 8373 55712
rect 8331 55663 8373 55672
rect 8236 55495 8276 55504
rect 8332 55544 8372 55663
rect 8332 55495 8372 55504
rect 8428 55544 8468 55553
rect 8524 55544 8564 56344
rect 8620 55805 8660 56344
rect 8716 56384 8756 56512
rect 8716 56335 8756 56344
rect 8812 56216 8852 57007
rect 9100 56813 9140 57016
rect 9099 56804 9141 56813
rect 9099 56764 9100 56804
rect 9140 56764 9141 56804
rect 9099 56755 9141 56764
rect 8908 56393 8948 56478
rect 8907 56384 8949 56393
rect 8907 56344 8908 56384
rect 8948 56344 8949 56384
rect 8907 56335 8949 56344
rect 9100 56384 9140 56393
rect 8908 56216 8948 56225
rect 8812 56176 8908 56216
rect 8908 56167 8948 56176
rect 8619 55796 8661 55805
rect 8619 55756 8620 55796
rect 8660 55756 8661 55796
rect 8619 55747 8661 55756
rect 9100 55721 9140 56344
rect 9099 55712 9141 55721
rect 9099 55672 9100 55712
rect 9140 55672 9141 55712
rect 9099 55663 9141 55672
rect 8619 55628 8661 55637
rect 8619 55588 8620 55628
rect 8660 55588 8661 55628
rect 8619 55579 8661 55588
rect 8468 55504 8564 55544
rect 8620 55544 8660 55579
rect 8428 55495 8468 55504
rect 8620 55493 8660 55504
rect 7948 55411 7988 55420
rect 8236 54872 8276 54881
rect 8236 54788 8276 54832
rect 9003 54872 9045 54881
rect 9003 54832 9004 54872
rect 9044 54832 9045 54872
rect 9003 54823 9045 54832
rect 8331 54788 8373 54797
rect 8236 54748 8332 54788
rect 8372 54748 8373 54788
rect 8331 54739 8373 54748
rect 8139 54704 8181 54713
rect 8139 54664 8140 54704
rect 8180 54664 8181 54704
rect 8139 54655 8181 54664
rect 7756 54412 7892 54452
rect 7756 53621 7796 54412
rect 7851 54284 7893 54293
rect 7851 54244 7852 54284
rect 7892 54244 7893 54284
rect 7851 54235 7893 54244
rect 7755 53612 7797 53621
rect 7755 53572 7756 53612
rect 7796 53572 7797 53612
rect 7755 53563 7797 53572
rect 7659 53444 7701 53453
rect 7659 53404 7660 53444
rect 7700 53404 7701 53444
rect 7659 53395 7701 53404
rect 7660 53360 7700 53395
rect 7660 53309 7700 53320
rect 7755 53360 7797 53369
rect 7755 53320 7756 53360
rect 7796 53320 7797 53360
rect 7755 53311 7797 53320
rect 7756 53226 7796 53311
rect 7852 53108 7892 54235
rect 7947 54032 7989 54041
rect 7947 53992 7948 54032
rect 7988 53992 7989 54032
rect 7947 53983 7989 53992
rect 7948 53285 7988 53983
rect 8044 53528 8084 53537
rect 7947 53276 7989 53285
rect 7947 53236 7948 53276
rect 7988 53236 7989 53276
rect 7947 53227 7989 53236
rect 7660 53068 7892 53108
rect 7563 51260 7605 51269
rect 7563 51220 7564 51260
rect 7604 51220 7605 51260
rect 7563 51211 7605 51220
rect 7660 51185 7700 53068
rect 7755 52688 7797 52697
rect 7755 52648 7756 52688
rect 7796 52648 7797 52688
rect 7755 52639 7797 52648
rect 7756 52109 7796 52639
rect 7755 52100 7797 52109
rect 7755 52060 7756 52100
rect 7796 52060 7797 52100
rect 7755 52051 7797 52060
rect 7756 51848 7796 52051
rect 7756 51799 7796 51808
rect 7852 51764 7892 51773
rect 7852 51605 7892 51724
rect 7851 51596 7893 51605
rect 7851 51556 7852 51596
rect 7892 51556 7893 51596
rect 7851 51547 7893 51556
rect 7948 51353 7988 53227
rect 8044 52865 8084 53488
rect 8140 53108 8180 54655
rect 9004 54461 9044 54823
rect 9003 54452 9045 54461
rect 9003 54412 9004 54452
rect 9044 54412 9045 54452
rect 9003 54403 9045 54412
rect 8619 54200 8661 54209
rect 8619 54160 8620 54200
rect 8660 54160 8661 54200
rect 8619 54151 8661 54160
rect 8523 54032 8565 54041
rect 8523 53992 8524 54032
rect 8564 53992 8565 54032
rect 8523 53983 8565 53992
rect 8524 53898 8564 53983
rect 8427 53864 8469 53873
rect 8427 53824 8428 53864
rect 8468 53824 8469 53864
rect 8427 53815 8469 53824
rect 8235 53360 8277 53369
rect 8235 53320 8236 53360
rect 8276 53320 8277 53360
rect 8235 53311 8277 53320
rect 8332 53360 8372 53369
rect 8236 53226 8276 53311
rect 8332 53117 8372 53320
rect 8331 53108 8373 53117
rect 8140 53068 8276 53108
rect 8139 52940 8181 52949
rect 8139 52900 8140 52940
rect 8180 52900 8181 52940
rect 8139 52891 8181 52900
rect 8043 52856 8085 52865
rect 8043 52816 8044 52856
rect 8084 52816 8085 52856
rect 8043 52807 8085 52816
rect 8043 52604 8085 52613
rect 8043 52564 8044 52604
rect 8084 52564 8085 52604
rect 8043 52555 8085 52564
rect 7947 51344 7989 51353
rect 7947 51304 7948 51344
rect 7988 51304 7989 51344
rect 7947 51295 7989 51304
rect 8044 51269 8084 52555
rect 8140 52520 8180 52891
rect 8140 52471 8180 52480
rect 8236 52361 8276 53068
rect 8331 53068 8332 53108
rect 8372 53068 8373 53108
rect 8331 53059 8373 53068
rect 8331 52772 8373 52781
rect 8331 52732 8332 52772
rect 8372 52732 8373 52772
rect 8331 52723 8373 52732
rect 8332 52520 8372 52723
rect 8332 52471 8372 52480
rect 8235 52352 8277 52361
rect 8235 52312 8236 52352
rect 8276 52312 8277 52352
rect 8235 52303 8277 52312
rect 8236 51848 8276 51857
rect 8043 51260 8085 51269
rect 8043 51220 8044 51260
rect 8084 51220 8085 51260
rect 8043 51211 8085 51220
rect 7659 51176 7701 51185
rect 7659 51136 7660 51176
rect 7700 51136 7701 51176
rect 7659 51127 7701 51136
rect 8236 51092 8276 51808
rect 8331 51848 8373 51857
rect 8331 51808 8332 51848
rect 8372 51808 8373 51848
rect 8331 51799 8373 51808
rect 8332 51714 8372 51799
rect 8140 51052 8372 51092
rect 7467 51008 7509 51017
rect 7467 50968 7468 51008
rect 7508 50968 7509 51008
rect 7467 50959 7509 50968
rect 7564 51008 7604 51017
rect 8044 51008 8084 51019
rect 7604 50968 7700 51008
rect 7564 50959 7604 50968
rect 7468 50840 7508 50959
rect 7468 50800 7604 50840
rect 7467 50588 7509 50597
rect 7467 50548 7468 50588
rect 7508 50548 7509 50588
rect 7467 50539 7509 50548
rect 7372 50287 7412 50296
rect 7276 49748 7316 49757
rect 7180 49708 7276 49748
rect 7083 49699 7125 49708
rect 7276 49699 7316 49708
rect 7084 49614 7124 49699
rect 7468 49337 7508 50539
rect 7564 49496 7604 50800
rect 7660 50681 7700 50968
rect 8044 50933 8084 50968
rect 8140 51008 8180 51052
rect 8140 50959 8180 50968
rect 8332 50933 8372 51052
rect 7755 50924 7797 50933
rect 7755 50884 7756 50924
rect 7796 50884 7797 50924
rect 7755 50875 7797 50884
rect 8043 50924 8085 50933
rect 8043 50884 8044 50924
rect 8084 50884 8085 50924
rect 8043 50875 8085 50884
rect 8331 50924 8373 50933
rect 8331 50884 8332 50924
rect 8372 50884 8373 50924
rect 8331 50875 8373 50884
rect 7756 50790 7796 50875
rect 8235 50840 8277 50849
rect 8235 50800 8236 50840
rect 8276 50800 8277 50840
rect 8235 50791 8277 50800
rect 7659 50672 7701 50681
rect 7659 50632 7660 50672
rect 7700 50632 7701 50672
rect 7659 50623 7701 50632
rect 8236 50513 8276 50791
rect 8235 50504 8277 50513
rect 8235 50464 8236 50504
rect 8276 50464 8277 50504
rect 8235 50455 8277 50464
rect 7947 50420 7989 50429
rect 7947 50380 7948 50420
rect 7988 50380 7989 50420
rect 7947 50371 7989 50380
rect 7660 50291 7700 50347
rect 7659 50212 7660 50261
rect 7756 50336 7796 50345
rect 7700 50212 7701 50261
rect 7659 50203 7701 50212
rect 7659 49664 7701 49673
rect 7659 49624 7660 49664
rect 7700 49624 7701 49664
rect 7659 49615 7701 49624
rect 7564 49447 7604 49456
rect 7660 49496 7700 49615
rect 7660 49447 7700 49456
rect 7467 49328 7509 49337
rect 7467 49288 7468 49328
rect 7508 49288 7509 49328
rect 7467 49279 7509 49288
rect 6987 48908 7029 48917
rect 6987 48868 6988 48908
rect 7028 48868 7029 48908
rect 6987 48859 7029 48868
rect 7468 48908 7508 48917
rect 7508 48868 7700 48908
rect 7468 48859 7508 48868
rect 6795 48824 6837 48833
rect 6795 48784 6796 48824
rect 6836 48784 6837 48824
rect 6795 48775 6837 48784
rect 7275 48824 7317 48833
rect 7275 48779 7276 48824
rect 7316 48779 7317 48824
rect 7275 48775 7317 48779
rect 7660 48824 7700 48868
rect 7660 48775 7700 48784
rect 6796 48690 6836 48775
rect 7276 48689 7316 48775
rect 7563 48740 7605 48749
rect 7563 48700 7564 48740
rect 7604 48700 7605 48740
rect 7563 48691 7605 48700
rect 7467 48656 7509 48665
rect 7467 48616 7468 48656
rect 7508 48616 7509 48656
rect 7467 48607 7509 48616
rect 7468 48413 7508 48607
rect 7467 48404 7509 48413
rect 7467 48364 7468 48404
rect 7508 48364 7509 48404
rect 7467 48355 7509 48364
rect 6987 48236 7029 48245
rect 6987 48196 6988 48236
rect 7028 48196 7029 48236
rect 6987 48187 7029 48196
rect 6796 48152 6836 48163
rect 6796 48077 6836 48112
rect 6795 48068 6837 48077
rect 6795 48028 6796 48068
rect 6836 48028 6837 48068
rect 6795 48019 6837 48028
rect 6891 47984 6933 47993
rect 6891 47944 6892 47984
rect 6932 47944 6933 47984
rect 6891 47935 6933 47944
rect 6988 47984 7028 48187
rect 7083 48068 7125 48077
rect 7083 48028 7084 48068
rect 7124 48028 7125 48068
rect 7083 48019 7125 48028
rect 6700 47860 6836 47900
rect 6603 47851 6645 47860
rect 6604 47312 6644 47321
rect 6604 46565 6644 47272
rect 6699 47312 6741 47321
rect 6699 47272 6700 47312
rect 6740 47272 6741 47312
rect 6699 47263 6741 47272
rect 6700 47178 6740 47263
rect 6796 47144 6836 47860
rect 6892 47312 6932 47935
rect 6988 47321 7028 47944
rect 7084 47984 7124 48019
rect 7084 47933 7124 47944
rect 7275 47984 7317 47993
rect 7275 47944 7276 47984
rect 7316 47944 7317 47984
rect 7275 47935 7317 47944
rect 7468 47984 7508 48355
rect 7564 48077 7604 48691
rect 7659 48656 7701 48665
rect 7659 48616 7660 48656
rect 7700 48616 7701 48656
rect 7659 48607 7701 48616
rect 7660 48522 7700 48607
rect 7563 48068 7605 48077
rect 7563 48028 7564 48068
rect 7604 48028 7605 48068
rect 7563 48019 7605 48028
rect 7468 47935 7508 47944
rect 7564 47984 7604 48019
rect 7276 47816 7316 47935
rect 7564 47934 7604 47944
rect 7659 47984 7701 47993
rect 7659 47944 7660 47984
rect 7700 47944 7701 47984
rect 7659 47935 7701 47944
rect 7756 47984 7796 50296
rect 7852 50336 7892 50345
rect 7852 49757 7892 50296
rect 7948 50286 7988 50371
rect 8236 50336 8276 50455
rect 8236 50287 8276 50296
rect 8235 49832 8277 49841
rect 8235 49792 8236 49832
rect 8276 49792 8277 49832
rect 8235 49783 8277 49792
rect 7851 49748 7893 49757
rect 7851 49708 7852 49748
rect 7892 49708 7893 49748
rect 7851 49699 7893 49708
rect 8236 49748 8276 49783
rect 7852 48824 7892 49699
rect 8236 49697 8276 49708
rect 8428 49673 8468 53815
rect 8523 53528 8565 53537
rect 8523 53488 8524 53528
rect 8564 53488 8565 53528
rect 8523 53479 8565 53488
rect 8524 53360 8564 53479
rect 8620 53369 8660 54151
rect 9099 54116 9141 54125
rect 9099 54076 9100 54116
rect 9140 54076 9141 54116
rect 9099 54067 9141 54076
rect 8715 54032 8757 54041
rect 8715 53992 8716 54032
rect 8756 53992 8757 54032
rect 8715 53983 8757 53992
rect 9003 54032 9045 54041
rect 9003 53992 9004 54032
rect 9044 53992 9045 54032
rect 9003 53983 9045 53992
rect 9100 54032 9140 54067
rect 8716 53948 8756 53983
rect 8716 53897 8756 53908
rect 9004 53864 9044 53983
rect 9100 53981 9140 53992
rect 9004 53824 9140 53864
rect 8907 53612 8949 53621
rect 8907 53572 8908 53612
rect 8948 53572 8949 53612
rect 8907 53563 8949 53572
rect 8812 53528 8852 53537
rect 8716 53488 8812 53528
rect 8524 53311 8564 53320
rect 8619 53360 8661 53369
rect 8619 53320 8620 53360
rect 8660 53320 8661 53360
rect 8619 53311 8661 53320
rect 8620 53226 8660 53311
rect 8619 53108 8661 53117
rect 8619 53068 8620 53108
rect 8660 53068 8661 53108
rect 8619 53059 8661 53068
rect 8523 51596 8565 51605
rect 8523 51556 8524 51596
rect 8564 51556 8565 51596
rect 8523 51547 8565 51556
rect 8524 51008 8564 51547
rect 8620 51512 8660 53059
rect 8716 52529 8756 53488
rect 8812 53479 8852 53488
rect 8715 52520 8757 52529
rect 8715 52480 8716 52520
rect 8756 52480 8757 52520
rect 8715 52471 8757 52480
rect 8620 51472 8852 51512
rect 8619 51344 8661 51353
rect 8619 51304 8620 51344
rect 8660 51304 8661 51344
rect 8619 51295 8661 51304
rect 8620 51185 8660 51295
rect 8619 51176 8661 51185
rect 8619 51136 8620 51176
rect 8660 51136 8661 51176
rect 8619 51127 8661 51136
rect 8620 51092 8660 51127
rect 8812 51092 8852 51472
rect 8620 51041 8660 51052
rect 8716 51052 8852 51092
rect 8524 50924 8564 50968
rect 8524 50884 8660 50924
rect 8620 50009 8660 50884
rect 8619 50000 8661 50009
rect 8619 49960 8620 50000
rect 8660 49960 8661 50000
rect 8619 49951 8661 49960
rect 8427 49664 8469 49673
rect 8427 49624 8428 49664
rect 8468 49624 8469 49664
rect 8427 49615 8469 49624
rect 7948 49496 7988 49505
rect 7948 48833 7988 49456
rect 8236 49496 8276 49505
rect 7852 48775 7892 48784
rect 7947 48824 7989 48833
rect 7947 48784 7948 48824
rect 7988 48784 7989 48824
rect 7947 48775 7989 48784
rect 8044 48824 8084 48833
rect 8044 48581 8084 48784
rect 8236 48665 8276 49456
rect 8427 49496 8469 49505
rect 8427 49456 8428 49496
rect 8468 49456 8469 49496
rect 8427 49447 8469 49456
rect 8428 49362 8468 49447
rect 8235 48656 8277 48665
rect 8235 48616 8236 48656
rect 8276 48616 8277 48656
rect 8235 48607 8277 48616
rect 8043 48572 8085 48581
rect 8043 48532 8044 48572
rect 8084 48532 8085 48572
rect 8043 48523 8085 48532
rect 8619 48572 8661 48581
rect 8619 48532 8620 48572
rect 8660 48532 8661 48572
rect 8619 48523 8661 48532
rect 8139 48068 8181 48077
rect 8139 48028 8140 48068
rect 8180 48028 8181 48068
rect 8139 48019 8181 48028
rect 7756 47935 7796 47944
rect 7660 47850 7700 47935
rect 7276 47767 7316 47776
rect 6892 47263 6932 47272
rect 6987 47312 7029 47321
rect 6987 47272 6988 47312
rect 7028 47272 7029 47312
rect 6987 47263 7029 47272
rect 8140 47312 8180 48019
rect 8620 47984 8660 48523
rect 8620 47935 8660 47944
rect 8716 47480 8756 51052
rect 8716 47440 8852 47480
rect 6796 47104 7028 47144
rect 6699 46724 6741 46733
rect 6699 46684 6700 46724
rect 6740 46684 6741 46724
rect 6699 46675 6741 46684
rect 6603 46556 6645 46565
rect 6603 46516 6604 46556
rect 6644 46516 6645 46556
rect 6603 46507 6645 46516
rect 6604 46397 6644 46507
rect 6700 46472 6740 46675
rect 6988 46640 7028 47104
rect 7563 46724 7605 46733
rect 7563 46684 7564 46724
rect 7604 46684 7605 46724
rect 7563 46675 7605 46684
rect 7083 46640 7125 46649
rect 6988 46600 7084 46640
rect 7124 46600 7125 46640
rect 7083 46591 7125 46600
rect 7276 46565 7316 46609
rect 7275 46556 7317 46565
rect 7275 46516 7276 46556
rect 7316 46516 7317 46556
rect 7275 46514 7317 46516
rect 7275 46507 7276 46514
rect 7084 46472 7124 46481
rect 6700 46423 6740 46432
rect 6796 46432 7084 46472
rect 6603 46388 6645 46397
rect 6603 46348 6604 46388
rect 6644 46348 6645 46388
rect 6603 46339 6645 46348
rect 6796 46313 6836 46432
rect 7084 46423 7124 46432
rect 7179 46472 7221 46481
rect 7179 46432 7180 46472
rect 7220 46432 7221 46472
rect 7316 46507 7317 46514
rect 7276 46465 7316 46474
rect 7179 46423 7221 46432
rect 7180 46338 7220 46423
rect 6795 46304 6837 46313
rect 6795 46264 6796 46304
rect 6836 46264 6837 46304
rect 6795 46255 6837 46264
rect 6892 46304 6932 46313
rect 7372 46304 7412 46313
rect 6932 46264 7124 46304
rect 6892 46255 6932 46264
rect 6604 46238 6644 46247
rect 6603 46180 6604 46229
rect 6644 46180 6645 46229
rect 6603 46171 6645 46180
rect 6604 46103 6644 46171
rect 6987 46136 7029 46145
rect 6987 46096 6988 46136
rect 7028 46096 7029 46136
rect 6987 46087 7029 46096
rect 6892 45800 6932 45809
rect 6508 45760 6892 45800
rect 6315 45632 6357 45641
rect 6315 45592 6316 45632
rect 6356 45592 6357 45632
rect 6315 45583 6357 45592
rect 6316 44456 6356 45583
rect 6412 45557 6452 45760
rect 6892 45751 6932 45760
rect 6699 45632 6741 45641
rect 6699 45592 6700 45632
rect 6740 45592 6741 45632
rect 6699 45583 6741 45592
rect 6411 45548 6453 45557
rect 6411 45508 6412 45548
rect 6452 45508 6453 45548
rect 6411 45499 6453 45508
rect 6507 44960 6549 44969
rect 6507 44920 6508 44960
rect 6548 44920 6549 44960
rect 6507 44911 6549 44920
rect 6316 44407 6356 44416
rect 6508 44297 6548 44911
rect 6507 44288 6549 44297
rect 6507 44248 6508 44288
rect 6548 44248 6549 44288
rect 6507 44239 6549 44248
rect 6508 43541 6548 44239
rect 6700 43700 6740 45583
rect 6988 45557 7028 46087
rect 6987 45548 7029 45557
rect 6987 45508 6988 45548
rect 7028 45508 7029 45548
rect 6987 45499 7029 45508
rect 6891 45464 6933 45473
rect 6891 45424 6892 45464
rect 6932 45424 6933 45464
rect 6891 45415 6933 45424
rect 6795 44960 6837 44969
rect 6795 44920 6796 44960
rect 6836 44920 6837 44960
rect 6795 44911 6837 44920
rect 6796 44826 6836 44911
rect 6892 44540 6932 45415
rect 6988 45212 7028 45499
rect 6988 45163 7028 45172
rect 7084 44792 7124 46264
rect 7372 45884 7412 46264
rect 7564 46304 7604 46675
rect 8140 46649 8180 47272
rect 8620 47312 8660 47321
rect 8332 47144 8372 47153
rect 8620 47144 8660 47272
rect 8715 47312 8757 47321
rect 8715 47272 8716 47312
rect 8756 47272 8757 47312
rect 8715 47263 8757 47272
rect 8716 47178 8756 47263
rect 8372 47104 8660 47144
rect 8332 47095 8372 47104
rect 8812 46901 8852 47440
rect 8811 46892 8853 46901
rect 8811 46852 8812 46892
rect 8852 46852 8853 46892
rect 8811 46843 8853 46852
rect 8619 46724 8661 46733
rect 8619 46684 8620 46724
rect 8660 46684 8661 46724
rect 8619 46675 8661 46684
rect 8139 46640 8181 46649
rect 8139 46600 8140 46640
rect 8180 46600 8181 46640
rect 8139 46591 8181 46600
rect 8236 46565 8276 46596
rect 8235 46556 8277 46565
rect 8235 46516 8236 46556
rect 8276 46516 8277 46556
rect 8235 46507 8277 46516
rect 7756 46472 7796 46483
rect 7756 46397 7796 46432
rect 7851 46472 7893 46481
rect 8044 46472 8084 46481
rect 7851 46432 7852 46472
rect 7892 46432 7893 46472
rect 7851 46423 7893 46432
rect 7948 46432 8044 46472
rect 7755 46388 7797 46397
rect 7755 46348 7756 46388
rect 7796 46348 7797 46388
rect 7755 46339 7797 46348
rect 7852 46338 7892 46423
rect 7564 46255 7604 46264
rect 7948 45968 7988 46432
rect 8044 46423 8084 46432
rect 8236 46472 8276 46507
rect 8140 46304 8180 46313
rect 7756 45928 7988 45968
rect 8044 46264 8140 46304
rect 7564 45884 7604 45895
rect 7372 45844 7508 45884
rect 7372 45786 7412 45795
rect 7372 45557 7412 45746
rect 7179 45548 7221 45557
rect 7179 45508 7180 45548
rect 7220 45508 7221 45548
rect 7179 45499 7221 45508
rect 7371 45548 7413 45557
rect 7371 45508 7372 45548
rect 7412 45508 7413 45548
rect 7371 45499 7413 45508
rect 7180 44960 7220 45499
rect 7275 45212 7317 45221
rect 7275 45172 7276 45212
rect 7316 45172 7317 45212
rect 7275 45163 7317 45172
rect 7180 44911 7220 44920
rect 7276 44960 7316 45163
rect 7468 45137 7508 45844
rect 7564 45809 7604 45844
rect 7756 45809 7796 45928
rect 7563 45800 7605 45809
rect 7563 45760 7564 45800
rect 7604 45760 7605 45800
rect 7563 45751 7605 45760
rect 7755 45800 7797 45809
rect 7755 45760 7756 45800
rect 7796 45760 7797 45800
rect 7755 45751 7797 45760
rect 7947 45800 7989 45809
rect 7947 45760 7948 45800
rect 7988 45760 7989 45800
rect 7947 45751 7989 45760
rect 7948 45666 7988 45751
rect 7467 45128 7509 45137
rect 7467 45088 7468 45128
rect 7508 45088 7509 45128
rect 7467 45079 7509 45088
rect 7276 44911 7316 44920
rect 7372 44960 7412 44969
rect 7372 44792 7412 44920
rect 7468 44960 7508 44969
rect 7660 44960 7700 44969
rect 7508 44920 7660 44960
rect 7468 44911 7508 44920
rect 7660 44911 7700 44920
rect 7755 44960 7797 44969
rect 7755 44920 7756 44960
rect 7796 44920 7797 44960
rect 7755 44911 7797 44920
rect 7948 44960 7988 44969
rect 8044 44960 8084 46264
rect 8140 46255 8180 46264
rect 8236 45641 8276 46432
rect 8428 46472 8468 46481
rect 8428 46313 8468 46432
rect 8427 46304 8469 46313
rect 8427 46264 8428 46304
rect 8468 46264 8469 46304
rect 8427 46255 8469 46264
rect 8523 45800 8565 45809
rect 8523 45760 8524 45800
rect 8564 45760 8565 45800
rect 8523 45751 8565 45760
rect 8235 45632 8277 45641
rect 8235 45592 8236 45632
rect 8276 45592 8277 45632
rect 8235 45583 8277 45592
rect 8139 45128 8181 45137
rect 8139 45088 8140 45128
rect 8180 45088 8181 45128
rect 8139 45079 8181 45088
rect 8331 45128 8373 45137
rect 8331 45088 8332 45128
rect 8372 45088 8373 45128
rect 8331 45079 8373 45088
rect 7988 44920 8084 44960
rect 8140 44960 8180 45079
rect 7948 44911 7988 44920
rect 8140 44911 8180 44920
rect 8235 44960 8277 44969
rect 8235 44920 8236 44960
rect 8276 44920 8277 44960
rect 8235 44911 8277 44920
rect 7756 44826 7796 44911
rect 8236 44826 8276 44911
rect 7084 44752 7412 44792
rect 7851 44792 7893 44801
rect 7851 44752 7852 44792
rect 7892 44752 7893 44792
rect 7851 44743 7893 44752
rect 8043 44792 8085 44801
rect 8043 44752 8044 44792
rect 8084 44752 8085 44792
rect 8043 44743 8085 44752
rect 7467 44708 7509 44717
rect 7467 44668 7468 44708
rect 7508 44668 7509 44708
rect 7467 44659 7509 44668
rect 6892 44500 7028 44540
rect 6891 44372 6933 44381
rect 6891 44332 6892 44372
rect 6932 44332 6933 44372
rect 6891 44323 6933 44332
rect 6892 44288 6932 44323
rect 6892 44213 6932 44248
rect 6891 44204 6933 44213
rect 6891 44164 6892 44204
rect 6932 44164 6933 44204
rect 6891 44155 6933 44164
rect 6795 44120 6837 44129
rect 6892 44124 6932 44155
rect 6795 44080 6796 44120
rect 6836 44080 6837 44120
rect 6795 44071 6837 44080
rect 6700 43651 6740 43660
rect 6507 43532 6549 43541
rect 6507 43492 6508 43532
rect 6548 43492 6549 43532
rect 6507 43483 6549 43492
rect 6219 43448 6261 43457
rect 6219 43408 6220 43448
rect 6260 43408 6261 43448
rect 6219 43399 6261 43408
rect 6508 43448 6548 43483
rect 6796 43448 6836 44071
rect 6892 43448 6932 43457
rect 6796 43408 6892 43448
rect 6028 41896 6164 41936
rect 5932 41768 5972 41777
rect 5972 41728 6068 41768
rect 5932 41719 5972 41728
rect 5931 41600 5973 41609
rect 5931 41560 5932 41600
rect 5972 41560 5973 41600
rect 5931 41551 5973 41560
rect 5835 38156 5877 38165
rect 5835 38116 5836 38156
rect 5876 38116 5877 38156
rect 5835 38107 5877 38116
rect 5548 37780 5876 37820
rect 5547 37652 5589 37661
rect 5547 37612 5548 37652
rect 5588 37612 5589 37652
rect 5547 37603 5589 37612
rect 5548 37518 5588 37603
rect 5740 37400 5780 37409
rect 5740 37157 5780 37360
rect 5739 37148 5781 37157
rect 5739 37108 5740 37148
rect 5780 37108 5781 37148
rect 5739 37099 5781 37108
rect 5547 36980 5589 36989
rect 5547 36940 5548 36980
rect 5588 36940 5589 36980
rect 5547 36931 5589 36940
rect 5548 36728 5588 36931
rect 5548 36679 5588 36688
rect 5300 35848 5780 35888
rect 5260 35839 5300 35848
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 4780 35167 4820 35176
rect 5068 35216 5108 35225
rect 5260 35216 5300 35225
rect 5452 35216 5492 35225
rect 5108 35176 5204 35216
rect 5068 35167 5108 35176
rect 5164 35048 5204 35176
rect 5300 35176 5396 35216
rect 5260 35167 5300 35176
rect 5260 35048 5300 35057
rect 5164 35008 5260 35048
rect 5260 34999 5300 35008
rect 5067 34964 5109 34973
rect 5067 34924 5068 34964
rect 5108 34924 5109 34964
rect 5067 34915 5109 34924
rect 5068 34830 5108 34915
rect 5259 34712 5301 34721
rect 5259 34672 5260 34712
rect 5300 34672 5301 34712
rect 5259 34663 5301 34672
rect 5260 34469 5300 34663
rect 5259 34460 5301 34469
rect 5259 34420 5260 34460
rect 5300 34420 5301 34460
rect 5259 34411 5301 34420
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 5260 33872 5300 33881
rect 5356 33872 5396 35176
rect 5452 35048 5492 35176
rect 5548 35216 5588 35225
rect 5588 35176 5684 35216
rect 5548 35167 5588 35176
rect 5452 35008 5588 35048
rect 5451 34880 5493 34889
rect 5451 34840 5452 34880
rect 5492 34840 5493 34880
rect 5451 34831 5493 34840
rect 5452 33965 5492 34831
rect 5548 34217 5588 35008
rect 5547 34208 5589 34217
rect 5547 34168 5548 34208
rect 5588 34168 5589 34208
rect 5547 34159 5589 34168
rect 5451 33956 5493 33965
rect 5451 33916 5452 33956
rect 5492 33916 5493 33956
rect 5451 33907 5493 33916
rect 5300 33832 5396 33872
rect 5260 33823 5300 33832
rect 5163 33788 5205 33797
rect 5163 33748 5164 33788
rect 5204 33748 5205 33788
rect 5163 33739 5205 33748
rect 4876 33704 4916 33713
rect 4876 33545 4916 33664
rect 4972 33704 5012 33713
rect 4875 33536 4917 33545
rect 4875 33496 4876 33536
rect 4916 33496 4917 33536
rect 4875 33487 4917 33496
rect 4876 33125 4916 33487
rect 4972 33293 5012 33664
rect 5164 33694 5204 33739
rect 5356 33704 5396 33713
rect 5164 33664 5356 33694
rect 5164 33654 5396 33664
rect 5452 33704 5492 33713
rect 5452 33461 5492 33664
rect 5548 33704 5588 34159
rect 5644 34049 5684 35176
rect 5740 34553 5780 35848
rect 5836 35393 5876 37780
rect 5932 37745 5972 41551
rect 6028 40433 6068 41728
rect 6027 40424 6069 40433
rect 6027 40384 6028 40424
rect 6068 40384 6069 40424
rect 6027 40375 6069 40384
rect 6124 40181 6164 41896
rect 6220 41441 6260 43399
rect 6508 43397 6548 43408
rect 6892 43399 6932 43408
rect 6603 42776 6645 42785
rect 6603 42736 6604 42776
rect 6644 42736 6645 42776
rect 6603 42727 6645 42736
rect 6796 42776 6836 42785
rect 6604 42533 6644 42727
rect 6603 42524 6645 42533
rect 6603 42484 6604 42524
rect 6644 42484 6645 42524
rect 6603 42475 6645 42484
rect 6699 42356 6741 42365
rect 6699 42316 6700 42356
rect 6740 42316 6741 42356
rect 6699 42307 6741 42316
rect 6700 41609 6740 42307
rect 6315 41600 6357 41609
rect 6315 41560 6316 41600
rect 6356 41560 6357 41600
rect 6315 41551 6357 41560
rect 6699 41600 6741 41609
rect 6699 41560 6700 41600
rect 6740 41560 6741 41600
rect 6699 41551 6741 41560
rect 6219 41432 6261 41441
rect 6219 41392 6220 41432
rect 6260 41392 6261 41432
rect 6219 41383 6261 41392
rect 6316 40508 6356 41551
rect 6700 41264 6740 41551
rect 6796 41525 6836 42736
rect 6891 41600 6933 41609
rect 6891 41560 6892 41600
rect 6932 41560 6933 41600
rect 6891 41551 6933 41560
rect 6795 41516 6837 41525
rect 6795 41476 6796 41516
rect 6836 41476 6837 41516
rect 6795 41467 6837 41476
rect 6796 41264 6836 41273
rect 6700 41224 6796 41264
rect 6796 41215 6836 41224
rect 6411 40928 6453 40937
rect 6411 40888 6412 40928
rect 6452 40888 6453 40928
rect 6411 40879 6453 40888
rect 6220 40468 6356 40508
rect 6123 40172 6165 40181
rect 6123 40132 6124 40172
rect 6164 40132 6165 40172
rect 6123 40123 6165 40132
rect 6220 39668 6260 40468
rect 6412 40424 6452 40879
rect 6795 40676 6837 40685
rect 6795 40636 6796 40676
rect 6836 40636 6837 40676
rect 6795 40627 6837 40636
rect 6412 40375 6452 40384
rect 6699 40424 6741 40433
rect 6699 40384 6700 40424
rect 6740 40384 6741 40424
rect 6699 40375 6741 40384
rect 6796 40424 6836 40627
rect 6796 40375 6836 40384
rect 6315 40340 6357 40349
rect 6315 40300 6316 40340
rect 6356 40300 6357 40340
rect 6315 40291 6357 40300
rect 6603 40340 6645 40349
rect 6603 40300 6604 40340
rect 6644 40300 6645 40340
rect 6603 40291 6645 40300
rect 6316 39752 6356 40291
rect 6604 40206 6644 40291
rect 6412 39752 6452 39761
rect 6316 39712 6412 39752
rect 6412 39703 6452 39712
rect 6508 39752 6548 39763
rect 6508 39677 6548 39712
rect 6507 39668 6549 39677
rect 6220 39628 6356 39668
rect 6123 39500 6165 39509
rect 6123 39460 6124 39500
rect 6164 39460 6165 39500
rect 6123 39451 6165 39460
rect 6027 39080 6069 39089
rect 6027 39040 6028 39080
rect 6068 39040 6069 39080
rect 6027 39031 6069 39040
rect 6028 38753 6068 39031
rect 6027 38744 6069 38753
rect 6027 38704 6028 38744
rect 6068 38704 6069 38744
rect 6027 38695 6069 38704
rect 5931 37736 5973 37745
rect 5931 37696 5932 37736
rect 5972 37696 5973 37736
rect 5931 37687 5973 37696
rect 5835 35384 5877 35393
rect 5835 35344 5836 35384
rect 5876 35344 5877 35384
rect 5835 35335 5877 35344
rect 5836 35216 5876 35225
rect 5836 34628 5876 35176
rect 5932 35216 5972 35225
rect 5932 34889 5972 35176
rect 5931 34880 5973 34889
rect 5931 34840 5932 34880
rect 5972 34840 5973 34880
rect 5931 34831 5973 34840
rect 5932 34628 5972 34637
rect 5836 34588 5932 34628
rect 5932 34579 5972 34588
rect 6028 34553 6068 38695
rect 6124 36653 6164 39451
rect 6316 39089 6356 39628
rect 6507 39628 6508 39668
rect 6548 39628 6549 39668
rect 6507 39619 6549 39628
rect 6700 39248 6740 40375
rect 6892 39752 6932 41551
rect 6988 39845 7028 44500
rect 7083 44288 7125 44297
rect 7083 44248 7084 44288
rect 7124 44248 7125 44288
rect 7083 44239 7125 44248
rect 6987 39836 7029 39845
rect 6987 39796 6988 39836
rect 7028 39796 7029 39836
rect 6987 39787 7029 39796
rect 6892 39703 6932 39712
rect 6988 39668 7028 39677
rect 6700 39208 6836 39248
rect 6315 39080 6357 39089
rect 6315 39040 6316 39080
rect 6356 39040 6357 39080
rect 6315 39031 6357 39040
rect 6699 38576 6741 38585
rect 6699 38536 6700 38576
rect 6740 38536 6741 38576
rect 6699 38527 6741 38536
rect 6603 38408 6645 38417
rect 6603 38368 6604 38408
rect 6644 38368 6645 38408
rect 6603 38359 6645 38368
rect 6220 38240 6260 38249
rect 6220 37661 6260 38200
rect 6315 38240 6357 38249
rect 6315 38200 6316 38240
rect 6356 38200 6357 38240
rect 6315 38191 6357 38200
rect 6316 38106 6356 38191
rect 6507 37904 6549 37913
rect 6507 37864 6508 37904
rect 6548 37864 6549 37904
rect 6507 37855 6549 37864
rect 6219 37652 6261 37661
rect 6219 37612 6220 37652
rect 6260 37612 6261 37652
rect 6219 37603 6261 37612
rect 6508 36989 6548 37855
rect 6507 36980 6549 36989
rect 6507 36940 6508 36980
rect 6548 36940 6549 36980
rect 6507 36931 6549 36940
rect 6123 36644 6165 36653
rect 6123 36604 6124 36644
rect 6164 36604 6165 36644
rect 6123 36595 6165 36604
rect 6124 34637 6164 36595
rect 6604 36056 6644 38359
rect 6700 38240 6740 38527
rect 6700 38081 6740 38200
rect 6796 38240 6836 39208
rect 6891 39164 6933 39173
rect 6891 39124 6892 39164
rect 6932 39124 6933 39164
rect 6891 39115 6933 39124
rect 6892 38912 6932 39115
rect 6988 39089 7028 39628
rect 6987 39080 7029 39089
rect 6987 39040 6988 39080
rect 7028 39040 7029 39080
rect 6987 39031 7029 39040
rect 6988 38912 7028 38921
rect 6892 38872 6988 38912
rect 6699 38072 6741 38081
rect 6699 38032 6700 38072
rect 6740 38032 6741 38072
rect 6699 38023 6741 38032
rect 6796 36905 6836 38200
rect 6988 37409 7028 38872
rect 6987 37400 7029 37409
rect 6987 37360 6988 37400
rect 7028 37360 7029 37400
rect 6987 37351 7029 37360
rect 6988 37266 7028 37351
rect 6795 36896 6837 36905
rect 6795 36856 6796 36896
rect 6836 36856 6837 36896
rect 6795 36847 6837 36856
rect 7084 36737 7124 44239
rect 7468 44129 7508 44659
rect 7852 44658 7892 44743
rect 7467 44120 7509 44129
rect 7467 44080 7468 44120
rect 7508 44080 7509 44120
rect 7467 44071 7509 44080
rect 8044 43373 8084 44743
rect 8332 44708 8372 45079
rect 8236 44668 8372 44708
rect 8139 44288 8181 44297
rect 8139 44248 8140 44288
rect 8180 44248 8181 44288
rect 8139 44239 8181 44248
rect 8140 44154 8180 44239
rect 8236 44045 8276 44668
rect 8331 44540 8373 44549
rect 8331 44500 8332 44540
rect 8372 44500 8373 44540
rect 8331 44491 8373 44500
rect 8332 44456 8372 44491
rect 8332 44405 8372 44416
rect 8331 44120 8373 44129
rect 8331 44080 8332 44120
rect 8372 44080 8373 44120
rect 8331 44071 8373 44080
rect 8235 44036 8277 44045
rect 8235 43996 8236 44036
rect 8276 43996 8277 44036
rect 8235 43987 8277 43996
rect 8332 43868 8372 44071
rect 8524 43877 8564 45751
rect 8620 45137 8660 46675
rect 8715 45548 8757 45557
rect 8715 45508 8716 45548
rect 8756 45508 8757 45548
rect 8715 45499 8757 45508
rect 8716 45212 8756 45499
rect 8716 45172 8804 45212
rect 8619 45128 8661 45137
rect 8619 45088 8620 45128
rect 8660 45088 8661 45128
rect 8619 45079 8661 45088
rect 8764 45002 8804 45172
rect 8764 44953 8804 44962
rect 8619 44876 8661 44885
rect 8619 44836 8620 44876
rect 8660 44836 8661 44876
rect 8619 44827 8661 44836
rect 8620 44742 8660 44827
rect 8620 44288 8660 44297
rect 8236 43828 8372 43868
rect 8523 43868 8565 43877
rect 8523 43828 8524 43868
rect 8564 43828 8565 43868
rect 8139 43532 8181 43541
rect 8139 43492 8140 43532
rect 8180 43492 8181 43532
rect 8139 43483 8181 43492
rect 8140 43448 8180 43483
rect 8140 43397 8180 43408
rect 8043 43364 8085 43373
rect 8043 43324 8044 43364
rect 8084 43324 8085 43364
rect 8043 43315 8085 43324
rect 7371 43028 7413 43037
rect 7371 42988 7372 43028
rect 7412 42988 7413 43028
rect 7371 42979 7413 42988
rect 7372 41936 7412 42979
rect 7275 40592 7317 40601
rect 7275 40552 7276 40592
rect 7316 40552 7317 40592
rect 7275 40543 7317 40552
rect 7276 39332 7316 40543
rect 7372 39509 7412 41896
rect 8044 42776 8084 43315
rect 8044 41609 8084 42736
rect 8236 42692 8276 43828
rect 8523 43819 8565 43828
rect 8332 43700 8372 43709
rect 8620 43700 8660 44248
rect 8716 44288 8756 44297
rect 8756 44248 8852 44288
rect 8716 44239 8756 44248
rect 8715 44036 8757 44045
rect 8715 43996 8716 44036
rect 8756 43996 8757 44036
rect 8715 43987 8757 43996
rect 8372 43660 8660 43700
rect 8332 43651 8372 43660
rect 8716 43448 8756 43987
rect 8812 43793 8852 44248
rect 8811 43784 8853 43793
rect 8811 43744 8812 43784
rect 8852 43744 8853 43784
rect 8811 43735 8853 43744
rect 8716 43399 8756 43408
rect 8140 42652 8276 42692
rect 8140 41861 8180 42652
rect 8236 42524 8276 42533
rect 8276 42484 8564 42524
rect 8236 42475 8276 42484
rect 8139 41852 8181 41861
rect 8139 41812 8140 41852
rect 8180 41812 8181 41852
rect 8139 41803 8181 41812
rect 8043 41600 8085 41609
rect 8043 41560 8044 41600
rect 8084 41560 8085 41600
rect 8043 41551 8085 41560
rect 7659 41516 7701 41525
rect 7659 41476 7660 41516
rect 7700 41476 7701 41516
rect 7659 41467 7701 41476
rect 7563 41012 7605 41021
rect 7563 40972 7564 41012
rect 7604 40972 7605 41012
rect 7563 40963 7605 40972
rect 7564 40769 7604 40963
rect 7563 40760 7605 40769
rect 7563 40720 7564 40760
rect 7604 40720 7605 40760
rect 7563 40711 7605 40720
rect 7468 39752 7508 39761
rect 7371 39500 7413 39509
rect 7371 39460 7372 39500
rect 7412 39460 7413 39500
rect 7371 39451 7413 39460
rect 7276 39292 7412 39332
rect 7179 39080 7221 39089
rect 7179 39040 7180 39080
rect 7220 39040 7221 39080
rect 7179 39031 7221 39040
rect 7180 38946 7220 39031
rect 7372 38912 7412 39292
rect 7468 39257 7508 39712
rect 7467 39248 7509 39257
rect 7467 39208 7468 39248
rect 7508 39208 7509 39248
rect 7467 39199 7509 39208
rect 7564 39173 7604 40711
rect 7660 40517 7700 41467
rect 8044 41264 8084 41551
rect 8235 41348 8277 41357
rect 8235 41308 8236 41348
rect 8276 41308 8277 41348
rect 8235 41299 8277 41308
rect 8044 40937 8084 41224
rect 8236 41214 8276 41299
rect 8524 41264 8564 42484
rect 8620 41936 8660 41945
rect 8620 41609 8660 41896
rect 8811 41852 8853 41861
rect 8811 41812 8812 41852
rect 8852 41812 8853 41852
rect 8811 41803 8853 41812
rect 8812 41718 8852 41803
rect 8619 41600 8661 41609
rect 8619 41560 8620 41600
rect 8660 41560 8661 41600
rect 8619 41551 8661 41560
rect 8524 41215 8564 41224
rect 8619 41264 8661 41273
rect 8619 41224 8620 41264
rect 8660 41224 8661 41264
rect 8619 41215 8661 41224
rect 8043 40928 8085 40937
rect 8043 40888 8044 40928
rect 8084 40888 8085 40928
rect 8043 40879 8085 40888
rect 7659 40508 7701 40517
rect 7659 40468 7660 40508
rect 7700 40468 7701 40508
rect 7659 40459 7701 40468
rect 7563 39164 7605 39173
rect 7563 39124 7564 39164
rect 7604 39124 7605 39164
rect 7563 39115 7605 39124
rect 7467 38996 7509 39005
rect 7467 38956 7468 38996
rect 7508 38956 7509 38996
rect 7467 38947 7509 38956
rect 7372 38863 7412 38872
rect 7275 38408 7317 38417
rect 7275 38368 7276 38408
rect 7316 38368 7317 38408
rect 7275 38359 7317 38368
rect 7276 38240 7316 38359
rect 7276 38191 7316 38200
rect 7275 37988 7317 37997
rect 7275 37948 7276 37988
rect 7316 37948 7317 37988
rect 7275 37939 7317 37948
rect 7179 37652 7221 37661
rect 7179 37612 7180 37652
rect 7220 37612 7221 37652
rect 7179 37603 7221 37612
rect 7180 37518 7220 37603
rect 6795 36728 6837 36737
rect 6316 36016 6644 36056
rect 6700 36688 6796 36728
rect 6836 36688 6837 36728
rect 6219 35300 6261 35309
rect 6316 35300 6356 36016
rect 6508 35888 6548 35897
rect 6700 35888 6740 36688
rect 6795 36679 6837 36688
rect 7083 36728 7125 36737
rect 7083 36688 7084 36728
rect 7124 36688 7125 36728
rect 7083 36679 7125 36688
rect 6796 36594 6836 36679
rect 6987 36560 7029 36569
rect 6987 36520 6988 36560
rect 7028 36520 7029 36560
rect 6987 36511 7029 36520
rect 6988 36426 7028 36511
rect 7179 36140 7221 36149
rect 7179 36100 7180 36140
rect 7220 36100 7221 36140
rect 7179 36091 7221 36100
rect 7180 36006 7220 36091
rect 6548 35848 6740 35888
rect 6892 35888 6932 35897
rect 6508 35839 6548 35848
rect 6219 35260 6220 35300
rect 6260 35260 6356 35300
rect 6219 35251 6261 35260
rect 6316 35174 6356 35183
rect 6356 35134 6357 35174
rect 6316 35125 6357 35134
rect 6317 35048 6357 35125
rect 6316 35008 6357 35048
rect 6412 35132 6452 35141
rect 6412 35048 6452 35092
rect 6412 35008 6548 35048
rect 6316 34964 6356 35008
rect 6316 34924 6357 34964
rect 6317 34796 6357 34924
rect 6316 34756 6357 34796
rect 6123 34628 6165 34637
rect 6123 34588 6124 34628
rect 6164 34588 6165 34628
rect 6123 34579 6165 34588
rect 5739 34544 5781 34553
rect 5739 34504 5740 34544
rect 5780 34504 5781 34544
rect 5739 34495 5781 34504
rect 6027 34544 6069 34553
rect 6027 34504 6028 34544
rect 6068 34504 6069 34544
rect 6027 34495 6069 34504
rect 6123 34460 6165 34469
rect 6123 34420 6124 34460
rect 6164 34420 6165 34460
rect 6123 34411 6165 34420
rect 5739 34376 5781 34385
rect 5739 34336 5740 34376
rect 5780 34336 5781 34376
rect 5739 34327 5781 34336
rect 6124 34376 6164 34411
rect 5740 34242 5780 34327
rect 6124 34325 6164 34336
rect 5932 34208 5972 34217
rect 5932 34124 5972 34168
rect 5932 34084 6068 34124
rect 5643 34040 5685 34049
rect 5643 34000 5644 34040
rect 5684 34000 5685 34040
rect 6028 34040 6068 34084
rect 6028 34000 6164 34040
rect 5643 33991 5685 34000
rect 5931 33956 5973 33965
rect 5931 33916 5932 33956
rect 5972 33916 5973 33956
rect 5931 33907 5973 33916
rect 5836 33704 5876 33713
rect 5548 33655 5588 33664
rect 5740 33664 5836 33704
rect 5451 33452 5493 33461
rect 5451 33412 5452 33452
rect 5492 33412 5493 33452
rect 5451 33403 5493 33412
rect 5355 33368 5397 33377
rect 5355 33328 5356 33368
rect 5396 33328 5397 33368
rect 5355 33319 5397 33328
rect 4971 33284 5013 33293
rect 4971 33244 4972 33284
rect 5012 33244 5013 33284
rect 4971 33235 5013 33244
rect 4875 33116 4917 33125
rect 4875 33076 4876 33116
rect 4916 33076 4917 33116
rect 4875 33067 4917 33076
rect 4683 32948 4725 32957
rect 4683 32908 4684 32948
rect 4724 32908 4725 32948
rect 4683 32899 4725 32908
rect 5356 32864 5396 33319
rect 5548 33116 5588 33125
rect 5740 33116 5780 33664
rect 5836 33655 5876 33664
rect 5932 33704 5972 33907
rect 6124 33797 6164 34000
rect 6123 33788 6165 33797
rect 6123 33748 6124 33788
rect 6164 33748 6165 33788
rect 6123 33739 6165 33748
rect 5932 33545 5972 33664
rect 5931 33536 5973 33545
rect 5931 33496 5932 33536
rect 5972 33496 5973 33536
rect 5931 33487 5973 33496
rect 5588 33076 5780 33116
rect 5548 33067 5588 33076
rect 5740 32864 5780 32873
rect 5356 32815 5396 32824
rect 5644 32824 5740 32864
rect 4588 32740 4724 32780
rect 3916 32320 4244 32360
rect 3531 32152 3532 32192
rect 3572 32152 3668 32192
rect 4108 32192 4148 32201
rect 3531 32143 3573 32152
rect 3243 32108 3285 32117
rect 3243 32068 3244 32108
rect 3284 32068 3285 32108
rect 3243 32059 3285 32068
rect 3244 30512 3284 32059
rect 3436 31352 3476 31361
rect 3340 30689 3380 30774
rect 3436 30773 3476 31312
rect 3435 30764 3477 30773
rect 3435 30724 3436 30764
rect 3476 30724 3477 30764
rect 3435 30715 3477 30724
rect 3339 30680 3381 30689
rect 3339 30640 3340 30680
rect 3380 30640 3381 30680
rect 3339 30631 3381 30640
rect 3244 30472 3380 30512
rect 3148 30388 3284 30428
rect 3147 30008 3189 30017
rect 3147 29968 3148 30008
rect 3188 29968 3189 30008
rect 3147 29959 3189 29968
rect 3148 29849 3188 29959
rect 3147 29840 3189 29849
rect 3147 29800 3148 29840
rect 3188 29800 3189 29840
rect 3147 29791 3189 29800
rect 3244 29840 3284 30388
rect 3340 29924 3380 30472
rect 3436 30092 3476 30101
rect 3532 30092 3572 32143
rect 4108 31940 4148 32152
rect 4204 32108 4244 32320
rect 4340 32320 4436 32360
rect 4300 32311 4340 32320
rect 4492 32201 4532 32286
rect 4491 32192 4533 32201
rect 4491 32152 4492 32192
rect 4532 32152 4533 32192
rect 4491 32143 4533 32152
rect 4588 32192 4628 32203
rect 4588 32117 4628 32152
rect 4587 32108 4629 32117
rect 4204 32068 4436 32108
rect 4396 32024 4436 32068
rect 4587 32068 4588 32108
rect 4628 32068 4629 32108
rect 4587 32059 4629 32068
rect 4492 32024 4532 32033
rect 4396 31984 4492 32024
rect 4492 31975 4532 31984
rect 4108 31900 4436 31940
rect 4396 31856 4436 31900
rect 4684 31856 4724 32740
rect 5644 32621 5684 32824
rect 5740 32815 5780 32824
rect 5643 32612 5685 32621
rect 5643 32572 5644 32612
rect 5684 32572 5685 32612
rect 5643 32563 5685 32572
rect 6027 32612 6069 32621
rect 6027 32572 6028 32612
rect 6068 32572 6069 32612
rect 6027 32563 6069 32572
rect 4779 32528 4821 32537
rect 4779 32488 4780 32528
rect 4820 32488 4821 32528
rect 4779 32479 4821 32488
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 4780 32360 4820 32479
rect 4972 32360 5012 32369
rect 4780 32320 4972 32360
rect 4972 32311 5012 32320
rect 4780 32192 4820 32201
rect 4780 31949 4820 32152
rect 5068 32192 5108 32201
rect 4779 31940 4821 31949
rect 4779 31900 4780 31940
rect 4820 31900 4821 31940
rect 4779 31891 4821 31900
rect 4396 31816 4724 31856
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 4300 31436 4340 31445
rect 3964 31361 4004 31370
rect 4004 31321 4052 31352
rect 3964 31312 4052 31321
rect 4012 30848 4052 31312
rect 4108 31268 4148 31277
rect 4300 31268 4340 31396
rect 4148 31228 4340 31268
rect 4108 31219 4148 31228
rect 4396 31184 4436 31816
rect 4683 31688 4725 31697
rect 4683 31648 4684 31688
rect 4724 31648 4725 31688
rect 4683 31639 4725 31648
rect 4587 31604 4629 31613
rect 4587 31564 4588 31604
rect 4628 31564 4629 31604
rect 4587 31555 4629 31564
rect 4300 31144 4436 31184
rect 4492 31184 4532 31193
rect 4012 30808 4244 30848
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 3476 30052 3572 30092
rect 3436 30043 3476 30052
rect 4107 30008 4149 30017
rect 4107 29968 4108 30008
rect 4148 29968 4149 30008
rect 4107 29959 4149 29968
rect 3340 29884 3476 29924
rect 3051 29084 3093 29093
rect 3051 29044 3052 29084
rect 3092 29044 3093 29084
rect 3051 29035 3093 29044
rect 2955 28916 2997 28925
rect 2955 28876 2956 28916
rect 2996 28876 2997 28916
rect 2955 28867 2997 28876
rect 2859 27992 2901 28001
rect 2859 27952 2860 27992
rect 2900 27952 2901 27992
rect 2859 27943 2901 27952
rect 2860 26741 2900 27943
rect 2956 27665 2996 28867
rect 3052 28328 3092 29035
rect 3147 28496 3189 28505
rect 3147 28456 3148 28496
rect 3188 28456 3189 28496
rect 3147 28447 3189 28456
rect 3052 27740 3092 28288
rect 3148 28328 3188 28447
rect 3148 28279 3188 28288
rect 3244 28001 3284 29800
rect 3339 29084 3381 29093
rect 3339 29044 3340 29084
rect 3380 29044 3381 29084
rect 3339 29035 3381 29044
rect 3243 27992 3285 28001
rect 3243 27952 3244 27992
rect 3284 27952 3285 27992
rect 3243 27943 3285 27952
rect 3147 27824 3189 27833
rect 3340 27824 3380 29035
rect 3147 27784 3148 27824
rect 3188 27784 3189 27824
rect 3147 27775 3189 27784
rect 3244 27784 3380 27824
rect 3047 27700 3092 27740
rect 2955 27656 2997 27665
rect 2955 27616 2956 27656
rect 2996 27616 2997 27656
rect 2955 27607 2997 27616
rect 3047 27572 3087 27700
rect 3148 27690 3188 27775
rect 3147 27572 3189 27581
rect 3047 27532 3092 27572
rect 2955 27488 2997 27497
rect 2955 27448 2956 27488
rect 2996 27448 2997 27488
rect 2955 27439 2997 27448
rect 2859 26732 2901 26741
rect 2859 26692 2860 26732
rect 2900 26692 2901 26732
rect 2859 26683 2901 26692
rect 2859 26060 2901 26069
rect 2859 26020 2860 26060
rect 2900 26020 2901 26060
rect 2859 26011 2901 26020
rect 2860 25397 2900 26011
rect 2859 25388 2901 25397
rect 2859 25348 2860 25388
rect 2900 25348 2901 25388
rect 2859 25339 2901 25348
rect 2859 25220 2901 25229
rect 2859 25180 2860 25220
rect 2900 25180 2901 25220
rect 2859 25171 2901 25180
rect 2763 23792 2805 23801
rect 2763 23752 2764 23792
rect 2804 23752 2805 23792
rect 2763 23743 2805 23752
rect 2860 23120 2900 25171
rect 2956 23288 2996 27439
rect 3052 26657 3092 27532
rect 3147 27532 3148 27572
rect 3188 27532 3189 27572
rect 3147 27523 3189 27532
rect 3051 26648 3093 26657
rect 3051 26608 3052 26648
rect 3092 26608 3093 26648
rect 3051 26599 3093 26608
rect 3148 26405 3188 27523
rect 3244 26984 3284 27784
rect 3340 27656 3380 27665
rect 3340 27497 3380 27616
rect 3339 27488 3381 27497
rect 3339 27448 3340 27488
rect 3380 27448 3381 27488
rect 3339 27439 3381 27448
rect 3436 27068 3476 29884
rect 3724 29840 3764 29849
rect 3627 29672 3669 29681
rect 3627 29632 3628 29672
rect 3668 29632 3669 29672
rect 3627 29623 3669 29632
rect 3628 29538 3668 29623
rect 3724 29345 3764 29800
rect 3819 29840 3861 29849
rect 3819 29800 3820 29840
rect 3860 29800 3861 29840
rect 3819 29791 3861 29800
rect 3916 29840 3956 29849
rect 3820 29706 3860 29791
rect 3819 29504 3861 29513
rect 3819 29464 3820 29504
rect 3860 29464 3861 29504
rect 3819 29455 3861 29464
rect 3723 29336 3765 29345
rect 3723 29296 3724 29336
rect 3764 29296 3765 29336
rect 3723 29287 3765 29296
rect 3724 29168 3764 29177
rect 3820 29168 3860 29455
rect 3916 29177 3956 29800
rect 4108 29840 4148 29959
rect 4108 29791 4148 29800
rect 4107 29672 4149 29681
rect 4107 29632 4108 29672
rect 4148 29632 4149 29672
rect 4107 29623 4149 29632
rect 4011 29588 4053 29597
rect 4011 29548 4012 29588
rect 4052 29548 4053 29588
rect 4011 29539 4053 29548
rect 3764 29128 3860 29168
rect 3915 29168 3957 29177
rect 3915 29128 3916 29168
rect 3956 29128 3957 29168
rect 3724 28925 3764 29128
rect 3915 29119 3957 29128
rect 3916 29000 3956 29009
rect 4012 29000 4052 29539
rect 3956 28960 4052 29000
rect 3916 28951 3956 28960
rect 3723 28916 3765 28925
rect 3723 28876 3724 28916
rect 3764 28876 3765 28916
rect 3723 28867 3765 28876
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 4108 28505 4148 29623
rect 4107 28496 4149 28505
rect 4107 28456 4108 28496
rect 4148 28456 4149 28496
rect 4107 28447 4149 28456
rect 3531 28412 3573 28421
rect 3531 28372 3532 28412
rect 3572 28372 3573 28412
rect 3531 28363 3573 28372
rect 3532 28278 3572 28363
rect 3627 28328 3669 28337
rect 3627 28288 3628 28328
rect 3668 28288 3669 28328
rect 3627 28279 3669 28288
rect 4107 28328 4149 28337
rect 4107 28288 4108 28328
rect 4148 28288 4149 28328
rect 4107 28279 4149 28288
rect 3628 28194 3668 28279
rect 4108 28194 4148 28279
rect 3627 27740 3669 27749
rect 3627 27700 3628 27740
rect 3668 27700 3764 27740
rect 3627 27691 3669 27700
rect 3531 27656 3573 27665
rect 3531 27616 3532 27656
rect 3572 27616 3573 27656
rect 3531 27607 3573 27616
rect 3724 27656 3764 27700
rect 3724 27607 3764 27616
rect 4107 27656 4149 27665
rect 4107 27616 4108 27656
rect 4148 27616 4149 27656
rect 4107 27607 4149 27616
rect 3532 27522 3572 27607
rect 3531 27404 3573 27413
rect 3531 27364 3532 27404
rect 3572 27364 3573 27404
rect 3531 27355 3573 27364
rect 3532 27270 3572 27355
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 3436 27019 3476 27028
rect 3627 26984 3669 26993
rect 3244 26944 3380 26984
rect 3244 26816 3284 26827
rect 3244 26741 3284 26776
rect 3243 26732 3285 26741
rect 3243 26692 3244 26732
rect 3284 26692 3285 26732
rect 3243 26683 3285 26692
rect 3147 26396 3189 26405
rect 3147 26356 3148 26396
rect 3188 26356 3189 26396
rect 3147 26347 3189 26356
rect 3147 26144 3189 26153
rect 3147 26104 3148 26144
rect 3188 26104 3189 26144
rect 3147 26095 3189 26104
rect 3244 26144 3284 26155
rect 3148 25397 3188 26095
rect 3244 26069 3284 26104
rect 3243 26060 3285 26069
rect 3243 26020 3244 26060
rect 3284 26020 3285 26060
rect 3243 26011 3285 26020
rect 3243 25892 3285 25901
rect 3243 25852 3244 25892
rect 3284 25852 3285 25892
rect 3243 25843 3285 25852
rect 3147 25388 3189 25397
rect 3147 25348 3148 25388
rect 3188 25348 3189 25388
rect 3147 25339 3189 25348
rect 3051 24800 3093 24809
rect 3051 24760 3052 24800
rect 3092 24760 3093 24800
rect 3051 24751 3093 24760
rect 3052 24053 3092 24751
rect 3051 24044 3093 24053
rect 3051 24004 3052 24044
rect 3092 24004 3093 24044
rect 3051 23995 3093 24004
rect 3148 23960 3188 25339
rect 3244 25229 3284 25843
rect 3243 25220 3285 25229
rect 3243 25180 3244 25220
rect 3284 25180 3285 25220
rect 3243 25171 3285 25180
rect 3244 24632 3284 25171
rect 3340 24800 3380 26944
rect 3627 26944 3628 26984
rect 3668 26944 3669 26984
rect 3627 26935 3669 26944
rect 3628 26816 3668 26935
rect 3628 26767 3668 26776
rect 3627 26648 3669 26657
rect 3627 26608 3628 26648
rect 3668 26608 3669 26648
rect 3627 26599 3669 26608
rect 3435 26312 3477 26321
rect 3435 26272 3436 26312
rect 3476 26272 3477 26312
rect 3435 26263 3477 26272
rect 3628 26312 3668 26599
rect 3819 26396 3861 26405
rect 3819 26356 3820 26396
rect 3860 26356 3861 26396
rect 3819 26347 3861 26356
rect 3628 26263 3668 26272
rect 3436 26178 3476 26263
rect 3820 26144 3860 26347
rect 3531 25976 3573 25985
rect 3531 25936 3532 25976
rect 3572 25936 3573 25976
rect 3531 25927 3573 25936
rect 3435 25304 3477 25313
rect 3435 25264 3436 25304
rect 3476 25264 3477 25304
rect 3435 25255 3477 25264
rect 3436 25170 3476 25255
rect 3532 24893 3572 25927
rect 3820 25901 3860 26104
rect 3819 25892 3861 25901
rect 3819 25852 3820 25892
rect 3860 25852 3861 25892
rect 3819 25843 3861 25852
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 4011 25556 4053 25565
rect 4011 25516 4012 25556
rect 4052 25516 4053 25556
rect 4011 25507 4053 25516
rect 4012 25318 4052 25507
rect 4012 25269 4052 25278
rect 3820 25220 3860 25229
rect 4108 25220 4148 27607
rect 4204 26321 4244 30808
rect 4300 28673 4340 31144
rect 4492 30941 4532 31144
rect 4491 30932 4533 30941
rect 4491 30892 4492 30932
rect 4532 30892 4533 30932
rect 4491 30883 4533 30892
rect 4395 30680 4437 30689
rect 4395 30640 4396 30680
rect 4436 30640 4437 30680
rect 4395 30631 4437 30640
rect 4588 30680 4628 31555
rect 4396 29597 4436 30631
rect 4588 29849 4628 30640
rect 4587 29840 4629 29849
rect 4587 29800 4588 29840
rect 4628 29800 4629 29840
rect 4587 29791 4629 29800
rect 4395 29588 4437 29597
rect 4395 29548 4396 29588
rect 4436 29548 4437 29588
rect 4395 29539 4437 29548
rect 4588 29513 4628 29791
rect 4684 29681 4724 31639
rect 5068 31520 5108 32152
rect 5452 31529 5492 31614
rect 5451 31520 5493 31529
rect 5068 31480 5396 31520
rect 4780 31352 4820 31361
rect 4780 30689 4820 31312
rect 5067 31352 5109 31361
rect 5067 31312 5068 31352
rect 5108 31312 5109 31352
rect 5067 31303 5109 31312
rect 5068 31218 5108 31303
rect 5163 31268 5205 31277
rect 5163 31228 5164 31268
rect 5204 31228 5205 31268
rect 5163 31219 5205 31228
rect 5164 31134 5204 31219
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 4779 30680 4821 30689
rect 4779 30640 4780 30680
rect 4820 30640 4821 30680
rect 4779 30631 4821 30640
rect 5067 30680 5109 30689
rect 5067 30640 5068 30680
rect 5108 30640 5109 30680
rect 5067 30631 5109 30640
rect 5164 30680 5204 30689
rect 5068 30546 5108 30631
rect 5164 30437 5204 30640
rect 5356 30521 5396 31480
rect 5451 31480 5452 31520
rect 5492 31480 5493 31520
rect 5451 31471 5493 31480
rect 5931 31520 5973 31529
rect 5931 31480 5932 31520
rect 5972 31480 5973 31520
rect 5931 31471 5973 31480
rect 5644 31352 5684 31361
rect 5644 31193 5684 31312
rect 5643 31184 5685 31193
rect 5643 31144 5644 31184
rect 5684 31144 5685 31184
rect 5643 31135 5685 31144
rect 5451 31016 5493 31025
rect 5451 30976 5452 31016
rect 5492 30976 5493 31016
rect 5451 30967 5493 30976
rect 5355 30512 5397 30521
rect 5355 30472 5356 30512
rect 5396 30472 5397 30512
rect 5355 30463 5397 30472
rect 4780 30428 4820 30437
rect 4780 30269 4820 30388
rect 5163 30428 5205 30437
rect 5163 30388 5164 30428
rect 5204 30388 5205 30428
rect 5163 30379 5205 30388
rect 4779 30260 4821 30269
rect 4779 30220 4780 30260
rect 4820 30220 4821 30260
rect 4779 30211 4821 30220
rect 5452 29933 5492 30967
rect 5547 30596 5589 30605
rect 5547 30556 5548 30596
rect 5588 30556 5589 30596
rect 5547 30547 5589 30556
rect 5644 30596 5684 30607
rect 5548 30462 5588 30547
rect 5644 30521 5684 30556
rect 5643 30512 5685 30521
rect 5643 30472 5644 30512
rect 5684 30472 5685 30512
rect 5643 30463 5685 30472
rect 5739 30428 5781 30437
rect 5739 30388 5740 30428
rect 5780 30388 5781 30428
rect 5739 30379 5781 30388
rect 5451 29924 5493 29933
rect 5451 29884 5452 29924
rect 5492 29884 5493 29924
rect 5451 29875 5493 29884
rect 5355 29840 5397 29849
rect 5355 29800 5356 29840
rect 5396 29800 5397 29840
rect 5355 29791 5397 29800
rect 5356 29706 5396 29791
rect 4683 29672 4725 29681
rect 4683 29632 4684 29672
rect 4724 29632 4725 29672
rect 4683 29623 4725 29632
rect 4587 29504 4629 29513
rect 4587 29464 4588 29504
rect 4628 29464 4629 29504
rect 4587 29455 4629 29464
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 5355 29504 5397 29513
rect 5355 29464 5356 29504
rect 5396 29464 5397 29504
rect 5355 29455 5397 29464
rect 4780 29336 4820 29345
rect 4396 29296 4780 29336
rect 4299 28664 4341 28673
rect 4299 28624 4300 28664
rect 4340 28624 4341 28664
rect 4299 28615 4341 28624
rect 4299 28496 4341 28505
rect 4299 28456 4300 28496
rect 4340 28456 4341 28496
rect 4299 28447 4341 28456
rect 4203 26312 4245 26321
rect 4203 26272 4204 26312
rect 4244 26272 4245 26312
rect 4203 26263 4245 26272
rect 3860 25180 4148 25220
rect 3820 25171 3860 25180
rect 4107 24968 4149 24977
rect 4107 24928 4108 24968
rect 4148 24928 4149 24968
rect 4107 24919 4149 24928
rect 3531 24884 3573 24893
rect 3531 24844 3532 24884
rect 3572 24844 3573 24884
rect 3531 24835 3573 24844
rect 3436 24800 3476 24809
rect 3340 24760 3436 24800
rect 3436 24751 3476 24760
rect 3724 24716 3764 24725
rect 3244 24583 3284 24592
rect 3532 24676 3724 24716
rect 3436 23960 3476 23969
rect 3148 23920 3436 23960
rect 3436 23911 3476 23920
rect 3532 23801 3572 24676
rect 3724 24667 3764 24676
rect 3915 24632 3957 24641
rect 3915 24587 3916 24632
rect 3956 24587 3957 24632
rect 3915 24583 3957 24587
rect 3916 24497 3956 24583
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 3627 24044 3669 24053
rect 3627 24004 3628 24044
rect 3668 24004 3669 24044
rect 3627 23995 3669 24004
rect 3628 23910 3668 23995
rect 3147 23792 3189 23801
rect 3147 23752 3148 23792
rect 3188 23752 3189 23792
rect 3147 23743 3189 23752
rect 3244 23792 3284 23801
rect 3531 23792 3573 23801
rect 3284 23752 3380 23792
rect 3244 23743 3284 23752
rect 3148 23624 3188 23743
rect 3148 23584 3284 23624
rect 2956 23248 3092 23288
rect 2956 23120 2996 23129
rect 2860 23080 2956 23120
rect 2667 22616 2709 22625
rect 2667 22576 2668 22616
rect 2708 22576 2709 22616
rect 2667 22567 2709 22576
rect 2668 22532 2708 22567
rect 2668 22481 2708 22492
rect 2860 22457 2900 23080
rect 2956 23071 2996 23080
rect 3052 22541 3092 23248
rect 3148 23204 3188 23215
rect 3148 23129 3188 23164
rect 3147 23120 3189 23129
rect 3147 23080 3148 23120
rect 3188 23080 3189 23120
rect 3147 23071 3189 23080
rect 3051 22532 3093 22541
rect 3051 22492 3052 22532
rect 3092 22492 3093 22532
rect 3051 22483 3093 22492
rect 2859 22448 2901 22457
rect 2859 22408 2860 22448
rect 2900 22408 2901 22448
rect 2859 22399 2901 22408
rect 2667 22364 2709 22373
rect 2667 22324 2668 22364
rect 2708 22324 2709 22364
rect 2667 22315 2709 22324
rect 2668 22112 2708 22315
rect 3052 22299 3092 22308
rect 2860 22259 3052 22285
rect 2860 22245 3092 22259
rect 3148 22280 3188 22289
rect 2668 22072 2804 22112
rect 2764 21608 2804 22072
rect 2764 21559 2804 21568
rect 2860 21533 2900 22245
rect 3148 22196 3188 22240
rect 3052 22156 3188 22196
rect 2955 21776 2997 21785
rect 2955 21736 2956 21776
rect 2996 21736 2997 21776
rect 2955 21727 2997 21736
rect 2956 21642 2996 21727
rect 2667 21524 2709 21533
rect 2667 21484 2668 21524
rect 2708 21484 2709 21524
rect 2667 21475 2709 21484
rect 2859 21524 2901 21533
rect 2859 21484 2860 21524
rect 2900 21484 2901 21524
rect 2859 21475 2901 21484
rect 2668 21020 2708 21475
rect 2668 20971 2708 20980
rect 2860 20852 2900 21475
rect 2668 20812 2900 20852
rect 2571 20516 2613 20525
rect 2571 20476 2572 20516
rect 2612 20476 2613 20516
rect 2571 20467 2613 20476
rect 2668 20348 2708 20812
rect 2956 20768 2996 20777
rect 2476 19256 2516 20056
rect 2572 20308 2708 20348
rect 2764 20728 2956 20768
rect 2572 19508 2612 20308
rect 2667 20180 2709 20189
rect 2667 20140 2668 20180
rect 2708 20140 2709 20180
rect 2667 20131 2709 20140
rect 2668 20046 2708 20131
rect 2668 19508 2708 19517
rect 2572 19468 2668 19508
rect 2668 19459 2708 19468
rect 2571 19340 2613 19349
rect 2571 19300 2572 19340
rect 2612 19300 2613 19340
rect 2571 19291 2613 19300
rect 2476 19207 2516 19216
rect 2475 18668 2517 18677
rect 2475 18628 2476 18668
rect 2516 18628 2517 18668
rect 2475 18619 2517 18628
rect 2476 18584 2516 18619
rect 2476 18533 2516 18544
rect 2475 17996 2517 18005
rect 2475 17956 2476 17996
rect 2516 17956 2517 17996
rect 2475 17947 2517 17956
rect 2380 17744 2420 17753
rect 2380 17408 2420 17704
rect 2476 17744 2516 17947
rect 2476 17669 2516 17704
rect 2475 17660 2517 17669
rect 2475 17620 2476 17660
rect 2516 17620 2517 17660
rect 2475 17611 2517 17620
rect 2572 17492 2612 19291
rect 2668 18752 2708 18761
rect 2764 18752 2804 20728
rect 2956 20719 2996 20728
rect 3052 20768 3092 22156
rect 3147 22028 3189 22037
rect 3147 21988 3148 22028
rect 3188 21988 3189 22028
rect 3147 21979 3189 21988
rect 2859 20600 2901 20609
rect 2859 20560 2860 20600
rect 2900 20560 2901 20600
rect 2859 20551 2901 20560
rect 2860 20096 2900 20551
rect 3052 20189 3092 20728
rect 3051 20180 3093 20189
rect 3051 20140 3052 20180
rect 3092 20140 3093 20180
rect 3051 20131 3093 20140
rect 2860 20047 2900 20056
rect 2708 18712 2804 18752
rect 3052 19256 3092 19265
rect 2668 18703 2708 18712
rect 3052 18416 3092 19216
rect 3052 18173 3092 18376
rect 3051 18164 3093 18173
rect 3051 18124 3052 18164
rect 3092 18124 3093 18164
rect 3051 18115 3093 18124
rect 3148 17996 3188 21979
rect 3052 17956 3188 17996
rect 3244 17996 3284 23584
rect 3340 23549 3380 23752
rect 3531 23752 3532 23792
rect 3572 23752 3573 23792
rect 3531 23743 3573 23752
rect 4011 23792 4053 23801
rect 4011 23752 4012 23792
rect 4052 23752 4053 23792
rect 4011 23743 4053 23752
rect 3915 23708 3957 23717
rect 3915 23668 3916 23708
rect 3956 23668 3957 23708
rect 3915 23659 3957 23668
rect 3916 23574 3956 23659
rect 4012 23658 4052 23743
rect 3339 23540 3381 23549
rect 3339 23500 3340 23540
rect 3380 23500 3381 23540
rect 3339 23491 3381 23500
rect 3435 23288 3477 23297
rect 3435 23248 3436 23288
rect 3476 23248 3477 23288
rect 3435 23239 3477 23248
rect 4012 23288 4052 23297
rect 4108 23288 4148 24919
rect 4300 24212 4340 28447
rect 4396 27077 4436 29296
rect 4780 29287 4820 29296
rect 4971 29336 5013 29345
rect 5163 29336 5205 29345
rect 4971 29296 4972 29336
rect 5012 29296 5013 29336
rect 4971 29287 5013 29296
rect 5068 29296 5164 29336
rect 5204 29296 5205 29336
rect 4972 29202 5012 29287
rect 4492 29168 4532 29177
rect 4492 29093 4532 29128
rect 4588 29168 4628 29177
rect 4628 29128 4724 29168
rect 4588 29119 4628 29128
rect 4484 29084 4532 29093
rect 4484 29044 4485 29084
rect 4525 29044 4532 29084
rect 4484 29035 4526 29044
rect 4587 29000 4629 29009
rect 4587 28960 4588 29000
rect 4628 28960 4629 29000
rect 4684 29000 4724 29128
rect 5068 29093 5108 29296
rect 5163 29287 5205 29296
rect 5163 29168 5205 29177
rect 5163 29128 5164 29168
rect 5204 29128 5205 29168
rect 5163 29119 5205 29128
rect 5260 29168 5300 29177
rect 5356 29168 5396 29455
rect 5300 29128 5396 29168
rect 5452 29168 5492 29875
rect 5547 29840 5589 29849
rect 5547 29800 5548 29840
rect 5588 29800 5589 29840
rect 5547 29791 5589 29800
rect 5548 29756 5588 29791
rect 5548 29705 5588 29716
rect 5260 29119 5300 29128
rect 5067 29084 5109 29093
rect 5067 29044 5068 29084
rect 5108 29044 5109 29084
rect 5067 29035 5109 29044
rect 4684 28960 4820 29000
rect 4587 28951 4629 28960
rect 4491 28664 4533 28673
rect 4491 28624 4492 28664
rect 4532 28624 4533 28664
rect 4491 28615 4533 28624
rect 4395 27068 4437 27077
rect 4395 27028 4396 27068
rect 4436 27028 4437 27068
rect 4395 27019 4437 27028
rect 4492 26816 4532 28615
rect 4588 28333 4628 28951
rect 4588 27833 4628 28293
rect 4780 28244 4820 28960
rect 5068 28328 5108 29035
rect 5164 29034 5204 29119
rect 5068 28279 5108 28288
rect 4780 28195 4820 28204
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 4587 27824 4629 27833
rect 4587 27784 4588 27824
rect 4628 27784 4629 27824
rect 5452 27824 5492 29128
rect 5643 29084 5685 29093
rect 5643 29044 5644 29084
rect 5684 29044 5685 29084
rect 5643 29035 5685 29044
rect 5644 27992 5684 29035
rect 5740 28253 5780 30379
rect 5835 29840 5877 29849
rect 5835 29800 5836 29840
rect 5876 29800 5877 29840
rect 5835 29791 5877 29800
rect 5932 29840 5972 31471
rect 6028 30428 6068 32563
rect 6124 32201 6164 33739
rect 6316 33620 6356 34756
rect 6411 34544 6453 34553
rect 6411 34504 6412 34544
rect 6452 34504 6453 34544
rect 6411 34495 6453 34504
rect 6412 34217 6452 34495
rect 6411 34208 6453 34217
rect 6411 34168 6412 34208
rect 6452 34168 6453 34208
rect 6411 34159 6453 34168
rect 6123 32192 6165 32201
rect 6123 32152 6124 32192
rect 6164 32152 6165 32192
rect 6123 32143 6165 32152
rect 6124 30680 6164 30689
rect 6316 30680 6356 33580
rect 6412 33620 6452 33631
rect 6412 33545 6452 33580
rect 6411 33536 6453 33545
rect 6411 33496 6412 33536
rect 6452 33496 6453 33536
rect 6411 33487 6453 33496
rect 6508 33368 6548 35008
rect 6604 34385 6644 35848
rect 6700 35720 6740 35729
rect 6700 35225 6740 35680
rect 6892 35552 6932 35848
rect 6988 35888 7028 35897
rect 7180 35888 7220 35897
rect 7276 35888 7316 37939
rect 7372 37400 7412 37409
rect 7372 37157 7412 37360
rect 7371 37148 7413 37157
rect 7371 37108 7372 37148
rect 7412 37108 7413 37148
rect 7371 37099 7413 37108
rect 7372 36728 7412 36737
rect 7372 36233 7412 36688
rect 7371 36224 7413 36233
rect 7371 36184 7372 36224
rect 7412 36184 7413 36224
rect 7371 36175 7413 36184
rect 7371 36056 7413 36065
rect 7371 36016 7372 36056
rect 7412 36016 7413 36056
rect 7371 36007 7413 36016
rect 7028 35848 7124 35888
rect 6988 35839 7028 35848
rect 7084 35720 7124 35848
rect 7220 35848 7316 35888
rect 7372 35888 7412 36007
rect 7180 35839 7220 35848
rect 7084 35680 7220 35720
rect 6796 35512 6932 35552
rect 6699 35216 6741 35225
rect 6699 35176 6700 35216
rect 6740 35176 6741 35216
rect 6699 35167 6741 35176
rect 6700 34553 6740 35167
rect 6796 34637 6836 35512
rect 6987 35384 7029 35393
rect 6987 35344 6988 35384
rect 7028 35344 7029 35384
rect 6987 35335 7029 35344
rect 6892 35216 6932 35225
rect 6892 34805 6932 35176
rect 6891 34796 6933 34805
rect 6891 34756 6892 34796
rect 6932 34756 6933 34796
rect 6891 34747 6933 34756
rect 6795 34628 6837 34637
rect 6795 34588 6796 34628
rect 6836 34588 6837 34628
rect 6795 34579 6837 34588
rect 6699 34544 6741 34553
rect 6699 34504 6700 34544
rect 6740 34504 6741 34544
rect 6699 34495 6741 34504
rect 6603 34376 6645 34385
rect 6603 34336 6604 34376
rect 6644 34336 6645 34376
rect 6603 34327 6645 34336
rect 6699 34292 6741 34301
rect 6699 34252 6700 34292
rect 6740 34252 6741 34292
rect 6699 34243 6741 34252
rect 6164 30640 6356 30680
rect 6124 30631 6164 30640
rect 6028 30388 6164 30428
rect 6027 30260 6069 30269
rect 6027 30220 6028 30260
rect 6068 30220 6069 30260
rect 6027 30211 6069 30220
rect 5932 29791 5972 29800
rect 6028 29840 6068 30211
rect 6028 29791 6068 29800
rect 5836 29706 5876 29791
rect 6124 29672 6164 30388
rect 6219 30176 6261 30185
rect 6219 30136 6220 30176
rect 6260 30136 6261 30176
rect 6219 30127 6261 30136
rect 6220 30092 6260 30127
rect 6220 30041 6260 30052
rect 6316 29840 6356 30640
rect 6412 33328 6548 33368
rect 6412 30437 6452 33328
rect 6700 31529 6740 34243
rect 6892 34217 6932 34747
rect 6891 34208 6933 34217
rect 6891 34168 6892 34208
rect 6932 34168 6933 34208
rect 6891 34159 6933 34168
rect 6891 33704 6933 33713
rect 6891 33664 6892 33704
rect 6932 33664 6933 33704
rect 6891 33655 6933 33664
rect 6892 33570 6932 33655
rect 6988 33032 7028 35335
rect 7180 35300 7220 35680
rect 7372 35645 7412 35848
rect 7371 35636 7413 35645
rect 7371 35596 7372 35636
rect 7412 35596 7413 35636
rect 7371 35587 7413 35596
rect 6892 32992 7028 33032
rect 7084 35260 7220 35300
rect 6795 32948 6837 32957
rect 6795 32908 6796 32948
rect 6836 32908 6837 32948
rect 6795 32899 6837 32908
rect 6699 31520 6741 31529
rect 6699 31480 6700 31520
rect 6740 31480 6741 31520
rect 6699 31471 6741 31480
rect 6796 30932 6836 32899
rect 6892 31361 6932 32992
rect 6988 32864 7028 32873
rect 6988 32117 7028 32824
rect 7084 32369 7124 35260
rect 7371 35216 7413 35225
rect 7371 35171 7372 35216
rect 7412 35171 7413 35216
rect 7371 35167 7413 35171
rect 7372 35081 7412 35167
rect 7371 34544 7413 34553
rect 7371 34504 7372 34544
rect 7412 34504 7413 34544
rect 7371 34495 7413 34504
rect 7372 34376 7412 34495
rect 7180 34336 7372 34376
rect 7180 33377 7220 34336
rect 7372 34327 7412 34336
rect 7468 34040 7508 38947
rect 7563 38240 7605 38249
rect 7563 38200 7564 38240
rect 7604 38200 7605 38240
rect 7563 38191 7605 38200
rect 7564 35300 7604 38191
rect 7660 37745 7700 40459
rect 8044 40433 8084 40879
rect 8235 40676 8277 40685
rect 8620 40676 8660 41215
rect 8811 40760 8853 40769
rect 8811 40720 8812 40760
rect 8852 40720 8853 40760
rect 8811 40711 8853 40720
rect 8235 40636 8236 40676
rect 8276 40636 8277 40676
rect 8235 40627 8277 40636
rect 8428 40636 8660 40676
rect 8236 40542 8276 40627
rect 8043 40424 8085 40433
rect 8043 40384 8044 40424
rect 8084 40384 8085 40424
rect 8043 40375 8085 40384
rect 8044 40290 8084 40375
rect 8428 40265 8468 40636
rect 8619 40424 8661 40433
rect 8619 40384 8620 40424
rect 8660 40384 8661 40424
rect 8619 40375 8661 40384
rect 8427 40256 8469 40265
rect 8427 40216 8428 40256
rect 8468 40216 8469 40256
rect 8427 40207 8469 40216
rect 8428 40122 8468 40207
rect 8139 39836 8181 39845
rect 8139 39796 8140 39836
rect 8180 39796 8181 39836
rect 8139 39787 8181 39796
rect 7948 39738 7988 39747
rect 8140 39702 8180 39787
rect 7948 39089 7988 39698
rect 7947 39080 7989 39089
rect 7947 39040 7948 39080
rect 7988 39040 7989 39080
rect 7947 39031 7989 39040
rect 8620 39005 8660 40375
rect 8812 39593 8852 40711
rect 8811 39584 8853 39593
rect 8811 39544 8812 39584
rect 8852 39544 8853 39584
rect 8811 39535 8853 39544
rect 8811 39080 8853 39089
rect 8811 39040 8812 39080
rect 8852 39040 8853 39080
rect 8811 39031 8853 39040
rect 8619 38996 8661 39005
rect 8619 38956 8620 38996
rect 8660 38956 8661 38996
rect 8619 38947 8661 38956
rect 8620 38912 8660 38947
rect 8812 38946 8852 39031
rect 7948 38324 7988 38333
rect 7756 38226 7796 38235
rect 7659 37736 7701 37745
rect 7659 37696 7660 37736
rect 7700 37696 7701 37736
rect 7659 37687 7701 37696
rect 7564 35251 7604 35260
rect 7660 34301 7700 37687
rect 7756 37661 7796 38186
rect 7755 37652 7797 37661
rect 7755 37612 7756 37652
rect 7796 37612 7797 37652
rect 7755 37603 7797 37612
rect 7948 37493 7988 38284
rect 8140 38249 8180 38334
rect 8139 38240 8181 38249
rect 8139 38200 8140 38240
rect 8180 38200 8181 38240
rect 8139 38191 8181 38200
rect 8332 38240 8372 38249
rect 8139 37988 8181 37997
rect 8139 37948 8140 37988
rect 8180 37948 8181 37988
rect 8139 37939 8181 37948
rect 8140 37854 8180 37939
rect 7947 37484 7989 37493
rect 7947 37444 7948 37484
rect 7988 37444 7989 37484
rect 7947 37435 7989 37444
rect 8332 36569 8372 38200
rect 8620 37400 8660 38872
rect 8908 38249 8948 53563
rect 9003 53528 9045 53537
rect 9003 53488 9004 53528
rect 9044 53488 9045 53528
rect 9003 53479 9045 53488
rect 9004 53360 9044 53479
rect 9004 53311 9044 53320
rect 9003 53108 9045 53117
rect 9003 53068 9004 53108
rect 9044 53068 9045 53108
rect 9003 53059 9045 53068
rect 9004 43793 9044 53059
rect 9100 52445 9140 53824
rect 9099 52436 9141 52445
rect 9099 52396 9100 52436
rect 9140 52396 9141 52436
rect 9099 52387 9141 52396
rect 9196 51689 9236 59872
rect 9388 59753 9428 66079
rect 9483 65624 9525 65633
rect 9483 65584 9484 65624
rect 9524 65584 9525 65624
rect 9483 65575 9525 65584
rect 9484 61769 9524 65575
rect 9580 64280 9620 69532
rect 9676 68489 9716 69952
rect 9772 69077 9812 79183
rect 9867 77552 9909 77561
rect 9867 77512 9868 77552
rect 9908 77512 9909 77552
rect 9867 77503 9909 77512
rect 9868 71504 9908 77503
rect 9964 76889 10004 81880
rect 10059 77552 10101 77561
rect 10059 77512 10060 77552
rect 10100 77512 10101 77552
rect 10059 77503 10101 77512
rect 10060 77418 10100 77503
rect 10156 77132 10196 82291
rect 10252 77645 10292 85936
rect 10347 83684 10389 83693
rect 10347 83644 10348 83684
rect 10388 83644 10389 83684
rect 10347 83635 10389 83644
rect 10348 83012 10388 83635
rect 10444 83189 10484 85936
rect 10636 84449 10676 85936
rect 10635 84440 10677 84449
rect 10635 84400 10636 84440
rect 10676 84400 10677 84440
rect 10635 84391 10677 84400
rect 10443 83180 10485 83189
rect 10443 83140 10444 83180
rect 10484 83140 10485 83180
rect 10443 83131 10485 83140
rect 10348 82972 10484 83012
rect 10444 81920 10484 82972
rect 10444 81880 10676 81920
rect 10539 79148 10581 79157
rect 10539 79108 10540 79148
rect 10580 79108 10581 79148
rect 10539 79099 10581 79108
rect 10348 79064 10388 79073
rect 10348 78065 10388 79024
rect 10540 79014 10580 79099
rect 10636 78140 10676 81880
rect 10732 79568 10772 79577
rect 10732 79409 10772 79528
rect 10731 79400 10773 79409
rect 10731 79360 10732 79400
rect 10772 79360 10773 79400
rect 10731 79351 10773 79360
rect 10732 78149 10772 79351
rect 10828 79325 10868 85936
rect 10923 83432 10965 83441
rect 10923 83392 10924 83432
rect 10964 83392 10965 83432
rect 10923 83383 10965 83392
rect 10827 79316 10869 79325
rect 10827 79276 10828 79316
rect 10868 79276 10869 79316
rect 10827 79267 10869 79276
rect 10827 79148 10869 79157
rect 10827 79108 10828 79148
rect 10868 79108 10869 79148
rect 10827 79099 10869 79108
rect 10828 79064 10868 79099
rect 10924 79073 10964 83383
rect 11020 82349 11060 85936
rect 11019 82340 11061 82349
rect 11019 82300 11020 82340
rect 11060 82300 11061 82340
rect 11019 82291 11061 82300
rect 11212 82088 11252 85936
rect 11404 83861 11444 85936
rect 11403 83852 11445 83861
rect 11403 83812 11404 83852
rect 11444 83812 11445 83852
rect 11403 83803 11445 83812
rect 11116 82048 11252 82088
rect 11019 79736 11061 79745
rect 11019 79696 11020 79736
rect 11060 79696 11061 79736
rect 11019 79687 11061 79696
rect 11020 79602 11060 79687
rect 11019 79148 11061 79157
rect 11019 79108 11020 79148
rect 11060 79108 11061 79148
rect 11019 79099 11061 79108
rect 10828 79013 10868 79024
rect 10923 79064 10965 79073
rect 10923 79024 10924 79064
rect 10964 79024 10965 79064
rect 10923 79015 10965 79024
rect 10924 78930 10964 79015
rect 10540 78100 10676 78140
rect 10731 78140 10773 78149
rect 10731 78100 10732 78140
rect 10772 78100 10773 78140
rect 10347 78056 10389 78065
rect 10347 78016 10348 78056
rect 10388 78016 10389 78056
rect 10347 78007 10389 78016
rect 10251 77636 10293 77645
rect 10251 77596 10252 77636
rect 10292 77596 10293 77636
rect 10251 77587 10293 77596
rect 10348 77561 10388 78007
rect 10347 77552 10389 77561
rect 10347 77512 10348 77552
rect 10388 77512 10389 77552
rect 10347 77503 10389 77512
rect 10540 77384 10580 78100
rect 10731 78091 10773 78100
rect 10732 78006 10772 78091
rect 10923 77636 10965 77645
rect 10923 77596 10924 77636
rect 10964 77596 10965 77636
rect 10923 77587 10965 77596
rect 10636 77552 10676 77561
rect 10676 77512 10868 77552
rect 10636 77503 10676 77512
rect 10540 77344 10676 77384
rect 10252 77300 10292 77309
rect 10292 77260 10484 77300
rect 10252 77251 10292 77260
rect 10156 77092 10292 77132
rect 9963 76880 10005 76889
rect 9963 76840 9964 76880
rect 10004 76840 10005 76880
rect 9963 76831 10005 76840
rect 9964 76717 10004 76726
rect 9964 76292 10004 76677
rect 10155 76544 10197 76553
rect 10155 76504 10156 76544
rect 10196 76504 10197 76544
rect 10155 76495 10197 76504
rect 10156 76410 10196 76495
rect 9964 76252 10196 76292
rect 10156 76208 10196 76252
rect 10156 76159 10196 76168
rect 9963 76040 10005 76049
rect 9963 76000 9964 76040
rect 10004 76000 10005 76040
rect 9963 75991 10005 76000
rect 10155 76040 10197 76049
rect 10155 76000 10156 76040
rect 10196 76000 10197 76040
rect 10155 75991 10197 76000
rect 9964 75906 10004 75991
rect 10156 75209 10196 75991
rect 10252 75629 10292 77092
rect 10347 76964 10389 76973
rect 10347 76924 10348 76964
rect 10388 76924 10389 76964
rect 10347 76915 10389 76924
rect 10348 76544 10388 76915
rect 10444 76712 10484 77260
rect 10444 76663 10484 76672
rect 10540 76712 10580 76721
rect 10636 76712 10676 77344
rect 10580 76672 10676 76712
rect 10540 76663 10580 76672
rect 10348 76504 10580 76544
rect 10443 76292 10485 76301
rect 10443 76252 10444 76292
rect 10484 76252 10485 76292
rect 10443 76243 10485 76252
rect 10347 75872 10389 75881
rect 10347 75832 10348 75872
rect 10388 75832 10389 75872
rect 10347 75823 10389 75832
rect 10348 75738 10388 75823
rect 10251 75620 10293 75629
rect 10444 75620 10484 76243
rect 10251 75580 10252 75620
rect 10292 75580 10293 75620
rect 10251 75571 10293 75580
rect 10348 75580 10484 75620
rect 10155 75200 10197 75209
rect 10155 75160 10156 75200
rect 10196 75160 10197 75200
rect 10155 75151 10197 75160
rect 10059 75032 10101 75041
rect 10059 74992 10060 75032
rect 10100 74992 10101 75032
rect 10059 74983 10101 74992
rect 10060 74523 10100 74983
rect 10251 74780 10293 74789
rect 10251 74740 10252 74780
rect 10292 74740 10293 74780
rect 10251 74731 10293 74740
rect 10252 74696 10292 74731
rect 10252 74645 10292 74656
rect 10060 74474 10100 74483
rect 10060 73693 10100 73702
rect 10060 73109 10100 73653
rect 10252 73520 10292 73529
rect 10059 73100 10101 73109
rect 10059 73060 10060 73100
rect 10100 73060 10101 73100
rect 10059 73051 10101 73060
rect 9964 73016 10004 73025
rect 9964 72437 10004 72976
rect 10155 72848 10197 72857
rect 10155 72808 10156 72848
rect 10196 72808 10197 72848
rect 10155 72799 10197 72808
rect 10156 72714 10196 72799
rect 9963 72428 10005 72437
rect 9963 72388 9964 72428
rect 10004 72388 10005 72428
rect 9963 72379 10005 72388
rect 10060 71504 10100 71513
rect 9868 71464 10060 71504
rect 10060 71455 10100 71464
rect 10252 70160 10292 73480
rect 10348 73193 10388 75580
rect 10443 75200 10485 75209
rect 10443 75160 10444 75200
rect 10484 75160 10485 75200
rect 10443 75151 10485 75160
rect 10444 75066 10484 75151
rect 10347 73184 10389 73193
rect 10347 73144 10348 73184
rect 10388 73144 10389 73184
rect 10347 73135 10389 73144
rect 10540 73100 10580 76504
rect 10636 75713 10676 76672
rect 10731 76544 10773 76553
rect 10731 76504 10732 76544
rect 10772 76504 10773 76544
rect 10731 76495 10773 76504
rect 10635 75704 10677 75713
rect 10635 75664 10636 75704
rect 10676 75664 10677 75704
rect 10635 75655 10677 75664
rect 10635 75032 10677 75041
rect 10635 74992 10636 75032
rect 10676 74992 10677 75032
rect 10635 74983 10677 74992
rect 10636 74898 10676 74983
rect 10635 74696 10677 74705
rect 10635 74656 10636 74696
rect 10676 74656 10677 74696
rect 10635 74647 10677 74656
rect 10444 73060 10580 73100
rect 10347 73016 10389 73025
rect 10347 72976 10348 73016
rect 10388 72976 10389 73016
rect 10347 72967 10389 72976
rect 10348 72882 10388 72967
rect 10347 72680 10389 72689
rect 10347 72640 10348 72680
rect 10388 72640 10389 72680
rect 10347 72631 10389 72640
rect 10348 72176 10388 72631
rect 10348 72127 10388 72136
rect 10347 71840 10389 71849
rect 10444 71840 10484 73060
rect 10636 72689 10676 74647
rect 10732 73100 10772 76495
rect 10828 75536 10868 77512
rect 10924 76796 10964 77587
rect 11020 76973 11060 79099
rect 11019 76964 11061 76973
rect 11019 76924 11020 76964
rect 11060 76924 11061 76964
rect 11019 76915 11061 76924
rect 10924 76553 10964 76756
rect 11020 76712 11060 76721
rect 10923 76544 10965 76553
rect 10923 76504 10924 76544
rect 10964 76504 10965 76544
rect 10923 76495 10965 76504
rect 11020 75881 11060 76672
rect 11019 75872 11061 75881
rect 11019 75832 11020 75872
rect 11060 75832 11061 75872
rect 11019 75823 11061 75832
rect 10828 75496 11060 75536
rect 10923 75368 10965 75377
rect 10923 75328 10924 75368
rect 10964 75328 10965 75368
rect 10923 75319 10965 75328
rect 10828 75200 10868 75209
rect 10828 74453 10868 75160
rect 10924 74528 10964 75319
rect 10924 74479 10964 74488
rect 10827 74444 10869 74453
rect 10827 74404 10828 74444
rect 10868 74404 10869 74444
rect 10827 74395 10869 74404
rect 10732 73060 10868 73100
rect 10635 72680 10677 72689
rect 10635 72640 10636 72680
rect 10676 72640 10677 72680
rect 10635 72631 10677 72640
rect 10347 71800 10348 71840
rect 10388 71800 10484 71840
rect 10347 71791 10389 71800
rect 10348 70664 10388 71791
rect 10731 71588 10773 71597
rect 10731 71548 10732 71588
rect 10772 71548 10773 71588
rect 10731 71539 10773 71548
rect 10540 71490 10580 71499
rect 10732 71454 10772 71539
rect 10540 70925 10580 71450
rect 10539 70916 10581 70925
rect 10539 70876 10540 70916
rect 10580 70876 10581 70916
rect 10539 70867 10581 70876
rect 10348 70615 10388 70624
rect 10539 70160 10581 70169
rect 10252 70120 10484 70160
rect 9868 70076 9908 70085
rect 9908 70036 10196 70076
rect 9868 70027 9908 70036
rect 10156 69992 10196 70036
rect 10156 69943 10196 69952
rect 10252 69992 10292 70001
rect 9868 69364 10196 69404
rect 9771 69068 9813 69077
rect 9771 69028 9772 69068
rect 9812 69028 9813 69068
rect 9771 69019 9813 69028
rect 9868 68900 9908 69364
rect 10059 69236 10101 69245
rect 10059 69196 10060 69236
rect 10100 69196 10101 69236
rect 10059 69187 10101 69196
rect 10060 68984 10100 69187
rect 10156 69152 10196 69364
rect 10156 69103 10196 69112
rect 10155 68984 10197 68993
rect 10060 68944 10156 68984
rect 10196 68944 10197 68984
rect 10155 68935 10197 68944
rect 9772 68860 9908 68900
rect 9675 68480 9717 68489
rect 9675 68440 9676 68480
rect 9716 68440 9717 68480
rect 9675 68431 9717 68440
rect 9676 68228 9716 68237
rect 9676 67640 9716 68188
rect 9772 67901 9812 68860
rect 9963 68480 10005 68489
rect 9963 68440 9964 68480
rect 10004 68440 10005 68480
rect 9963 68431 10005 68440
rect 9867 68396 9909 68405
rect 9867 68356 9868 68396
rect 9908 68356 9909 68396
rect 9867 68347 9909 68356
rect 9771 67892 9813 67901
rect 9771 67852 9772 67892
rect 9812 67852 9813 67892
rect 9771 67843 9813 67852
rect 9772 67649 9812 67734
rect 9676 67591 9716 67600
rect 9771 67640 9813 67649
rect 9771 67600 9772 67640
rect 9812 67600 9813 67640
rect 9771 67591 9813 67600
rect 9868 67472 9908 68347
rect 9676 67432 9908 67472
rect 9676 67136 9716 67432
rect 9676 67087 9716 67096
rect 9771 64616 9813 64625
rect 9771 64576 9772 64616
rect 9812 64576 9813 64616
rect 9771 64567 9813 64576
rect 9868 64616 9908 64625
rect 9964 64616 10004 68431
rect 10059 67808 10101 67817
rect 10059 67768 10060 67808
rect 10100 67768 10101 67808
rect 10156 67808 10196 68935
rect 10252 68489 10292 69952
rect 10347 68984 10389 68993
rect 10347 68944 10348 68984
rect 10388 68944 10389 68984
rect 10347 68935 10389 68944
rect 10348 68850 10388 68935
rect 10251 68480 10293 68489
rect 10251 68440 10252 68480
rect 10292 68440 10293 68480
rect 10251 68431 10293 68440
rect 10444 67985 10484 70120
rect 10539 70120 10540 70160
rect 10580 70120 10581 70160
rect 10539 70111 10581 70120
rect 10443 67976 10485 67985
rect 10443 67936 10444 67976
rect 10484 67936 10485 67976
rect 10443 67927 10485 67936
rect 10156 67768 10292 67808
rect 10059 67759 10101 67768
rect 10060 66968 10100 67759
rect 10252 67724 10292 67768
rect 10156 67640 10196 67649
rect 10156 66977 10196 67600
rect 10060 66919 10100 66928
rect 10155 66968 10197 66977
rect 10155 66928 10156 66968
rect 10196 66928 10197 66968
rect 10155 66919 10197 66928
rect 10252 66800 10292 67684
rect 10444 67640 10484 67927
rect 10540 67817 10580 70111
rect 10636 69908 10676 69917
rect 10636 69245 10676 69868
rect 10731 69908 10773 69917
rect 10731 69868 10732 69908
rect 10772 69868 10773 69908
rect 10731 69859 10773 69868
rect 10732 69774 10772 69859
rect 10635 69236 10677 69245
rect 10635 69196 10636 69236
rect 10676 69196 10677 69236
rect 10635 69187 10677 69196
rect 10731 69152 10773 69161
rect 10731 69112 10732 69152
rect 10772 69112 10773 69152
rect 10731 69103 10773 69112
rect 10732 69018 10772 69103
rect 10635 68984 10677 68993
rect 10635 68944 10636 68984
rect 10676 68944 10677 68984
rect 10635 68935 10677 68944
rect 10636 68480 10676 68935
rect 10636 68431 10676 68440
rect 10731 68480 10773 68489
rect 10731 68440 10732 68480
rect 10772 68440 10773 68480
rect 10731 68431 10773 68440
rect 10732 68346 10772 68431
rect 10828 67985 10868 73060
rect 10923 73016 10965 73025
rect 10923 72976 10924 73016
rect 10964 72976 10965 73016
rect 10923 72967 10965 72976
rect 10924 70076 10964 72967
rect 11020 72941 11060 75496
rect 11116 73697 11156 82048
rect 11596 81920 11636 85936
rect 11500 81880 11636 81920
rect 11211 81836 11253 81845
rect 11211 81796 11212 81836
rect 11252 81796 11253 81836
rect 11211 81787 11253 81796
rect 11212 77468 11252 81787
rect 11307 79988 11349 79997
rect 11307 79948 11308 79988
rect 11348 79948 11349 79988
rect 11307 79939 11349 79948
rect 11308 79157 11348 79939
rect 11403 79400 11445 79409
rect 11403 79360 11404 79400
rect 11444 79360 11445 79400
rect 11403 79351 11445 79360
rect 11307 79148 11349 79157
rect 11307 79108 11308 79148
rect 11348 79108 11349 79148
rect 11307 79099 11349 79108
rect 11404 79064 11444 79351
rect 11404 79015 11444 79024
rect 11307 78980 11349 78989
rect 11307 78940 11308 78980
rect 11348 78940 11349 78980
rect 11307 78931 11349 78940
rect 11308 78846 11348 78931
rect 11212 77428 11348 77468
rect 11211 76460 11253 76469
rect 11211 76420 11212 76460
rect 11252 76420 11253 76460
rect 11211 76411 11253 76420
rect 11115 73688 11157 73697
rect 11115 73648 11116 73688
rect 11156 73648 11157 73688
rect 11115 73639 11157 73648
rect 11019 72932 11061 72941
rect 11019 72892 11020 72932
rect 11060 72892 11061 72932
rect 11019 72883 11061 72892
rect 11020 72689 11060 72883
rect 11019 72680 11061 72689
rect 11019 72640 11020 72680
rect 11060 72640 11061 72680
rect 11019 72631 11061 72640
rect 11115 71588 11157 71597
rect 11115 71548 11116 71588
rect 11156 71548 11157 71588
rect 11115 71539 11157 71548
rect 10924 70036 11060 70076
rect 10923 69908 10965 69917
rect 10923 69868 10924 69908
rect 10964 69868 10965 69908
rect 10923 69859 10965 69868
rect 10924 68489 10964 69859
rect 10923 68480 10965 68489
rect 10923 68440 10924 68480
rect 10964 68440 10965 68480
rect 10923 68431 10965 68440
rect 10827 67976 10869 67985
rect 10827 67936 10828 67976
rect 10868 67936 10869 67976
rect 10827 67927 10869 67936
rect 10539 67808 10581 67817
rect 10924 67808 10964 68431
rect 10539 67768 10540 67808
rect 10580 67768 10581 67808
rect 10539 67759 10581 67768
rect 10828 67768 10964 67808
rect 10732 67640 10772 67649
rect 10444 67600 10732 67640
rect 10732 67591 10772 67600
rect 9908 64576 10004 64616
rect 10156 66760 10292 66800
rect 9772 64482 9812 64567
rect 9580 64240 9812 64280
rect 9772 61769 9812 64240
rect 9483 61760 9525 61769
rect 9483 61720 9484 61760
rect 9524 61720 9525 61760
rect 9483 61711 9525 61720
rect 9771 61760 9813 61769
rect 9771 61720 9772 61760
rect 9812 61720 9813 61760
rect 9771 61711 9813 61720
rect 9771 61172 9813 61181
rect 9771 61132 9772 61172
rect 9812 61132 9813 61172
rect 9771 61123 9813 61132
rect 9387 59744 9429 59753
rect 9387 59704 9388 59744
rect 9428 59704 9429 59744
rect 9387 59695 9429 59704
rect 9675 59660 9717 59669
rect 9675 59620 9676 59660
rect 9716 59620 9717 59660
rect 9675 59611 9717 59620
rect 9292 59492 9332 59501
rect 9332 59452 9524 59492
rect 9292 59443 9332 59452
rect 9484 59408 9524 59452
rect 9580 59408 9620 59417
rect 9484 59368 9580 59408
rect 9580 59359 9620 59368
rect 9676 59408 9716 59611
rect 9676 59359 9716 59368
rect 9772 59240 9812 61123
rect 9868 59921 9908 64576
rect 9963 64364 10005 64373
rect 9963 64324 9964 64364
rect 10004 64324 10005 64364
rect 9963 64315 10005 64324
rect 9964 61601 10004 64315
rect 10059 63860 10101 63869
rect 10059 63820 10060 63860
rect 10100 63820 10101 63860
rect 10059 63811 10101 63820
rect 10060 63449 10100 63811
rect 10059 63440 10101 63449
rect 10059 63400 10060 63440
rect 10100 63400 10101 63440
rect 10059 63391 10101 63400
rect 10060 63113 10100 63391
rect 10059 63104 10101 63113
rect 10059 63064 10060 63104
rect 10100 63064 10101 63104
rect 10059 63055 10101 63064
rect 9963 61592 10005 61601
rect 9963 61552 9964 61592
rect 10004 61552 10005 61592
rect 9963 61543 10005 61552
rect 10060 61592 10100 63055
rect 10060 61543 10100 61552
rect 10059 60920 10101 60929
rect 10059 60880 10060 60920
rect 10100 60880 10101 60920
rect 10059 60871 10101 60880
rect 10060 60786 10100 60871
rect 9867 59912 9909 59921
rect 9867 59872 9868 59912
rect 9908 59872 9909 59912
rect 9867 59863 9909 59872
rect 9676 59200 9812 59240
rect 9291 58904 9333 58913
rect 9291 58864 9292 58904
rect 9332 58864 9333 58904
rect 9291 58855 9333 58864
rect 9292 58484 9332 58855
rect 9387 58736 9429 58745
rect 9387 58696 9388 58736
rect 9428 58696 9429 58736
rect 9387 58687 9429 58696
rect 9292 58435 9332 58444
rect 9388 57476 9428 58687
rect 9676 57728 9716 59200
rect 9868 58745 9908 59863
rect 9963 59744 10005 59753
rect 9963 59704 9964 59744
rect 10004 59704 10005 59744
rect 9963 59695 10005 59704
rect 9964 58913 10004 59695
rect 10060 59324 10100 59335
rect 10060 59249 10100 59284
rect 10156 59324 10196 66760
rect 10731 66464 10773 66473
rect 10731 66424 10732 66464
rect 10772 66424 10773 66464
rect 10731 66415 10773 66424
rect 10347 66128 10389 66137
rect 10732 66128 10772 66415
rect 10828 66389 10868 67768
rect 10923 67640 10965 67649
rect 10923 67600 10924 67640
rect 10964 67600 10965 67640
rect 10923 67591 10965 67600
rect 10827 66380 10869 66389
rect 10827 66340 10828 66380
rect 10868 66340 10869 66380
rect 10827 66331 10869 66340
rect 10347 66088 10348 66128
rect 10388 66088 10389 66128
rect 10347 66079 10389 66088
rect 10444 66088 10732 66128
rect 10251 65540 10293 65549
rect 10251 65500 10252 65540
rect 10292 65500 10293 65540
rect 10251 65491 10293 65500
rect 10252 64700 10292 65491
rect 10348 65456 10388 66079
rect 10444 65717 10484 66088
rect 10732 66079 10772 66088
rect 10540 65960 10580 65969
rect 10580 65920 10868 65960
rect 10540 65911 10580 65920
rect 10443 65708 10485 65717
rect 10443 65668 10444 65708
rect 10484 65668 10485 65708
rect 10443 65659 10485 65668
rect 10828 65456 10868 65920
rect 10388 65416 10484 65456
rect 10348 65407 10388 65416
rect 10347 65288 10389 65297
rect 10347 65248 10348 65288
rect 10388 65248 10389 65288
rect 10347 65239 10389 65248
rect 10252 63272 10292 64660
rect 10348 64700 10388 65239
rect 10348 64651 10388 64660
rect 10444 64280 10484 65416
rect 10828 65407 10868 65416
rect 10924 65456 10964 67591
rect 10539 65204 10581 65213
rect 10539 65164 10540 65204
rect 10580 65164 10581 65204
rect 10539 65155 10581 65164
rect 10540 65070 10580 65155
rect 10827 64616 10869 64625
rect 10827 64576 10828 64616
rect 10868 64576 10869 64616
rect 10827 64567 10869 64576
rect 10828 64482 10868 64567
rect 10924 64280 10964 65416
rect 11020 64709 11060 70036
rect 11116 69992 11156 71539
rect 11212 70169 11252 76411
rect 11211 70160 11253 70169
rect 11211 70120 11212 70160
rect 11252 70120 11253 70160
rect 11211 70111 11253 70120
rect 11212 69992 11252 70001
rect 11116 69952 11212 69992
rect 11116 69329 11156 69952
rect 11212 69943 11252 69952
rect 11115 69320 11157 69329
rect 11115 69280 11116 69320
rect 11156 69280 11157 69320
rect 11115 69271 11157 69280
rect 11212 69320 11252 69329
rect 11308 69320 11348 77428
rect 11500 76880 11540 81880
rect 11788 79316 11828 85936
rect 11980 83273 12020 85936
rect 12172 84449 12212 85936
rect 12171 84440 12213 84449
rect 12171 84400 12172 84440
rect 12212 84400 12213 84440
rect 12171 84391 12213 84400
rect 11979 83264 12021 83273
rect 11979 83224 11980 83264
rect 12020 83224 12021 83264
rect 11979 83215 12021 83224
rect 12364 82508 12404 85936
rect 12172 82468 12404 82508
rect 12172 81920 12212 82468
rect 12556 81920 12596 85936
rect 12748 82013 12788 85936
rect 12747 82004 12789 82013
rect 12747 81964 12748 82004
rect 12788 81964 12789 82004
rect 12747 81955 12789 81964
rect 11404 76840 11540 76880
rect 11596 79276 11828 79316
rect 11884 81880 12212 81920
rect 12364 81880 12596 81920
rect 11404 76721 11444 76840
rect 11403 76712 11445 76721
rect 11403 76672 11404 76712
rect 11444 76672 11445 76712
rect 11403 76663 11445 76672
rect 11500 76712 11540 76721
rect 11596 76712 11636 79276
rect 11691 79148 11733 79157
rect 11691 79108 11692 79148
rect 11732 79108 11733 79148
rect 11691 79099 11733 79108
rect 11540 76672 11636 76712
rect 11692 78224 11732 79099
rect 11884 79064 11924 81880
rect 11979 79820 12021 79829
rect 11979 79780 11980 79820
rect 12020 79780 12021 79820
rect 11979 79771 12021 79780
rect 12267 79820 12309 79829
rect 12267 79780 12268 79820
rect 12308 79780 12309 79820
rect 12267 79771 12309 79780
rect 11884 79015 11924 79024
rect 11500 76663 11540 76672
rect 11499 76040 11541 76049
rect 11499 76000 11500 76040
rect 11540 76000 11541 76040
rect 11692 76040 11732 78184
rect 11980 78065 12020 79771
rect 12171 79736 12213 79745
rect 12171 79696 12172 79736
rect 12212 79696 12213 79736
rect 12171 79687 12213 79696
rect 12268 79736 12308 79771
rect 11979 78056 12021 78065
rect 11979 78016 11980 78056
rect 12020 78016 12021 78056
rect 11979 78007 12021 78016
rect 11884 77552 11924 77561
rect 11980 77552 12020 78007
rect 11924 77512 12020 77552
rect 11884 76301 11924 77512
rect 12076 77300 12116 77309
rect 12076 76796 12116 77260
rect 12028 76756 12116 76796
rect 12028 76754 12068 76756
rect 12028 76705 12068 76714
rect 12172 76712 12212 79687
rect 12268 79685 12308 79696
rect 12364 79148 12404 81880
rect 12940 81257 12980 85936
rect 12939 81248 12981 81257
rect 12939 81208 12940 81248
rect 12980 81208 12981 81248
rect 12939 81199 12981 81208
rect 12268 79108 12404 79148
rect 12460 79568 12500 79577
rect 12268 76880 12308 79108
rect 12460 79064 12500 79528
rect 12747 79400 12789 79409
rect 12747 79360 12748 79400
rect 12788 79360 12789 79400
rect 12747 79351 12789 79360
rect 12556 79148 12596 79157
rect 12596 79108 12692 79148
rect 12556 79099 12596 79108
rect 12412 79054 12500 79064
rect 12452 79024 12500 79054
rect 12412 79005 12452 79014
rect 12268 76840 12500 76880
rect 12172 76672 12308 76712
rect 12171 76544 12213 76553
rect 12171 76504 12172 76544
rect 12212 76504 12213 76544
rect 12171 76495 12213 76504
rect 12172 76410 12212 76495
rect 11883 76292 11925 76301
rect 11883 76252 11884 76292
rect 11924 76252 11925 76292
rect 11883 76243 11925 76252
rect 12171 76292 12213 76301
rect 12171 76252 12172 76292
rect 12212 76252 12213 76292
rect 12171 76243 12213 76252
rect 11979 76208 12021 76217
rect 11979 76168 11980 76208
rect 12020 76168 12021 76208
rect 11979 76159 12021 76168
rect 11692 76000 11828 76040
rect 11499 75991 11541 76000
rect 11500 75906 11540 75991
rect 11691 75872 11733 75881
rect 11691 75832 11692 75872
rect 11732 75832 11733 75872
rect 11691 75823 11733 75832
rect 11595 75200 11637 75209
rect 11595 75160 11596 75200
rect 11636 75160 11637 75200
rect 11595 75151 11637 75160
rect 11403 75032 11445 75041
rect 11403 74992 11404 75032
rect 11444 74992 11445 75032
rect 11403 74983 11445 74992
rect 11404 73688 11444 74983
rect 11499 74696 11541 74705
rect 11499 74656 11500 74696
rect 11540 74656 11541 74696
rect 11499 74647 11541 74656
rect 11404 73639 11444 73648
rect 11500 73688 11540 74647
rect 11500 73639 11540 73648
rect 11499 73436 11541 73445
rect 11499 73396 11500 73436
rect 11540 73396 11541 73436
rect 11499 73387 11541 73396
rect 11403 73016 11445 73025
rect 11403 72976 11404 73016
rect 11444 72976 11445 73016
rect 11403 72967 11445 72976
rect 11252 69280 11348 69320
rect 11212 69271 11252 69280
rect 11211 68480 11253 68489
rect 11211 68440 11212 68480
rect 11252 68440 11253 68480
rect 11211 68431 11253 68440
rect 11116 68396 11156 68405
rect 11116 65549 11156 68356
rect 11212 68346 11252 68431
rect 11260 67682 11300 67691
rect 11300 67642 11348 67654
rect 11260 67614 11348 67642
rect 11211 67556 11253 67565
rect 11211 67516 11212 67556
rect 11252 67516 11253 67556
rect 11211 67507 11253 67516
rect 11212 66968 11252 67507
rect 11308 67388 11348 67614
rect 11404 67556 11444 72967
rect 11500 67556 11540 73387
rect 11596 73016 11636 75151
rect 11596 72437 11636 72976
rect 11595 72428 11637 72437
rect 11595 72388 11596 72428
rect 11636 72388 11637 72428
rect 11595 72379 11637 72388
rect 11596 72176 11636 72379
rect 11596 72017 11636 72136
rect 11595 72008 11637 72017
rect 11595 71968 11596 72008
rect 11636 71968 11637 72008
rect 11595 71959 11637 71968
rect 11692 71588 11732 75823
rect 11788 74033 11828 76000
rect 11883 74360 11925 74369
rect 11883 74320 11884 74360
rect 11924 74320 11925 74360
rect 11883 74311 11925 74320
rect 11787 74024 11829 74033
rect 11787 73984 11788 74024
rect 11828 73984 11829 74024
rect 11787 73975 11829 73984
rect 11788 73445 11828 73975
rect 11884 73772 11924 74311
rect 11980 74285 12020 76159
rect 12075 75200 12117 75209
rect 12075 75160 12076 75200
rect 12116 75160 12117 75200
rect 12075 75151 12117 75160
rect 12076 75066 12116 75151
rect 12075 74696 12117 74705
rect 12075 74656 12076 74696
rect 12116 74656 12117 74696
rect 12075 74647 12117 74656
rect 11979 74276 12021 74285
rect 11979 74236 11980 74276
rect 12020 74236 12021 74276
rect 11979 74227 12021 74236
rect 11979 73856 12021 73865
rect 11979 73816 11980 73856
rect 12020 73816 12021 73856
rect 11979 73807 12021 73816
rect 11884 73723 11924 73732
rect 11980 73772 12020 73807
rect 12076 73772 12116 74647
rect 12172 74528 12212 76243
rect 12268 76217 12308 76672
rect 12267 76208 12309 76217
rect 12267 76168 12268 76208
rect 12308 76168 12309 76208
rect 12267 76159 12309 76168
rect 12268 75032 12308 75041
rect 12268 74537 12308 74992
rect 12172 74479 12212 74488
rect 12267 74528 12309 74537
rect 12267 74488 12268 74528
rect 12308 74488 12309 74528
rect 12267 74479 12309 74488
rect 12267 74276 12309 74285
rect 12267 74236 12268 74276
rect 12308 74236 12309 74276
rect 12267 74227 12309 74236
rect 12364 74276 12404 74285
rect 12076 73732 12212 73772
rect 11980 73721 12020 73732
rect 11979 73604 12021 73613
rect 11979 73564 11980 73604
rect 12020 73564 12021 73604
rect 11979 73555 12021 73564
rect 11787 73436 11829 73445
rect 11787 73396 11788 73436
rect 11828 73396 11829 73436
rect 11787 73387 11829 73396
rect 11787 72764 11829 72773
rect 11787 72724 11788 72764
rect 11828 72724 11829 72764
rect 11787 72715 11829 72724
rect 11788 72630 11828 72715
rect 11980 72176 12020 73555
rect 12076 73016 12116 73025
rect 12076 72857 12116 72976
rect 12172 73016 12212 73732
rect 12075 72848 12117 72857
rect 12075 72808 12076 72848
rect 12116 72808 12117 72848
rect 12075 72799 12117 72808
rect 11980 72127 12020 72136
rect 11788 72008 11828 72017
rect 11828 71968 12020 72008
rect 11788 71959 11828 71968
rect 11692 71548 11924 71588
rect 11596 70673 11636 70758
rect 11595 70664 11637 70673
rect 11595 70624 11596 70664
rect 11636 70624 11637 70664
rect 11595 70615 11637 70624
rect 11788 70496 11828 70505
rect 11788 69992 11828 70456
rect 11884 70160 11924 71548
rect 11980 71504 12020 71968
rect 11980 71455 12020 71464
rect 12076 71504 12116 71513
rect 12172 71504 12212 72976
rect 12116 71464 12212 71504
rect 11979 71168 12021 71177
rect 11979 71128 11980 71168
rect 12020 71128 12021 71168
rect 11979 71119 12021 71128
rect 11980 71009 12020 71119
rect 11979 71000 12021 71009
rect 11979 70960 11980 71000
rect 12020 70960 12021 71000
rect 11979 70951 12021 70960
rect 11980 70664 12020 70951
rect 11980 70615 12020 70624
rect 11884 70111 11924 70120
rect 11740 69982 11828 69992
rect 11780 69952 11828 69982
rect 11740 69933 11780 69942
rect 11883 69152 11925 69161
rect 11883 69112 11884 69152
rect 11924 69112 11925 69152
rect 11883 69103 11925 69112
rect 11884 69018 11924 69103
rect 11692 68480 11732 68489
rect 11692 68321 11732 68440
rect 11691 68312 11733 68321
rect 11691 68272 11692 68312
rect 11732 68272 11733 68312
rect 11691 68263 11733 68272
rect 11595 68144 11637 68153
rect 11595 68104 11596 68144
rect 11636 68104 11637 68144
rect 11595 68095 11637 68104
rect 11596 67892 11636 68095
rect 11596 67843 11636 67852
rect 11787 67808 11829 67817
rect 11787 67768 11788 67808
rect 11828 67768 11829 67808
rect 11787 67759 11829 67768
rect 11788 67640 11828 67759
rect 11788 67591 11828 67600
rect 11500 67516 11732 67556
rect 11404 67507 11444 67516
rect 11308 67348 11540 67388
rect 11500 67136 11540 67348
rect 11500 67087 11540 67096
rect 11308 66968 11348 66977
rect 11692 66968 11732 67516
rect 11788 66968 11828 66977
rect 11212 66928 11308 66968
rect 11115 65540 11157 65549
rect 11115 65500 11116 65540
rect 11156 65500 11157 65540
rect 11115 65491 11157 65500
rect 11019 64700 11061 64709
rect 11019 64660 11020 64700
rect 11060 64660 11061 64700
rect 11019 64651 11061 64660
rect 10348 64240 10484 64280
rect 10732 64240 10964 64280
rect 11020 64280 11060 64651
rect 11212 64373 11252 66928
rect 11308 66919 11348 66928
rect 11596 66928 11788 66968
rect 11499 66212 11541 66221
rect 11499 66172 11500 66212
rect 11540 66172 11541 66212
rect 11499 66163 11541 66172
rect 11307 65540 11349 65549
rect 11307 65500 11308 65540
rect 11348 65500 11349 65540
rect 11307 65491 11349 65500
rect 11308 65456 11348 65491
rect 11308 65405 11348 65416
rect 11403 65456 11445 65465
rect 11403 65416 11404 65456
rect 11444 65416 11445 65456
rect 11403 65407 11445 65416
rect 11307 65204 11349 65213
rect 11307 65164 11308 65204
rect 11348 65164 11349 65204
rect 11307 65155 11349 65164
rect 11308 64630 11348 65155
rect 11308 64581 11348 64590
rect 11211 64364 11253 64373
rect 11211 64324 11212 64364
rect 11252 64324 11253 64364
rect 11211 64315 11253 64324
rect 11020 64240 11156 64280
rect 10348 63944 10388 64240
rect 10348 63869 10388 63904
rect 10347 63860 10389 63869
rect 10347 63820 10348 63860
rect 10388 63820 10389 63860
rect 10347 63811 10389 63820
rect 10539 63776 10581 63785
rect 10539 63736 10540 63776
rect 10580 63736 10581 63776
rect 10539 63727 10581 63736
rect 10443 63692 10485 63701
rect 10443 63652 10444 63692
rect 10484 63652 10485 63692
rect 10443 63643 10485 63652
rect 10444 63356 10484 63643
rect 10540 63642 10580 63727
rect 10635 63524 10677 63533
rect 10635 63484 10636 63524
rect 10676 63484 10677 63524
rect 10635 63475 10677 63484
rect 10444 63307 10484 63316
rect 10252 63232 10388 63272
rect 10251 63104 10293 63113
rect 10251 63064 10252 63104
rect 10292 63064 10293 63104
rect 10251 63055 10293 63064
rect 10252 62970 10292 63055
rect 10251 61760 10293 61769
rect 10251 61720 10252 61760
rect 10292 61720 10293 61760
rect 10251 61711 10293 61720
rect 10252 61626 10292 61711
rect 10348 61685 10388 63232
rect 10539 63188 10581 63197
rect 10539 63148 10540 63188
rect 10580 63148 10581 63188
rect 10539 63139 10581 63148
rect 10540 62936 10580 63139
rect 10636 63104 10676 63475
rect 10732 63197 10772 64240
rect 11019 64028 11061 64037
rect 11019 63988 11020 64028
rect 11060 63988 11061 64028
rect 11019 63979 11061 63988
rect 10828 63944 10868 63953
rect 10828 63701 10868 63904
rect 10924 63944 10964 63953
rect 10827 63692 10869 63701
rect 10827 63652 10828 63692
rect 10868 63652 10869 63692
rect 10827 63643 10869 63652
rect 10731 63188 10773 63197
rect 10924 63188 10964 63904
rect 11020 63785 11060 63979
rect 11019 63776 11061 63785
rect 11019 63736 11020 63776
rect 11060 63736 11061 63776
rect 11019 63727 11061 63736
rect 10731 63148 10732 63188
rect 10772 63148 10773 63188
rect 10731 63139 10773 63148
rect 10828 63148 10964 63188
rect 10636 63055 10676 63064
rect 10731 63020 10773 63029
rect 10731 62980 10732 63020
rect 10772 62980 10773 63020
rect 10731 62971 10773 62980
rect 10540 62896 10676 62936
rect 10443 61844 10485 61853
rect 10443 61804 10444 61844
rect 10484 61804 10485 61844
rect 10443 61795 10485 61804
rect 10347 61676 10389 61685
rect 10347 61636 10348 61676
rect 10388 61636 10389 61676
rect 10347 61627 10389 61636
rect 10251 61340 10293 61349
rect 10251 61300 10252 61340
rect 10292 61300 10293 61340
rect 10251 61291 10293 61300
rect 10252 59669 10292 61291
rect 10444 60668 10484 61795
rect 10539 61760 10581 61769
rect 10539 61720 10540 61760
rect 10580 61720 10581 61760
rect 10539 61711 10581 61720
rect 10540 61611 10580 61711
rect 10540 61562 10580 61571
rect 10636 61592 10676 62896
rect 10636 61508 10676 61552
rect 10540 61468 10676 61508
rect 10540 61349 10580 61468
rect 10732 61424 10772 62971
rect 10636 61384 10772 61424
rect 10539 61340 10581 61349
rect 10539 61300 10540 61340
rect 10580 61300 10581 61340
rect 10539 61291 10581 61300
rect 10539 61088 10581 61097
rect 10539 61048 10540 61088
rect 10580 61048 10581 61088
rect 10539 61039 10581 61048
rect 10540 60845 10580 61039
rect 10539 60836 10581 60845
rect 10539 60796 10540 60836
rect 10580 60796 10581 60836
rect 10539 60787 10581 60796
rect 10444 60628 10580 60668
rect 10347 60584 10389 60593
rect 10347 60544 10348 60584
rect 10388 60544 10389 60584
rect 10347 60535 10389 60544
rect 10251 59660 10293 59669
rect 10251 59620 10252 59660
rect 10292 59620 10293 59660
rect 10251 59611 10293 59620
rect 10196 59284 10292 59324
rect 10156 59275 10196 59284
rect 10059 59240 10101 59249
rect 10059 59200 10060 59240
rect 10100 59200 10101 59240
rect 10059 59191 10101 59200
rect 9963 58904 10005 58913
rect 9963 58864 9964 58904
rect 10004 58864 10005 58904
rect 9963 58855 10005 58864
rect 9867 58736 9909 58745
rect 9867 58696 9868 58736
rect 9908 58696 9909 58736
rect 9867 58687 9909 58696
rect 9963 58568 10005 58577
rect 9963 58528 9964 58568
rect 10004 58528 10005 58568
rect 9963 58519 10005 58528
rect 9964 58434 10004 58519
rect 10155 58484 10197 58493
rect 10155 58444 10156 58484
rect 10196 58444 10197 58484
rect 10155 58435 10197 58444
rect 9867 57980 9909 57989
rect 9867 57940 9868 57980
rect 9908 57940 9909 57980
rect 9867 57931 9909 57940
rect 9772 57854 9812 57863
rect 9772 57812 9812 57814
rect 9868 57812 9908 57931
rect 9772 57772 9908 57812
rect 9676 57688 9812 57728
rect 9388 57436 9716 57476
rect 9580 57056 9620 57065
rect 9292 56972 9332 56981
rect 9580 56972 9620 57016
rect 9676 57056 9716 57436
rect 9676 57007 9716 57016
rect 9332 56932 9620 56972
rect 9292 56923 9332 56932
rect 9483 56804 9525 56813
rect 9483 56764 9484 56804
rect 9524 56764 9525 56804
rect 9483 56755 9525 56764
rect 9484 56309 9524 56755
rect 9675 56384 9717 56393
rect 9675 56344 9676 56384
rect 9716 56344 9717 56384
rect 9675 56335 9717 56344
rect 9483 56300 9525 56309
rect 9483 56260 9484 56300
rect 9524 56260 9525 56300
rect 9483 56251 9525 56260
rect 9291 56132 9333 56141
rect 9291 56092 9292 56132
rect 9332 56092 9333 56132
rect 9291 56083 9333 56092
rect 9292 53537 9332 56083
rect 9484 54872 9524 56251
rect 9676 55301 9716 56335
rect 9675 55292 9717 55301
rect 9675 55252 9676 55292
rect 9716 55252 9717 55292
rect 9675 55243 9717 55252
rect 9388 54832 9484 54872
rect 9291 53528 9333 53537
rect 9291 53488 9292 53528
rect 9332 53488 9333 53528
rect 9291 53479 9333 53488
rect 9388 53369 9428 54832
rect 9484 54823 9524 54832
rect 9676 54797 9716 55243
rect 9675 54788 9717 54797
rect 9675 54748 9676 54788
rect 9716 54748 9717 54788
rect 9675 54739 9717 54748
rect 9676 54620 9716 54629
rect 9483 54536 9525 54545
rect 9483 54496 9484 54536
rect 9524 54496 9525 54536
rect 9483 54487 9525 54496
rect 9484 54032 9524 54487
rect 9676 54209 9716 54580
rect 9675 54200 9717 54209
rect 9675 54160 9676 54200
rect 9716 54160 9717 54200
rect 9580 54125 9620 54156
rect 9675 54151 9717 54160
rect 9579 54116 9621 54125
rect 9579 54076 9580 54116
rect 9620 54076 9621 54116
rect 9579 54067 9621 54076
rect 9387 53360 9429 53369
rect 9387 53320 9388 53360
rect 9428 53320 9429 53360
rect 9387 53311 9429 53320
rect 9484 53192 9524 53992
rect 9580 54032 9620 54067
rect 9580 53789 9620 53992
rect 9675 54032 9717 54041
rect 9675 53992 9676 54032
rect 9716 53992 9717 54032
rect 9675 53983 9717 53992
rect 9579 53780 9621 53789
rect 9579 53740 9580 53780
rect 9620 53740 9621 53780
rect 9579 53731 9621 53740
rect 9292 53152 9524 53192
rect 9195 51680 9237 51689
rect 9195 51640 9196 51680
rect 9236 51640 9237 51680
rect 9195 51631 9237 51640
rect 9292 51101 9332 53152
rect 9676 53117 9716 53983
rect 9675 53108 9717 53117
rect 9675 53068 9676 53108
rect 9716 53068 9717 53108
rect 9675 53059 9717 53068
rect 9772 52688 9812 57688
rect 9868 56141 9908 57772
rect 10059 57140 10101 57149
rect 10059 57100 10060 57140
rect 10100 57100 10101 57140
rect 10059 57091 10101 57100
rect 10156 57140 10196 58435
rect 10156 57091 10196 57100
rect 10060 57006 10100 57091
rect 9867 56132 9909 56141
rect 9867 56092 9868 56132
rect 9908 56092 9909 56132
rect 9867 56083 9909 56092
rect 10059 55712 10101 55721
rect 10059 55672 10060 55712
rect 10100 55672 10101 55712
rect 10059 55663 10101 55672
rect 10060 55578 10100 55663
rect 10252 55553 10292 59284
rect 10348 58829 10388 60535
rect 10443 60080 10485 60089
rect 10443 60040 10444 60080
rect 10484 60040 10485 60080
rect 10443 60031 10485 60040
rect 10347 58820 10389 58829
rect 10347 58780 10348 58820
rect 10388 58780 10389 58820
rect 10347 58771 10389 58780
rect 10444 58493 10484 60031
rect 10443 58484 10485 58493
rect 10443 58444 10444 58484
rect 10484 58444 10485 58484
rect 10443 58435 10485 58444
rect 10347 55712 10389 55721
rect 10347 55672 10348 55712
rect 10388 55672 10389 55712
rect 10347 55663 10389 55672
rect 9868 55544 9908 55553
rect 9868 55049 9908 55504
rect 10251 55544 10293 55553
rect 10251 55504 10252 55544
rect 10292 55504 10293 55544
rect 10251 55495 10293 55504
rect 10348 55544 10388 55663
rect 10348 55495 10388 55504
rect 10444 55544 10484 55553
rect 9867 55040 9909 55049
rect 9867 55000 9868 55040
rect 9908 55000 9909 55040
rect 9867 54991 9909 55000
rect 10155 54956 10197 54965
rect 10155 54916 10156 54956
rect 10196 54916 10197 54956
rect 10155 54907 10197 54916
rect 10060 54872 10100 54881
rect 10060 54293 10100 54832
rect 10156 54872 10196 54907
rect 10156 54821 10196 54832
rect 10251 54872 10293 54881
rect 10251 54832 10252 54872
rect 10292 54832 10293 54872
rect 10251 54823 10293 54832
rect 10348 54872 10388 54881
rect 10252 54738 10292 54823
rect 10155 54704 10197 54713
rect 10155 54664 10156 54704
rect 10196 54664 10197 54704
rect 10155 54655 10197 54664
rect 10059 54284 10101 54293
rect 10059 54244 10060 54284
rect 10100 54244 10101 54284
rect 10059 54235 10101 54244
rect 10060 54041 10100 54126
rect 10059 54032 10101 54041
rect 10059 53992 10060 54032
rect 10100 53992 10101 54032
rect 10059 53983 10101 53992
rect 10156 53864 10196 54655
rect 10060 53824 10196 53864
rect 9963 53780 10005 53789
rect 9963 53740 9964 53780
rect 10004 53740 10005 53780
rect 9963 53731 10005 53740
rect 9867 53024 9909 53033
rect 9867 52984 9868 53024
rect 9908 52984 9909 53024
rect 9867 52975 9909 52984
rect 9388 52648 9812 52688
rect 9291 51092 9333 51101
rect 9291 51052 9292 51092
rect 9332 51052 9333 51092
rect 9291 51043 9333 51052
rect 9099 51008 9141 51017
rect 9099 50968 9100 51008
rect 9140 50968 9141 51008
rect 9099 50959 9141 50968
rect 9100 50874 9140 50959
rect 9195 50756 9237 50765
rect 9195 50716 9196 50756
rect 9236 50716 9237 50756
rect 9195 50707 9237 50716
rect 9196 48161 9236 50707
rect 9291 49328 9333 49337
rect 9291 49288 9292 49328
rect 9332 49288 9333 49328
rect 9291 49279 9333 49288
rect 9292 48824 9332 49279
rect 9195 48152 9237 48161
rect 9195 48112 9196 48152
rect 9236 48112 9237 48152
rect 9195 48103 9237 48112
rect 9292 47825 9332 48784
rect 9291 47816 9333 47825
rect 9291 47776 9292 47816
rect 9332 47776 9333 47816
rect 9291 47767 9333 47776
rect 9292 47489 9332 47767
rect 9291 47480 9333 47489
rect 9291 47440 9292 47480
rect 9332 47440 9333 47480
rect 9291 47431 9333 47440
rect 9100 47228 9140 47239
rect 9100 47153 9140 47188
rect 9196 47228 9236 47237
rect 9388 47228 9428 52648
rect 9580 52520 9620 52529
rect 9580 52361 9620 52480
rect 9579 52352 9621 52361
rect 9579 52312 9580 52352
rect 9620 52312 9621 52352
rect 9579 52303 9621 52312
rect 9772 52352 9812 52361
rect 9628 51017 9668 51026
rect 9772 51008 9812 52312
rect 9868 51857 9908 52975
rect 9867 51848 9909 51857
rect 9867 51808 9868 51848
rect 9908 51808 9909 51848
rect 9867 51799 9909 51808
rect 9868 51714 9908 51799
rect 9668 50977 9812 51008
rect 9628 50968 9812 50977
rect 9771 50840 9813 50849
rect 9771 50800 9772 50840
rect 9812 50800 9813 50840
rect 9771 50791 9813 50800
rect 9772 50706 9812 50791
rect 9484 50429 9524 50460
rect 9483 50420 9525 50429
rect 9483 50380 9484 50420
rect 9524 50380 9525 50420
rect 9483 50371 9525 50380
rect 9484 50336 9524 50371
rect 9484 50261 9524 50296
rect 9483 50252 9525 50261
rect 9483 50212 9484 50252
rect 9524 50212 9525 50252
rect 9483 50203 9525 50212
rect 9676 50084 9716 50093
rect 9716 50044 9812 50084
rect 9676 50035 9716 50044
rect 9580 49496 9620 49505
rect 9484 48992 9524 49001
rect 9580 48992 9620 49456
rect 9524 48952 9620 48992
rect 9676 49496 9716 49505
rect 9484 48943 9524 48952
rect 9676 48320 9716 49456
rect 9772 48824 9812 50044
rect 9772 48775 9812 48784
rect 9868 48824 9908 48833
rect 9868 48320 9908 48784
rect 9580 48280 9908 48320
rect 9388 47188 9524 47228
rect 9099 47144 9141 47153
rect 9099 47104 9100 47144
rect 9140 47104 9141 47144
rect 9196 47144 9236 47188
rect 9196 47104 9428 47144
rect 9099 47095 9141 47104
rect 9291 46892 9333 46901
rect 9291 46852 9292 46892
rect 9332 46852 9333 46892
rect 9291 46843 9333 46852
rect 9195 46640 9237 46649
rect 9195 46600 9196 46640
rect 9236 46600 9237 46640
rect 9195 46591 9237 46600
rect 9196 45800 9236 46591
rect 9100 45760 9196 45800
rect 9100 44465 9140 45760
rect 9196 45751 9236 45760
rect 9195 45128 9237 45137
rect 9195 45088 9196 45128
rect 9236 45088 9237 45128
rect 9195 45079 9237 45088
rect 9099 44456 9141 44465
rect 9099 44416 9100 44456
rect 9140 44416 9141 44456
rect 9099 44407 9141 44416
rect 9099 44288 9141 44297
rect 9099 44248 9100 44288
rect 9140 44248 9141 44288
rect 9099 44239 9141 44248
rect 9196 44288 9236 45079
rect 9292 44969 9332 46843
rect 9388 45716 9428 47104
rect 9484 46229 9524 47188
rect 9483 46220 9525 46229
rect 9483 46180 9484 46220
rect 9524 46180 9525 46220
rect 9483 46171 9525 46180
rect 9580 46061 9620 48280
rect 9675 48152 9717 48161
rect 9675 48112 9676 48152
rect 9716 48112 9717 48152
rect 9675 48103 9717 48112
rect 9676 47312 9716 48103
rect 9867 48068 9909 48077
rect 9867 48028 9868 48068
rect 9908 48028 9909 48068
rect 9867 48019 9909 48028
rect 9868 47984 9908 48019
rect 9868 47933 9908 47944
rect 9676 47263 9716 47272
rect 9964 46556 10004 53731
rect 10060 51092 10100 53824
rect 10348 53528 10388 54832
rect 10156 53488 10388 53528
rect 10156 53369 10196 53488
rect 10155 53360 10197 53369
rect 10155 53320 10156 53360
rect 10196 53320 10197 53360
rect 10155 53311 10197 53320
rect 10252 53360 10292 53371
rect 10252 53285 10292 53320
rect 10251 53276 10293 53285
rect 10444 53276 10484 55504
rect 10540 55040 10580 60628
rect 10636 60509 10676 61384
rect 10828 61097 10868 63148
rect 10923 62936 10965 62945
rect 10923 62896 10924 62936
rect 10964 62896 10965 62936
rect 10923 62887 10965 62896
rect 10924 62432 10964 62887
rect 10924 62383 10964 62392
rect 11116 62180 11156 64240
rect 11404 63944 11444 65407
rect 11500 64532 11540 66163
rect 11500 64483 11540 64492
rect 11307 63860 11349 63869
rect 10924 62140 11156 62180
rect 11212 63820 11308 63860
rect 11348 63820 11349 63860
rect 10827 61088 10869 61097
rect 10827 61048 10828 61088
rect 10868 61048 10869 61088
rect 10827 61039 10869 61048
rect 10732 60920 10772 60929
rect 10635 60500 10677 60509
rect 10635 60460 10636 60500
rect 10676 60460 10677 60500
rect 10635 60451 10677 60460
rect 10636 60332 10676 60341
rect 10732 60332 10772 60880
rect 10828 60920 10868 61039
rect 10828 60871 10868 60880
rect 10827 60752 10869 60761
rect 10827 60712 10828 60752
rect 10868 60712 10869 60752
rect 10827 60703 10869 60712
rect 10676 60292 10772 60332
rect 10636 60283 10676 60292
rect 10636 59408 10676 59417
rect 10636 59165 10676 59368
rect 10635 59156 10677 59165
rect 10635 59116 10636 59156
rect 10676 59116 10677 59156
rect 10635 59107 10677 59116
rect 10636 57056 10676 59107
rect 10636 57007 10676 57016
rect 10828 56729 10868 60703
rect 10924 59249 10964 62140
rect 11115 61844 11157 61853
rect 11115 61804 11116 61844
rect 11156 61804 11157 61844
rect 11115 61795 11157 61804
rect 11116 61676 11156 61795
rect 11116 61625 11156 61636
rect 11019 61592 11061 61601
rect 11019 61552 11020 61592
rect 11060 61552 11061 61592
rect 11019 61543 11061 61552
rect 11020 61458 11060 61543
rect 11212 60845 11252 63820
rect 11307 63811 11349 63820
rect 11308 63726 11348 63811
rect 11404 61853 11444 63904
rect 11403 61844 11445 61853
rect 11403 61804 11404 61844
rect 11444 61804 11445 61844
rect 11403 61795 11445 61804
rect 11404 60920 11444 61795
rect 11596 61760 11636 66928
rect 11788 66919 11828 66928
rect 12076 66809 12116 71464
rect 12268 69161 12308 74227
rect 12364 73949 12404 74236
rect 12363 73940 12405 73949
rect 12363 73900 12364 73940
rect 12404 73900 12405 73940
rect 12363 73891 12405 73900
rect 12460 73688 12500 76840
rect 12652 76133 12692 79108
rect 12748 76637 12788 79351
rect 13132 79325 13172 85936
rect 13227 84860 13269 84869
rect 13227 84820 13228 84860
rect 13268 84820 13269 84860
rect 13227 84811 13269 84820
rect 13228 83768 13268 84811
rect 13324 84449 13364 85936
rect 13323 84440 13365 84449
rect 13323 84400 13324 84440
rect 13364 84400 13365 84440
rect 13323 84391 13365 84400
rect 13324 83768 13364 83777
rect 13228 83728 13324 83768
rect 13324 83719 13364 83728
rect 13516 83684 13556 85936
rect 13708 84449 13748 85936
rect 13900 84449 13940 85936
rect 14092 84533 14132 85936
rect 14091 84524 14133 84533
rect 14091 84484 14092 84524
rect 14132 84484 14133 84524
rect 14091 84475 14133 84484
rect 14284 84449 14324 85936
rect 14476 84953 14516 85936
rect 14475 84944 14517 84953
rect 14475 84904 14476 84944
rect 14516 84904 14517 84944
rect 14475 84895 14517 84904
rect 14668 84617 14708 85936
rect 14667 84608 14709 84617
rect 14667 84568 14668 84608
rect 14708 84568 14709 84608
rect 14667 84559 14709 84568
rect 14860 84533 14900 85936
rect 14859 84524 14901 84533
rect 14859 84484 14860 84524
rect 14900 84484 14901 84524
rect 14859 84475 14901 84484
rect 15052 84449 15092 85936
rect 15244 84449 15284 85936
rect 15436 85625 15476 85936
rect 15435 85616 15477 85625
rect 15435 85576 15436 85616
rect 15476 85576 15477 85616
rect 15435 85567 15477 85576
rect 13707 84440 13749 84449
rect 13707 84400 13708 84440
rect 13748 84400 13749 84440
rect 13707 84391 13749 84400
rect 13899 84440 13941 84449
rect 13899 84400 13900 84440
rect 13940 84400 13941 84440
rect 13899 84391 13941 84400
rect 14283 84440 14325 84449
rect 14283 84400 14284 84440
rect 14324 84400 14325 84440
rect 14283 84391 14325 84400
rect 15051 84440 15093 84449
rect 15051 84400 15052 84440
rect 15092 84400 15093 84440
rect 15051 84391 15093 84400
rect 15243 84440 15285 84449
rect 15243 84400 15244 84440
rect 15284 84400 15285 84440
rect 15243 84391 15285 84400
rect 14955 83768 14997 83777
rect 14955 83728 14956 83768
rect 14996 83728 14997 83768
rect 14955 83719 14997 83728
rect 15532 83768 15572 83777
rect 15628 83768 15668 85936
rect 15723 85868 15765 85877
rect 15723 85828 15724 85868
rect 15764 85828 15765 85868
rect 15723 85819 15765 85828
rect 15572 83728 15668 83768
rect 15724 83768 15764 85819
rect 15532 83719 15572 83728
rect 15724 83719 15764 83728
rect 13516 83644 13652 83684
rect 13515 83516 13557 83525
rect 13515 83476 13516 83516
rect 13556 83476 13557 83516
rect 13515 83467 13557 83476
rect 13516 83382 13556 83467
rect 13612 81920 13652 83644
rect 14956 83634 14996 83719
rect 15147 83516 15189 83525
rect 15147 83476 15148 83516
rect 15188 83476 15189 83516
rect 15147 83467 15189 83476
rect 15340 83516 15380 83525
rect 15148 83382 15188 83467
rect 13899 82844 13941 82853
rect 13899 82804 13900 82844
rect 13940 82804 13941 82844
rect 13899 82795 13941 82804
rect 13516 81880 13652 81920
rect 13227 80576 13269 80585
rect 13227 80536 13228 80576
rect 13268 80536 13364 80576
rect 13227 80527 13269 80536
rect 13228 80442 13268 80527
rect 13131 79316 13173 79325
rect 13131 79276 13132 79316
rect 13172 79276 13173 79316
rect 13131 79267 13173 79276
rect 13132 79064 13172 79073
rect 13132 78476 13172 79024
rect 13132 78427 13172 78436
rect 13228 79064 13268 79073
rect 12940 78224 12980 78235
rect 12940 78149 12980 78184
rect 12939 78140 12981 78149
rect 12939 78100 12940 78140
rect 12980 78100 12981 78140
rect 12939 78091 12981 78100
rect 13036 77552 13076 77561
rect 13036 77225 13076 77512
rect 13035 77216 13077 77225
rect 13035 77176 13036 77216
rect 13076 77176 13077 77216
rect 13035 77167 13077 77176
rect 12843 76880 12885 76889
rect 12843 76840 12844 76880
rect 12884 76840 12885 76880
rect 12843 76831 12885 76840
rect 12747 76628 12789 76637
rect 12747 76588 12748 76628
rect 12788 76588 12789 76628
rect 12747 76579 12789 76588
rect 12747 76292 12789 76301
rect 12747 76252 12748 76292
rect 12788 76252 12789 76292
rect 12747 76243 12789 76252
rect 12651 76124 12693 76133
rect 12651 76084 12652 76124
rect 12692 76084 12693 76124
rect 12651 76075 12693 76084
rect 12748 76040 12788 76243
rect 12748 75991 12788 76000
rect 12747 74696 12789 74705
rect 12747 74656 12748 74696
rect 12788 74656 12789 74696
rect 12747 74647 12789 74656
rect 12651 74528 12693 74537
rect 12651 74488 12652 74528
rect 12692 74488 12693 74528
rect 12651 74479 12693 74488
rect 12748 74528 12788 74647
rect 12748 74479 12788 74488
rect 12652 74394 12692 74479
rect 12555 74360 12597 74369
rect 12555 74320 12556 74360
rect 12596 74320 12597 74360
rect 12555 74311 12597 74320
rect 12460 73445 12500 73648
rect 12459 73436 12501 73445
rect 12459 73396 12460 73436
rect 12500 73396 12501 73436
rect 12459 73387 12501 73396
rect 12556 73100 12596 74311
rect 12747 74192 12789 74201
rect 12747 74152 12748 74192
rect 12788 74152 12789 74192
rect 12747 74143 12789 74152
rect 12651 73856 12693 73865
rect 12651 73816 12652 73856
rect 12692 73816 12693 73856
rect 12651 73807 12693 73816
rect 12460 73060 12596 73100
rect 12460 72932 12500 73060
rect 12556 72932 12596 72941
rect 12460 72892 12556 72932
rect 12363 71420 12405 71429
rect 12363 71380 12364 71420
rect 12404 71380 12405 71420
rect 12363 71371 12405 71380
rect 12460 71420 12500 72892
rect 12556 72883 12596 72892
rect 12652 72932 12692 73807
rect 12652 71840 12692 72892
rect 12748 72185 12788 74143
rect 12747 72176 12789 72185
rect 12747 72136 12748 72176
rect 12788 72136 12789 72176
rect 12747 72127 12789 72136
rect 12267 69152 12309 69161
rect 12267 69112 12268 69152
rect 12308 69112 12309 69152
rect 12267 69103 12309 69112
rect 12172 68466 12212 68475
rect 12172 68153 12212 68426
rect 12171 68144 12213 68153
rect 12171 68104 12172 68144
rect 12212 68104 12213 68144
rect 12171 68095 12213 68104
rect 12075 66800 12117 66809
rect 12075 66760 12076 66800
rect 12116 66760 12117 66800
rect 12075 66751 12117 66760
rect 11980 66137 12020 66222
rect 11979 66128 12021 66137
rect 12268 66128 12308 69103
rect 12364 68648 12404 71371
rect 12460 71345 12500 71380
rect 12556 71800 12692 71840
rect 12556 71420 12596 71800
rect 12459 71336 12501 71345
rect 12459 71296 12460 71336
rect 12500 71296 12501 71336
rect 12459 71287 12501 71296
rect 12556 70412 12596 71380
rect 12651 71000 12693 71009
rect 12651 70960 12652 71000
rect 12692 70960 12693 71000
rect 12651 70951 12693 70960
rect 12364 68599 12404 68608
rect 12460 70372 12596 70412
rect 12364 66128 12404 66137
rect 11979 66088 11980 66128
rect 12020 66088 12021 66128
rect 11979 66079 12021 66088
rect 12076 66088 12364 66128
rect 12076 65960 12116 66088
rect 12364 66079 12404 66088
rect 11788 65920 12116 65960
rect 12172 65960 12212 65969
rect 12212 65920 12404 65960
rect 11788 64112 11828 65920
rect 12172 65911 12212 65920
rect 12267 65708 12309 65717
rect 12267 65668 12268 65708
rect 12308 65668 12309 65708
rect 12267 65659 12309 65668
rect 11692 64072 11828 64112
rect 11884 65456 11924 65465
rect 11692 61769 11732 64072
rect 11787 63944 11829 63953
rect 11884 63944 11924 65416
rect 12268 64616 12308 65659
rect 12364 65451 12404 65920
rect 12364 65402 12404 65411
rect 12364 64616 12404 64625
rect 12268 64576 12364 64616
rect 12364 64280 12404 64576
rect 11787 63904 11788 63944
rect 11828 63904 11884 63944
rect 11787 63895 11829 63904
rect 11884 63895 11924 63904
rect 11980 64240 12404 64280
rect 11500 61720 11636 61760
rect 11691 61760 11733 61769
rect 11691 61720 11692 61760
rect 11732 61720 11733 61760
rect 11500 61433 11540 61720
rect 11691 61711 11733 61720
rect 11596 61592 11636 61601
rect 11788 61592 11828 63895
rect 11883 63440 11925 63449
rect 11883 63400 11884 63440
rect 11924 63400 11925 63440
rect 11883 63391 11925 63400
rect 11884 63104 11924 63391
rect 11884 63055 11924 63064
rect 11636 61552 11828 61592
rect 11499 61424 11541 61433
rect 11499 61384 11500 61424
rect 11540 61384 11541 61424
rect 11499 61375 11541 61384
rect 11308 60880 11444 60920
rect 11596 60920 11636 61552
rect 11788 60920 11828 60929
rect 11596 60880 11788 60920
rect 11828 60880 11924 60920
rect 11211 60836 11253 60845
rect 11211 60796 11212 60836
rect 11252 60796 11253 60836
rect 11211 60787 11253 60796
rect 11308 60836 11348 60880
rect 11788 60871 11828 60880
rect 11212 60702 11252 60787
rect 11308 60761 11348 60796
rect 11307 60752 11349 60761
rect 11307 60712 11308 60752
rect 11348 60712 11349 60752
rect 11307 60703 11349 60712
rect 11500 60080 11540 60091
rect 11500 60005 11540 60040
rect 11499 59996 11541 60005
rect 11499 59956 11500 59996
rect 11540 59956 11541 59996
rect 11499 59947 11541 59956
rect 11403 59660 11445 59669
rect 11308 59620 11404 59660
rect 11444 59620 11445 59660
rect 11308 59576 11348 59620
rect 11403 59611 11445 59620
rect 11308 59527 11348 59536
rect 11116 59394 11156 59403
rect 10923 59240 10965 59249
rect 10923 59200 10924 59240
rect 10964 59200 10965 59240
rect 10923 59191 10965 59200
rect 11019 58988 11061 58997
rect 11019 58948 11020 58988
rect 11060 58948 11061 58988
rect 11019 58939 11061 58948
rect 10923 58484 10965 58493
rect 10923 58444 10924 58484
rect 10964 58444 10965 58484
rect 10923 58435 10965 58444
rect 10924 57905 10964 58435
rect 10923 57896 10965 57905
rect 10923 57856 10924 57896
rect 10964 57856 10965 57896
rect 10923 57847 10965 57856
rect 11020 57896 11060 58939
rect 11116 57980 11156 59354
rect 11212 58568 11252 58579
rect 11212 58493 11252 58528
rect 11692 58568 11732 58577
rect 11211 58484 11253 58493
rect 11211 58444 11212 58484
rect 11252 58444 11253 58484
rect 11211 58435 11253 58444
rect 11404 58484 11444 58493
rect 11692 58484 11732 58528
rect 11787 58568 11829 58577
rect 11787 58528 11788 58568
rect 11828 58528 11829 58568
rect 11787 58519 11829 58528
rect 11444 58444 11732 58484
rect 11404 58435 11444 58444
rect 11788 58434 11828 58519
rect 11884 58316 11924 60880
rect 11692 58276 11924 58316
rect 11212 57980 11252 57989
rect 11116 57940 11212 57980
rect 11212 57931 11252 57940
rect 10635 56720 10677 56729
rect 10635 56680 10636 56720
rect 10676 56680 10677 56720
rect 10635 56671 10677 56680
rect 10827 56720 10869 56729
rect 10827 56680 10828 56720
rect 10868 56680 10869 56720
rect 10827 56671 10869 56680
rect 10636 55217 10676 56671
rect 10924 56384 10964 57847
rect 11020 57812 11060 57856
rect 11020 57772 11252 57812
rect 11116 57061 11156 57070
rect 11019 56636 11061 56645
rect 11019 56596 11020 56636
rect 11060 56596 11061 56636
rect 11019 56587 11061 56596
rect 10924 56309 10964 56344
rect 10923 56300 10965 56309
rect 10923 56260 10924 56300
rect 10964 56260 10965 56300
rect 10923 56251 10965 56260
rect 11020 55973 11060 56587
rect 11116 56552 11156 57021
rect 11212 56804 11252 57772
rect 11403 57392 11445 57401
rect 11403 57352 11404 57392
rect 11444 57352 11445 57392
rect 11403 57343 11445 57352
rect 11320 56981 11360 57000
rect 11308 56972 11360 56981
rect 11404 56972 11444 57343
rect 11348 56932 11444 56972
rect 11308 56923 11348 56932
rect 11212 56764 11348 56804
rect 11116 56503 11156 56512
rect 11019 55964 11061 55973
rect 11019 55924 11020 55964
rect 11060 55924 11061 55964
rect 11019 55915 11061 55924
rect 10924 55628 10964 55637
rect 11020 55628 11060 55915
rect 10964 55588 11060 55628
rect 11211 55628 11253 55637
rect 11211 55588 11212 55628
rect 11252 55588 11253 55628
rect 10924 55579 10964 55588
rect 11211 55579 11253 55588
rect 10828 55544 10868 55553
rect 10828 55460 10868 55504
rect 10828 55420 10964 55460
rect 10635 55208 10677 55217
rect 10635 55168 10636 55208
rect 10676 55168 10677 55208
rect 10635 55159 10677 55168
rect 10827 55208 10869 55217
rect 10827 55168 10828 55208
rect 10868 55168 10869 55208
rect 10827 55159 10869 55168
rect 10540 55000 10676 55040
rect 10540 54872 10580 54883
rect 10540 54797 10580 54832
rect 10539 54788 10581 54797
rect 10539 54748 10540 54788
rect 10580 54748 10581 54788
rect 10539 54739 10581 54748
rect 10539 54200 10581 54209
rect 10539 54160 10540 54200
rect 10580 54160 10581 54200
rect 10539 54151 10581 54160
rect 10251 53236 10252 53276
rect 10292 53236 10293 53276
rect 10251 53227 10293 53236
rect 10348 53236 10484 53276
rect 10540 54037 10580 54151
rect 10155 52940 10197 52949
rect 10348 52940 10388 53236
rect 10540 53117 10580 53997
rect 10155 52900 10156 52940
rect 10196 52900 10388 52940
rect 10444 53108 10484 53117
rect 10155 52891 10197 52900
rect 10444 52772 10484 53068
rect 10539 53108 10581 53117
rect 10539 53068 10540 53108
rect 10580 53068 10581 53108
rect 10539 53059 10581 53068
rect 10348 52732 10484 52772
rect 10348 52613 10388 52732
rect 10347 52604 10389 52613
rect 10347 52564 10348 52604
rect 10388 52564 10389 52604
rect 10347 52562 10389 52564
rect 10347 52555 10348 52562
rect 10156 52520 10196 52531
rect 10156 52445 10196 52480
rect 10252 52520 10292 52529
rect 10388 52555 10389 52562
rect 10348 52513 10388 52522
rect 10636 52520 10676 55000
rect 10731 53864 10773 53873
rect 10731 53824 10732 53864
rect 10772 53824 10773 53864
rect 10731 53815 10773 53824
rect 10732 53730 10772 53815
rect 10828 53528 10868 55159
rect 10924 54209 10964 55420
rect 10923 54200 10965 54209
rect 10923 54160 10924 54200
rect 10964 54160 10965 54200
rect 10923 54151 10965 54160
rect 10924 54032 10964 54041
rect 11212 54032 11252 55579
rect 10964 53992 11156 54032
rect 10924 53983 10964 53992
rect 11020 53864 11060 53873
rect 10732 53488 10868 53528
rect 10924 53824 11020 53864
rect 10732 52949 10772 53488
rect 10827 53360 10869 53369
rect 10827 53320 10828 53360
rect 10868 53320 10869 53360
rect 10827 53311 10869 53320
rect 10924 53360 10964 53824
rect 11020 53815 11060 53824
rect 11116 53528 11156 53992
rect 11212 53957 11252 53992
rect 11211 53948 11253 53957
rect 11211 53908 11212 53948
rect 11252 53908 11253 53948
rect 11211 53899 11253 53908
rect 11212 53868 11252 53899
rect 11308 53528 11348 56764
rect 11404 55544 11444 55553
rect 11404 55460 11444 55504
rect 11692 55460 11732 58276
rect 11883 57980 11925 57989
rect 11883 57940 11884 57980
rect 11924 57940 11925 57980
rect 11883 57931 11925 57940
rect 11884 57896 11924 57931
rect 11884 57845 11924 57856
rect 11883 57728 11925 57737
rect 11883 57688 11884 57728
rect 11924 57688 11925 57728
rect 11883 57679 11925 57688
rect 11884 56384 11924 57679
rect 11980 57065 12020 64240
rect 12364 63953 12404 64034
rect 12363 63944 12405 63953
rect 12363 63899 12364 63944
rect 12404 63899 12405 63944
rect 12363 63895 12405 63899
rect 12364 63890 12404 63895
rect 12076 62936 12116 62945
rect 12076 61606 12116 62896
rect 12076 61557 12116 61566
rect 12172 62432 12212 62441
rect 12172 61349 12212 62392
rect 12364 62180 12404 62189
rect 12267 61676 12309 61685
rect 12267 61636 12268 61676
rect 12308 61636 12309 61676
rect 12267 61627 12309 61636
rect 12268 61508 12308 61627
rect 12268 61459 12308 61468
rect 12171 61340 12213 61349
rect 12171 61300 12172 61340
rect 12212 61300 12213 61340
rect 12171 61291 12213 61300
rect 12172 60836 12212 61291
rect 12364 60920 12404 62140
rect 12460 61760 12500 70372
rect 12555 69320 12597 69329
rect 12555 69280 12556 69320
rect 12596 69280 12597 69320
rect 12555 69271 12597 69280
rect 12556 65717 12596 69271
rect 12652 67649 12692 70951
rect 12747 69152 12789 69161
rect 12747 69112 12748 69152
rect 12788 69112 12789 69152
rect 12747 69103 12789 69112
rect 12748 68489 12788 69103
rect 12747 68480 12789 68489
rect 12747 68440 12748 68480
rect 12788 68440 12789 68480
rect 12747 68431 12789 68440
rect 12748 67817 12788 68431
rect 12747 67808 12789 67817
rect 12747 67768 12748 67808
rect 12788 67768 12789 67808
rect 12747 67759 12789 67768
rect 12652 67609 12788 67649
rect 12555 65708 12597 65717
rect 12555 65668 12556 65708
rect 12596 65668 12597 65708
rect 12555 65659 12597 65668
rect 12556 65540 12596 65549
rect 12596 65500 12692 65540
rect 12556 65491 12596 65500
rect 12652 65297 12692 65500
rect 12651 65288 12693 65297
rect 12651 65248 12652 65288
rect 12692 65248 12693 65288
rect 12651 65239 12693 65248
rect 12556 64028 12596 64037
rect 12651 64028 12693 64037
rect 12596 63988 12652 64028
rect 12692 63988 12693 64028
rect 12556 63979 12596 63988
rect 12651 63979 12693 63988
rect 12748 63281 12788 67609
rect 12747 63272 12789 63281
rect 12747 63232 12748 63272
rect 12788 63232 12789 63272
rect 12747 63223 12789 63232
rect 12748 63113 12788 63223
rect 12747 63104 12789 63113
rect 12747 63064 12748 63104
rect 12788 63064 12789 63104
rect 12747 63055 12789 63064
rect 12460 61720 12596 61760
rect 12460 61592 12500 61603
rect 12460 61517 12500 61552
rect 12459 61508 12501 61517
rect 12459 61468 12460 61508
rect 12500 61468 12501 61508
rect 12459 61459 12501 61468
rect 12459 61172 12501 61181
rect 12459 61132 12460 61172
rect 12500 61132 12501 61172
rect 12459 61123 12501 61132
rect 12460 61088 12500 61123
rect 12460 61037 12500 61048
rect 12316 60910 12404 60920
rect 12356 60880 12404 60910
rect 12316 60861 12356 60870
rect 12076 60796 12212 60836
rect 12076 60089 12116 60796
rect 12171 60668 12213 60677
rect 12556 60668 12596 61720
rect 12171 60628 12172 60668
rect 12212 60628 12213 60668
rect 12171 60619 12213 60628
rect 12268 60628 12596 60668
rect 12075 60080 12117 60089
rect 12075 60040 12076 60080
rect 12116 60040 12117 60080
rect 12075 60031 12117 60040
rect 12172 58652 12212 60619
rect 12172 58603 12212 58612
rect 12268 58652 12308 60628
rect 12459 60500 12501 60509
rect 12459 60460 12460 60500
rect 12500 60460 12501 60500
rect 12459 60451 12501 60460
rect 12460 59324 12500 60451
rect 12651 60416 12693 60425
rect 12651 60376 12652 60416
rect 12692 60376 12693 60416
rect 12651 60367 12693 60376
rect 12460 59284 12596 59324
rect 12171 57980 12213 57989
rect 12171 57940 12172 57980
rect 12212 57940 12213 57980
rect 12171 57931 12213 57940
rect 11979 57056 12021 57065
rect 11979 57016 11980 57056
rect 12020 57016 12021 57056
rect 11979 57007 12021 57016
rect 11980 56922 12020 57007
rect 11980 56384 12020 56393
rect 11884 56344 11980 56384
rect 11980 56335 12020 56344
rect 12075 55628 12117 55637
rect 12075 55588 12076 55628
rect 12116 55588 12117 55628
rect 12075 55579 12117 55588
rect 11932 55553 11972 55562
rect 11972 55513 12020 55544
rect 11932 55504 12020 55513
rect 11404 55420 11732 55460
rect 11403 54872 11445 54881
rect 11403 54832 11404 54872
rect 11444 54832 11445 54872
rect 11403 54823 11445 54832
rect 10924 53311 10964 53320
rect 11020 53488 11156 53528
rect 11212 53488 11348 53528
rect 10828 53226 10868 53311
rect 10827 53108 10869 53117
rect 10827 53068 10828 53108
rect 10868 53068 10869 53108
rect 10827 53059 10869 53068
rect 10731 52940 10773 52949
rect 10731 52900 10732 52940
rect 10772 52900 10773 52940
rect 10731 52891 10773 52900
rect 10155 52436 10197 52445
rect 10155 52396 10156 52436
rect 10196 52396 10197 52436
rect 10155 52387 10197 52396
rect 10252 52361 10292 52480
rect 10540 52480 10676 52520
rect 10731 52520 10773 52529
rect 10731 52480 10732 52520
rect 10772 52480 10773 52520
rect 10251 52352 10293 52361
rect 10251 52312 10252 52352
rect 10292 52312 10293 52352
rect 10251 52303 10293 52312
rect 10444 52352 10484 52363
rect 10444 52277 10484 52312
rect 10443 52268 10485 52277
rect 10443 52228 10444 52268
rect 10484 52228 10485 52268
rect 10443 52219 10485 52228
rect 10443 51932 10485 51941
rect 10443 51892 10444 51932
rect 10484 51892 10485 51932
rect 10443 51883 10485 51892
rect 10060 51052 10292 51092
rect 10155 49832 10197 49841
rect 10155 49792 10156 49832
rect 10196 49792 10197 49832
rect 10155 49783 10197 49792
rect 10156 49589 10196 49783
rect 10155 49580 10197 49589
rect 10155 49540 10156 49580
rect 10196 49540 10197 49580
rect 10155 49531 10197 49540
rect 10060 49496 10100 49505
rect 10060 48833 10100 49456
rect 10156 49446 10196 49531
rect 10252 49328 10292 51052
rect 10156 49288 10292 49328
rect 10059 48824 10101 48833
rect 10059 48784 10060 48824
rect 10100 48784 10101 48824
rect 10059 48775 10101 48784
rect 10156 48572 10196 49288
rect 10251 48824 10293 48833
rect 10251 48784 10252 48824
rect 10292 48784 10293 48824
rect 10251 48775 10293 48784
rect 10348 48824 10388 48833
rect 10444 48824 10484 51883
rect 10388 48784 10484 48824
rect 10348 48775 10388 48784
rect 10252 48690 10292 48775
rect 10156 48532 10484 48572
rect 10251 48236 10293 48245
rect 10251 48196 10252 48236
rect 10292 48196 10293 48236
rect 10251 48187 10293 48196
rect 10252 47993 10292 48187
rect 10251 47984 10293 47993
rect 10251 47944 10252 47984
rect 10292 47944 10293 47984
rect 10251 47935 10293 47944
rect 10252 47850 10292 47935
rect 10060 47816 10100 47825
rect 10100 47776 10196 47816
rect 10060 47767 10100 47776
rect 10156 47307 10196 47776
rect 10348 47396 10388 47405
rect 10156 47258 10196 47267
rect 10252 47356 10348 47396
rect 10252 46901 10292 47356
rect 10348 47347 10388 47356
rect 10347 47144 10389 47153
rect 10347 47104 10348 47144
rect 10388 47104 10389 47144
rect 10347 47095 10389 47104
rect 10251 46892 10293 46901
rect 10251 46852 10252 46892
rect 10292 46852 10293 46892
rect 10251 46843 10293 46852
rect 9772 46516 10004 46556
rect 9676 46472 9716 46481
rect 9579 46052 9621 46061
rect 9579 46012 9580 46052
rect 9620 46012 9621 46052
rect 9579 46003 9621 46012
rect 9676 45893 9716 46432
rect 9675 45884 9717 45893
rect 9675 45844 9676 45884
rect 9716 45844 9717 45884
rect 9675 45835 9717 45844
rect 9579 45800 9621 45809
rect 9579 45760 9580 45800
rect 9620 45760 9621 45800
rect 9579 45751 9621 45760
rect 9388 45676 9524 45716
rect 9387 45548 9429 45557
rect 9387 45508 9388 45548
rect 9428 45508 9429 45548
rect 9387 45499 9429 45508
rect 9388 45414 9428 45499
rect 9291 44960 9333 44969
rect 9291 44920 9292 44960
rect 9332 44920 9333 44960
rect 9291 44911 9333 44920
rect 9292 44826 9332 44911
rect 9196 44239 9236 44248
rect 9100 44154 9140 44239
rect 9003 43784 9045 43793
rect 9003 43744 9004 43784
rect 9044 43744 9045 43784
rect 9003 43735 9045 43744
rect 9099 42692 9141 42701
rect 9099 42652 9100 42692
rect 9140 42652 9141 42692
rect 9099 42643 9141 42652
rect 9100 42104 9140 42643
rect 9140 42064 9236 42104
rect 9100 42055 9140 42064
rect 9004 41180 9044 41189
rect 9004 40433 9044 41140
rect 9100 41180 9140 41189
rect 9100 40517 9140 41140
rect 9099 40508 9141 40517
rect 9099 40468 9100 40508
rect 9140 40468 9141 40508
rect 9099 40459 9141 40468
rect 9003 40424 9045 40433
rect 9003 40384 9004 40424
rect 9044 40384 9045 40424
rect 9003 40375 9045 40384
rect 9100 40256 9140 40265
rect 9196 40256 9236 42064
rect 9484 40592 9524 45676
rect 9580 45666 9620 45751
rect 9772 45548 9812 46516
rect 10156 46472 10196 46481
rect 9868 46388 9908 46397
rect 10156 46388 10196 46432
rect 10252 46472 10292 46483
rect 10252 46397 10292 46432
rect 9908 46348 10196 46388
rect 10251 46388 10293 46397
rect 10251 46348 10252 46388
rect 10292 46348 10293 46388
rect 9868 46339 9908 46348
rect 10251 46339 10293 46348
rect 10059 46220 10101 46229
rect 10059 46180 10060 46220
rect 10100 46180 10101 46220
rect 10059 46171 10101 46180
rect 9867 46052 9909 46061
rect 9867 46012 9868 46052
rect 9908 46012 9909 46052
rect 9867 46003 9909 46012
rect 9580 45508 9812 45548
rect 9580 43952 9620 45508
rect 9868 45389 9908 46003
rect 9867 45380 9909 45389
rect 9867 45340 9868 45380
rect 9908 45340 9909 45380
rect 9867 45331 9909 45340
rect 9963 45212 10005 45221
rect 9963 45172 9964 45212
rect 10004 45172 10005 45212
rect 9963 45163 10005 45172
rect 9867 45128 9909 45137
rect 9867 45088 9868 45128
rect 9908 45088 9909 45128
rect 9867 45079 9909 45088
rect 9771 45044 9813 45053
rect 9771 45004 9772 45044
rect 9812 45004 9813 45044
rect 9771 44995 9813 45004
rect 9868 45044 9908 45079
rect 9675 44960 9717 44969
rect 9675 44920 9676 44960
rect 9716 44920 9717 44960
rect 9675 44911 9717 44920
rect 9676 44288 9716 44911
rect 9772 44910 9812 44995
rect 9868 44993 9908 45004
rect 9676 44239 9716 44248
rect 9580 43912 9716 43952
rect 9579 42860 9621 42869
rect 9579 42820 9580 42860
rect 9620 42820 9621 42860
rect 9579 42811 9621 42820
rect 9580 42726 9620 42811
rect 9676 42608 9716 43912
rect 9964 43700 10004 45163
rect 9868 43660 10004 43700
rect 9771 42860 9813 42869
rect 9771 42820 9772 42860
rect 9812 42820 9813 42860
rect 9771 42811 9813 42820
rect 9580 42568 9716 42608
rect 9580 41264 9620 42568
rect 9676 41936 9716 41947
rect 9772 41945 9812 42811
rect 9676 41861 9716 41896
rect 9771 41936 9813 41945
rect 9771 41896 9772 41936
rect 9812 41896 9813 41936
rect 9771 41887 9813 41896
rect 9675 41852 9717 41861
rect 9675 41812 9676 41852
rect 9716 41812 9717 41852
rect 9675 41803 9717 41812
rect 9772 41802 9812 41887
rect 9580 41215 9620 41224
rect 9484 40552 9620 40592
rect 9387 40340 9429 40349
rect 9387 40300 9388 40340
rect 9428 40300 9429 40340
rect 9387 40291 9429 40300
rect 9140 40216 9236 40256
rect 9100 39920 9140 40216
rect 9100 39871 9140 39880
rect 9388 39752 9428 40291
rect 9388 39703 9428 39712
rect 9484 39752 9524 39761
rect 9580 39752 9620 40552
rect 9868 39920 9908 43660
rect 9963 43532 10005 43541
rect 9963 43492 9964 43532
rect 10004 43492 10005 43532
rect 9963 43483 10005 43492
rect 9964 43448 10004 43483
rect 9964 43397 10004 43408
rect 10060 42701 10100 46171
rect 10348 45128 10388 47095
rect 10444 45212 10484 48532
rect 10540 45296 10580 52480
rect 10731 52471 10773 52480
rect 10828 52520 10868 53059
rect 10923 52688 10965 52697
rect 10923 52648 10924 52688
rect 10964 52648 10965 52688
rect 10923 52639 10965 52648
rect 10924 52529 10964 52639
rect 10828 52471 10868 52480
rect 10923 52520 10965 52529
rect 10923 52480 10924 52520
rect 10964 52480 10965 52520
rect 10923 52471 10965 52480
rect 10732 52386 10772 52471
rect 10635 52352 10677 52361
rect 10635 52312 10636 52352
rect 10676 52312 10677 52352
rect 10635 52303 10677 52312
rect 10923 52352 10965 52361
rect 10923 52312 10924 52352
rect 10964 52312 10965 52352
rect 10923 52303 10965 52312
rect 10636 52218 10676 52303
rect 10635 52100 10677 52109
rect 10635 52060 10636 52100
rect 10676 52060 10677 52100
rect 10635 52051 10677 52060
rect 10636 49496 10676 52051
rect 10676 49456 10868 49496
rect 10636 49447 10676 49456
rect 10635 49328 10677 49337
rect 10635 49288 10636 49328
rect 10676 49288 10677 49328
rect 10635 49279 10677 49288
rect 10636 46472 10676 49279
rect 10828 48824 10868 49456
rect 10828 48775 10868 48784
rect 10924 47825 10964 52303
rect 11020 52277 11060 53488
rect 11115 53360 11157 53369
rect 11115 53320 11116 53360
rect 11156 53320 11157 53360
rect 11115 53311 11157 53320
rect 11116 53226 11156 53311
rect 11115 53108 11157 53117
rect 11115 53068 11116 53108
rect 11156 53068 11157 53108
rect 11115 53059 11157 53068
rect 11116 52974 11156 53059
rect 11115 52856 11157 52865
rect 11115 52816 11116 52856
rect 11156 52816 11157 52856
rect 11115 52807 11157 52816
rect 11116 52520 11156 52807
rect 11212 52688 11252 53488
rect 11308 53360 11348 53371
rect 11308 53285 11348 53320
rect 11307 53276 11349 53285
rect 11307 53236 11308 53276
rect 11348 53236 11349 53276
rect 11307 53227 11349 53236
rect 11404 52772 11444 54823
rect 11500 54041 11540 55420
rect 11980 55040 12020 55504
rect 12076 55460 12116 55579
rect 12076 55411 12116 55420
rect 11980 54991 12020 55000
rect 11787 54956 11829 54965
rect 11787 54916 11788 54956
rect 11828 54916 11829 54956
rect 11787 54907 11829 54916
rect 11788 54872 11828 54907
rect 11499 54032 11541 54041
rect 11499 53992 11500 54032
rect 11540 53992 11541 54032
rect 11499 53983 11541 53992
rect 11595 53864 11637 53873
rect 11595 53824 11596 53864
rect 11636 53824 11637 53864
rect 11595 53815 11637 53824
rect 11499 53696 11541 53705
rect 11499 53656 11500 53696
rect 11540 53656 11541 53696
rect 11499 53647 11541 53656
rect 11404 52723 11444 52732
rect 11212 52648 11348 52688
rect 11212 52520 11252 52529
rect 11116 52480 11212 52520
rect 11212 52471 11252 52480
rect 11115 52352 11157 52361
rect 11115 52312 11116 52352
rect 11156 52312 11157 52352
rect 11115 52303 11157 52312
rect 11019 52268 11061 52277
rect 11019 52228 11020 52268
rect 11060 52228 11061 52268
rect 11019 52219 11061 52228
rect 11116 52218 11156 52303
rect 11308 52016 11348 52648
rect 11500 52016 11540 53647
rect 11596 52520 11636 53815
rect 11691 53360 11733 53369
rect 11691 53320 11692 53360
rect 11732 53320 11733 53360
rect 11691 53311 11733 53320
rect 11692 52604 11732 53311
rect 11788 52697 11828 54832
rect 12075 54032 12117 54041
rect 12075 53992 12076 54032
rect 12116 53992 12117 54032
rect 12075 53983 12117 53992
rect 11979 52940 12021 52949
rect 11979 52900 11980 52940
rect 12020 52900 12021 52940
rect 11979 52891 12021 52900
rect 11787 52688 11829 52697
rect 11787 52648 11788 52688
rect 11828 52648 11924 52688
rect 11787 52639 11829 52648
rect 11692 52555 11732 52564
rect 11596 52471 11636 52480
rect 11787 52520 11829 52529
rect 11787 52480 11788 52520
rect 11828 52480 11829 52520
rect 11787 52471 11829 52480
rect 11788 52386 11828 52471
rect 11884 52109 11924 52648
rect 11883 52100 11925 52109
rect 11883 52060 11884 52100
rect 11924 52060 11925 52100
rect 11883 52051 11925 52060
rect 11020 51976 11348 52016
rect 11404 51976 11540 52016
rect 10731 47816 10773 47825
rect 10731 47776 10732 47816
rect 10772 47776 10773 47816
rect 10731 47767 10773 47776
rect 10923 47816 10965 47825
rect 10923 47776 10924 47816
rect 10964 47776 10965 47816
rect 10923 47767 10965 47776
rect 10732 46556 10772 47767
rect 10923 47396 10965 47405
rect 10923 47356 10924 47396
rect 10964 47356 10965 47396
rect 10923 47347 10965 47356
rect 10827 47312 10869 47321
rect 10827 47272 10828 47312
rect 10868 47272 10869 47312
rect 10827 47263 10869 47272
rect 10924 47312 10964 47347
rect 10828 46901 10868 47263
rect 10924 47237 10964 47272
rect 10923 47228 10965 47237
rect 10923 47188 10924 47228
rect 10964 47188 10965 47228
rect 10923 47179 10965 47188
rect 10924 47148 10964 47179
rect 10827 46892 10869 46901
rect 10827 46852 10828 46892
rect 10868 46852 10869 46892
rect 10827 46843 10869 46852
rect 11020 46640 11060 51976
rect 11116 51848 11156 51857
rect 11404 51848 11444 51976
rect 11156 51808 11444 51848
rect 11499 51848 11541 51857
rect 11499 51808 11500 51848
rect 11540 51808 11541 51848
rect 11116 50261 11156 51808
rect 11499 51799 11541 51808
rect 11500 51714 11540 51799
rect 11308 51596 11348 51605
rect 11212 51556 11308 51596
rect 11212 50588 11252 51556
rect 11308 51547 11348 51556
rect 11320 51017 11360 51036
rect 11308 51008 11360 51017
rect 11348 50968 11444 51008
rect 11308 50959 11348 50968
rect 11212 50548 11348 50588
rect 11211 50336 11253 50345
rect 11211 50296 11212 50336
rect 11252 50296 11253 50336
rect 11211 50287 11253 50296
rect 11115 50252 11157 50261
rect 11115 50212 11116 50252
rect 11156 50212 11157 50252
rect 11115 50203 11157 50212
rect 11212 50202 11252 50287
rect 11308 49580 11348 50548
rect 11404 50513 11444 50968
rect 11403 50504 11445 50513
rect 11403 50464 11404 50504
rect 11444 50464 11445 50504
rect 11403 50455 11445 50464
rect 11787 49664 11829 49673
rect 11787 49624 11788 49664
rect 11828 49624 11829 49664
rect 11787 49615 11829 49624
rect 11308 49540 11444 49580
rect 11116 49501 11156 49510
rect 11116 49169 11156 49461
rect 11307 49412 11349 49421
rect 11307 49372 11308 49412
rect 11348 49372 11349 49412
rect 11307 49363 11349 49372
rect 11308 49278 11348 49363
rect 11115 49160 11157 49169
rect 11404 49160 11444 49540
rect 11115 49120 11116 49160
rect 11156 49120 11157 49160
rect 11115 49111 11157 49120
rect 11356 49120 11444 49160
rect 11595 49160 11637 49169
rect 11595 49120 11596 49160
rect 11636 49120 11637 49160
rect 11356 48814 11396 49120
rect 11595 49111 11637 49120
rect 11499 48908 11541 48917
rect 11499 48868 11500 48908
rect 11540 48868 11541 48908
rect 11499 48859 11541 48868
rect 11500 48774 11540 48859
rect 11356 48765 11396 48774
rect 11499 48320 11541 48329
rect 11499 48280 11500 48320
rect 11540 48280 11541 48320
rect 11499 48271 11541 48280
rect 11500 47984 11540 48271
rect 11596 48236 11636 49111
rect 11692 48824 11732 48833
rect 11692 48581 11732 48784
rect 11691 48572 11733 48581
rect 11691 48532 11692 48572
rect 11732 48532 11733 48572
rect 11691 48523 11733 48532
rect 11692 48236 11732 48245
rect 11596 48196 11692 48236
rect 11692 48187 11732 48196
rect 11403 47900 11445 47909
rect 11500 47900 11540 47944
rect 11403 47860 11404 47900
rect 11444 47860 11540 47900
rect 11403 47851 11445 47860
rect 11788 47816 11828 49615
rect 11883 48488 11925 48497
rect 11883 48448 11884 48488
rect 11924 48448 11925 48488
rect 11883 48439 11925 48448
rect 11500 47776 11828 47816
rect 11020 46600 11156 46640
rect 10732 46507 10772 46516
rect 10636 46388 10676 46432
rect 10923 46388 10965 46397
rect 10636 46348 10772 46388
rect 10540 45256 10676 45296
rect 10444 45172 10580 45212
rect 10348 45088 10484 45128
rect 10252 44960 10292 44969
rect 10252 44801 10292 44920
rect 10348 44960 10388 44969
rect 10251 44792 10293 44801
rect 10251 44752 10252 44792
rect 10292 44752 10293 44792
rect 10251 44743 10293 44752
rect 10252 44297 10292 44743
rect 10348 44549 10388 44920
rect 10347 44540 10389 44549
rect 10347 44500 10348 44540
rect 10388 44500 10389 44540
rect 10347 44491 10389 44500
rect 10348 44372 10388 44381
rect 10251 44288 10293 44297
rect 10156 44274 10196 44283
rect 10251 44248 10252 44288
rect 10292 44248 10293 44288
rect 10251 44239 10293 44248
rect 10156 43700 10196 44234
rect 10156 43651 10196 43660
rect 10059 42692 10101 42701
rect 10059 42652 10060 42692
rect 10100 42652 10101 42692
rect 10059 42643 10101 42652
rect 9963 41936 10005 41945
rect 9963 41896 9964 41936
rect 10004 41896 10005 41936
rect 9963 41887 10005 41896
rect 9524 39712 9620 39752
rect 9676 39880 9908 39920
rect 9964 39920 10004 41887
rect 10060 41861 10100 42643
rect 10251 42272 10293 42281
rect 10251 42232 10252 42272
rect 10292 42232 10293 42272
rect 10251 42223 10293 42232
rect 10252 42020 10292 42223
rect 10252 41971 10292 41980
rect 10155 41936 10197 41945
rect 10155 41896 10156 41936
rect 10196 41896 10197 41936
rect 10155 41887 10197 41896
rect 10059 41852 10101 41861
rect 10059 41812 10060 41852
rect 10100 41812 10101 41852
rect 10059 41803 10101 41812
rect 10156 41802 10196 41887
rect 10348 41516 10388 44332
rect 10156 41476 10388 41516
rect 10059 41348 10101 41357
rect 10059 41308 10060 41348
rect 10100 41308 10101 41348
rect 10059 41299 10101 41308
rect 10060 41259 10100 41299
rect 10060 41210 10100 41219
rect 9964 39880 10100 39920
rect 9004 39584 9044 39593
rect 9004 38912 9044 39544
rect 9099 39584 9141 39593
rect 9099 39544 9100 39584
rect 9140 39544 9141 39584
rect 9099 39535 9141 39544
rect 9004 38408 9044 38872
rect 8907 38240 8949 38249
rect 8907 38200 8908 38240
rect 8948 38200 8949 38240
rect 8907 38191 8949 38200
rect 8811 37652 8853 37661
rect 8811 37612 8812 37652
rect 8852 37612 8853 37652
rect 8811 37603 8853 37612
rect 8812 37518 8852 37603
rect 8620 36728 8660 37360
rect 8331 36560 8373 36569
rect 8331 36520 8332 36560
rect 8372 36520 8373 36560
rect 8331 36511 8373 36520
rect 8620 35981 8660 36688
rect 9004 37232 9044 38368
rect 8811 36560 8853 36569
rect 8811 36520 8812 36560
rect 8852 36520 8853 36560
rect 8811 36511 8853 36520
rect 9004 36560 9044 37192
rect 8812 36426 8852 36511
rect 8811 36056 8853 36065
rect 8811 36016 8812 36056
rect 8852 36016 8853 36056
rect 8811 36007 8853 36016
rect 8619 35972 8661 35981
rect 8619 35932 8620 35972
rect 8660 35932 8661 35972
rect 8619 35923 8661 35932
rect 8620 35888 8660 35923
rect 8812 35922 8852 36007
rect 8620 35837 8660 35848
rect 9004 35720 9044 36520
rect 8235 35300 8277 35309
rect 8235 35260 8236 35300
rect 8276 35260 8277 35300
rect 8235 35251 8277 35260
rect 8619 35300 8661 35309
rect 8619 35260 8620 35300
rect 8660 35260 8661 35300
rect 8619 35251 8661 35260
rect 7851 35216 7893 35225
rect 7851 35176 7852 35216
rect 7892 35176 7893 35216
rect 7851 35167 7893 35176
rect 8140 35216 8180 35225
rect 7852 35082 7892 35167
rect 8140 35048 8180 35176
rect 8236 35166 8276 35251
rect 8235 35048 8277 35057
rect 8140 35008 8236 35048
rect 8276 35008 8277 35048
rect 8235 34999 8277 35008
rect 7851 34964 7893 34973
rect 7851 34924 7852 34964
rect 7892 34924 7893 34964
rect 7851 34915 7893 34924
rect 7755 34376 7797 34385
rect 7755 34336 7756 34376
rect 7796 34336 7797 34376
rect 7755 34327 7797 34336
rect 7659 34292 7701 34301
rect 7659 34252 7660 34292
rect 7700 34252 7701 34292
rect 7659 34243 7701 34252
rect 7756 34242 7796 34327
rect 7276 34000 7508 34040
rect 7564 34208 7604 34217
rect 7179 33368 7221 33377
rect 7179 33328 7180 33368
rect 7220 33328 7221 33368
rect 7179 33319 7221 33328
rect 7179 32780 7221 32789
rect 7179 32740 7180 32780
rect 7220 32740 7221 32780
rect 7179 32731 7221 32740
rect 7180 32646 7220 32731
rect 7083 32360 7125 32369
rect 7083 32320 7084 32360
rect 7124 32320 7125 32360
rect 7083 32311 7125 32320
rect 6987 32108 7029 32117
rect 6987 32068 6988 32108
rect 7028 32068 7029 32108
rect 6987 32059 7029 32068
rect 6988 31613 7028 32059
rect 7276 31940 7316 34000
rect 7564 33956 7604 34168
rect 7755 34124 7797 34133
rect 7755 34084 7756 34124
rect 7796 34084 7797 34124
rect 7755 34075 7797 34084
rect 7468 33916 7604 33956
rect 7468 33704 7508 33916
rect 7659 33872 7701 33881
rect 7659 33832 7660 33872
rect 7700 33832 7701 33872
rect 7659 33823 7701 33832
rect 7563 33788 7605 33797
rect 7563 33748 7564 33788
rect 7604 33748 7605 33788
rect 7563 33739 7605 33748
rect 7420 33694 7508 33704
rect 7460 33664 7508 33694
rect 7564 33654 7604 33739
rect 7420 33645 7460 33654
rect 7468 32864 7508 32875
rect 7468 32789 7508 32824
rect 7564 32864 7604 32873
rect 7467 32780 7509 32789
rect 7467 32740 7468 32780
rect 7508 32740 7509 32780
rect 7467 32731 7509 32740
rect 7276 31900 7508 31940
rect 6987 31604 7029 31613
rect 6987 31564 6988 31604
rect 7028 31564 7029 31604
rect 6987 31555 7029 31564
rect 7275 31520 7317 31529
rect 7275 31480 7276 31520
rect 7316 31480 7317 31520
rect 7275 31471 7317 31480
rect 6891 31352 6933 31361
rect 6891 31312 6892 31352
rect 6932 31312 6933 31352
rect 6891 31303 6933 31312
rect 7276 31352 7316 31471
rect 7316 31312 7412 31352
rect 7276 31303 7316 31312
rect 6892 31218 6932 31303
rect 7083 31184 7125 31193
rect 7083 31144 7084 31184
rect 7124 31144 7125 31184
rect 7083 31135 7125 31144
rect 7084 31050 7124 31135
rect 6796 30892 6932 30932
rect 6796 30764 6836 30773
rect 6508 30724 6796 30764
rect 6411 30428 6453 30437
rect 6411 30388 6412 30428
rect 6452 30388 6453 30428
rect 6411 30379 6453 30388
rect 6411 30092 6453 30101
rect 6411 30052 6412 30092
rect 6452 30052 6453 30092
rect 6411 30043 6453 30052
rect 6412 29958 6452 30043
rect 6508 29840 6548 30724
rect 6796 30715 6836 30724
rect 6604 30666 6644 30675
rect 6604 29849 6644 30626
rect 6699 30344 6741 30353
rect 6699 30304 6700 30344
rect 6740 30304 6741 30344
rect 6699 30295 6741 30304
rect 6316 29800 6452 29840
rect 6028 29632 6164 29672
rect 6219 29672 6261 29681
rect 6219 29632 6220 29672
rect 6260 29632 6261 29672
rect 5931 29420 5973 29429
rect 5931 29380 5932 29420
rect 5972 29380 5973 29420
rect 5931 29371 5973 29380
rect 5739 28244 5781 28253
rect 5739 28204 5740 28244
rect 5780 28204 5781 28244
rect 5739 28195 5781 28204
rect 5644 27952 5780 27992
rect 5740 27833 5780 27952
rect 5739 27824 5781 27833
rect 5452 27784 5588 27824
rect 4587 27775 4629 27784
rect 4972 27656 5012 27665
rect 5452 27656 5492 27665
rect 4684 27616 4972 27642
rect 4684 27602 5012 27616
rect 5068 27616 5452 27656
rect 4587 26816 4629 26825
rect 4492 26776 4588 26816
rect 4628 26776 4629 26816
rect 4587 26767 4629 26776
rect 4491 25304 4533 25313
rect 4491 25264 4492 25304
rect 4532 25264 4533 25304
rect 4491 25255 4533 25264
rect 4395 25220 4437 25229
rect 4395 25180 4396 25220
rect 4436 25180 4437 25220
rect 4395 25171 4437 25180
rect 4396 24632 4436 25171
rect 4492 25170 4532 25255
rect 4396 24389 4436 24592
rect 4395 24380 4437 24389
rect 4395 24340 4396 24380
rect 4436 24340 4437 24380
rect 4395 24331 4437 24340
rect 4588 24212 4628 26767
rect 4300 24172 4436 24212
rect 4052 23248 4148 23288
rect 4300 23792 4340 23801
rect 4012 23239 4052 23248
rect 3340 23120 3380 23129
rect 3340 22373 3380 23080
rect 3436 23120 3476 23239
rect 3627 23204 3669 23213
rect 3627 23164 3628 23204
rect 3668 23164 3669 23204
rect 3627 23155 3669 23164
rect 4203 23204 4245 23213
rect 4203 23164 4204 23204
rect 4244 23164 4245 23204
rect 4203 23155 4245 23164
rect 3436 23071 3476 23080
rect 3532 23120 3572 23129
rect 3532 22448 3572 23080
rect 3628 23070 3668 23155
rect 3819 23120 3861 23129
rect 3819 23080 3820 23120
rect 3860 23080 3861 23120
rect 3819 23071 3861 23080
rect 4108 23120 4148 23129
rect 3820 22986 3860 23071
rect 4108 22961 4148 23080
rect 4107 22952 4149 22961
rect 4107 22912 4108 22952
rect 4148 22912 4149 22952
rect 4107 22903 4149 22912
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 4011 22532 4053 22541
rect 4011 22492 4012 22532
rect 4052 22492 4053 22532
rect 4011 22483 4053 22492
rect 3436 22408 3572 22448
rect 3915 22448 3957 22457
rect 3915 22408 3916 22448
rect 3956 22408 3957 22448
rect 3339 22364 3381 22373
rect 3339 22324 3340 22364
rect 3380 22324 3381 22364
rect 3339 22315 3381 22324
rect 3340 21617 3380 22315
rect 3436 21776 3476 22408
rect 3915 22399 3957 22408
rect 3532 22280 3572 22291
rect 3532 22205 3572 22240
rect 3627 22280 3669 22289
rect 3627 22240 3628 22280
rect 3668 22240 3669 22280
rect 3627 22231 3669 22240
rect 3819 22280 3861 22289
rect 3819 22240 3820 22280
rect 3860 22240 3861 22280
rect 3819 22231 3861 22240
rect 3531 22196 3573 22205
rect 3531 22156 3532 22196
rect 3572 22156 3573 22196
rect 3531 22147 3573 22156
rect 3628 22146 3668 22231
rect 3436 21727 3476 21736
rect 3531 21692 3573 21701
rect 3531 21652 3532 21692
rect 3572 21652 3573 21692
rect 3531 21643 3573 21652
rect 3723 21692 3765 21701
rect 3723 21652 3724 21692
rect 3764 21652 3765 21692
rect 3723 21643 3765 21652
rect 3339 21608 3381 21617
rect 3339 21568 3340 21608
rect 3380 21568 3381 21608
rect 3532 21598 3572 21643
rect 3339 21559 3381 21568
rect 3436 21558 3572 21598
rect 3627 21608 3669 21617
rect 3627 21568 3628 21608
rect 3668 21568 3669 21608
rect 3627 21559 3669 21568
rect 3724 21608 3764 21643
rect 3436 20852 3476 21558
rect 3628 21474 3668 21559
rect 3724 21557 3764 21568
rect 3820 21440 3860 22231
rect 3916 21776 3956 22399
rect 3916 21727 3956 21736
rect 4012 21608 4052 22483
rect 4107 22280 4149 22289
rect 4107 22240 4108 22280
rect 4148 22240 4149 22280
rect 4107 22231 4149 22240
rect 4108 22146 4148 22231
rect 4204 22028 4244 23155
rect 4300 22625 4340 23752
rect 4299 22616 4341 22625
rect 4299 22576 4300 22616
rect 4340 22576 4341 22616
rect 4299 22567 4341 22576
rect 4396 22037 4436 24172
rect 4492 24172 4628 24212
rect 4492 23549 4532 24172
rect 4588 23969 4628 24054
rect 4587 23960 4629 23969
rect 4587 23920 4588 23960
rect 4628 23920 4629 23960
rect 4587 23911 4629 23920
rect 4588 23792 4628 23801
rect 4588 23633 4628 23752
rect 4587 23624 4629 23633
rect 4587 23584 4588 23624
rect 4628 23584 4629 23624
rect 4587 23575 4629 23584
rect 4491 23540 4533 23549
rect 4491 23500 4492 23540
rect 4532 23500 4533 23540
rect 4491 23491 4533 23500
rect 4587 23456 4629 23465
rect 4587 23416 4588 23456
rect 4628 23416 4629 23456
rect 4587 23407 4629 23416
rect 4491 23204 4533 23213
rect 4491 23164 4492 23204
rect 4532 23164 4533 23204
rect 4491 23155 4533 23164
rect 4492 23120 4532 23155
rect 4492 23069 4532 23080
rect 4588 22952 4628 23407
rect 4492 22912 4628 22952
rect 4012 21559 4052 21568
rect 4108 21988 4244 22028
rect 4395 22028 4437 22037
rect 4395 21988 4396 22028
rect 4436 21988 4437 22028
rect 4108 21608 4148 21988
rect 4395 21979 4437 21988
rect 4203 21776 4245 21785
rect 4203 21736 4204 21776
rect 4244 21736 4245 21776
rect 4203 21727 4245 21736
rect 4108 21559 4148 21568
rect 4204 21608 4244 21727
rect 4204 21559 4244 21568
rect 4396 21608 4436 21619
rect 4396 21533 4436 21568
rect 4492 21608 4532 22912
rect 4588 22373 4628 22389
rect 4587 22364 4629 22373
rect 4587 22324 4588 22364
rect 4628 22324 4629 22364
rect 4587 22315 4629 22324
rect 4588 22294 4628 22315
rect 4588 22245 4628 22254
rect 4684 21944 4724 27602
rect 5068 27068 5108 27616
rect 5452 27607 5492 27616
rect 5163 27488 5205 27497
rect 5163 27448 5164 27488
rect 5204 27448 5205 27488
rect 5163 27439 5205 27448
rect 5355 27488 5397 27497
rect 5355 27448 5356 27488
rect 5396 27448 5397 27488
rect 5355 27439 5397 27448
rect 5164 27354 5204 27439
rect 5068 27019 5108 27028
rect 4876 26825 4916 26910
rect 4875 26816 4917 26825
rect 4875 26776 4876 26816
rect 4916 26776 4917 26816
rect 4875 26767 4917 26776
rect 5356 26816 5396 27439
rect 5356 26767 5396 26776
rect 5068 26648 5108 26657
rect 4780 26608 5068 26648
rect 4780 25565 4820 26608
rect 5068 26599 5108 26608
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 5067 26312 5109 26321
rect 5067 26272 5068 26312
rect 5108 26272 5109 26312
rect 5067 26263 5109 26272
rect 5068 26144 5108 26263
rect 5452 26144 5492 26153
rect 5548 26144 5588 27784
rect 5739 27784 5740 27824
rect 5780 27784 5781 27824
rect 5739 27775 5781 27784
rect 5740 27656 5780 27665
rect 5740 27245 5780 27616
rect 5836 27656 5876 27665
rect 5739 27236 5781 27245
rect 5739 27196 5740 27236
rect 5780 27196 5781 27236
rect 5739 27187 5781 27196
rect 5644 27077 5684 27162
rect 5643 27068 5685 27077
rect 5643 27028 5644 27068
rect 5684 27028 5685 27068
rect 5643 27019 5685 27028
rect 5068 26095 5108 26104
rect 5356 26104 5452 26144
rect 5492 26104 5588 26144
rect 5644 26816 5684 26825
rect 4779 25556 4821 25565
rect 4779 25516 4780 25556
rect 4820 25516 4821 25556
rect 4779 25507 4821 25516
rect 4780 23792 4820 25507
rect 4972 25304 5012 25313
rect 4972 25145 5012 25264
rect 5068 25304 5108 25315
rect 5068 25229 5108 25264
rect 5356 25229 5396 26104
rect 5452 26095 5492 26104
rect 5547 25388 5589 25397
rect 5547 25348 5548 25388
rect 5588 25348 5589 25388
rect 5547 25339 5589 25348
rect 5452 25304 5492 25313
rect 5067 25220 5109 25229
rect 5067 25180 5068 25220
rect 5108 25180 5109 25220
rect 5067 25171 5109 25180
rect 5355 25220 5397 25229
rect 5355 25180 5356 25220
rect 5396 25180 5397 25220
rect 5355 25171 5397 25180
rect 4971 25136 5013 25145
rect 4971 25096 4972 25136
rect 5012 25096 5013 25136
rect 4971 25087 5013 25096
rect 5452 24977 5492 25264
rect 5548 25304 5588 25339
rect 5548 25253 5588 25264
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 5451 24968 5493 24977
rect 5451 24928 5452 24968
rect 5492 24928 5493 24968
rect 5451 24919 5493 24928
rect 5355 24632 5397 24641
rect 5355 24592 5356 24632
rect 5396 24592 5397 24632
rect 5355 24583 5397 24592
rect 5452 24632 5492 24641
rect 5492 24592 5588 24632
rect 5452 24583 5492 24592
rect 4875 24548 4917 24557
rect 4875 24508 4876 24548
rect 4916 24508 4917 24548
rect 4875 24499 4917 24508
rect 4972 24548 5012 24557
rect 4876 24414 4916 24499
rect 4972 24305 5012 24508
rect 5356 24498 5396 24583
rect 4971 24296 5013 24305
rect 4971 24256 4972 24296
rect 5012 24256 5013 24296
rect 4971 24247 5013 24256
rect 4780 23743 4820 23752
rect 4876 23792 4916 23801
rect 4876 23624 4916 23752
rect 5068 23792 5108 23801
rect 5068 23633 5108 23752
rect 5164 23792 5204 23801
rect 5204 23752 5492 23792
rect 5164 23743 5204 23752
rect 4780 23584 4916 23624
rect 5067 23624 5109 23633
rect 5067 23584 5068 23624
rect 5108 23584 5109 23624
rect 4780 22877 4820 23584
rect 5067 23575 5109 23584
rect 5356 23624 5396 23633
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 4779 22868 4821 22877
rect 4779 22828 4780 22868
rect 4820 22828 4821 22868
rect 4779 22819 4821 22828
rect 4779 22700 4821 22709
rect 4779 22660 4780 22700
rect 4820 22660 4821 22700
rect 4779 22651 4821 22660
rect 4780 22196 4820 22651
rect 5356 22541 5396 23584
rect 5452 22709 5492 23752
rect 5548 23129 5588 24592
rect 5644 23969 5684 26776
rect 5836 26657 5876 27616
rect 5932 27329 5972 29371
rect 5931 27320 5973 27329
rect 5931 27280 5932 27320
rect 5972 27280 5973 27320
rect 5931 27271 5973 27280
rect 6028 26825 6068 29632
rect 6219 29623 6261 29632
rect 6124 27404 6164 27413
rect 6027 26816 6069 26825
rect 6027 26776 6028 26816
rect 6068 26776 6069 26816
rect 6027 26767 6069 26776
rect 6028 26682 6068 26767
rect 5835 26648 5877 26657
rect 5835 26608 5836 26648
rect 5876 26608 5877 26648
rect 5835 26599 5877 26608
rect 6124 26312 6164 27364
rect 5932 26272 6164 26312
rect 5835 25388 5877 25397
rect 5835 25348 5836 25388
rect 5876 25348 5877 25388
rect 5835 25339 5877 25348
rect 5836 25304 5876 25339
rect 5836 25253 5876 25264
rect 5932 25304 5972 26272
rect 6027 25724 6069 25733
rect 6027 25684 6028 25724
rect 6068 25684 6069 25724
rect 6027 25675 6069 25684
rect 5932 25255 5972 25264
rect 6028 25220 6068 25675
rect 6028 25180 6164 25220
rect 6124 25136 6164 25180
rect 6124 25087 6164 25096
rect 5739 24884 5781 24893
rect 5739 24844 5740 24884
rect 5780 24844 5781 24884
rect 5739 24835 5781 24844
rect 5643 23960 5685 23969
rect 5643 23920 5644 23960
rect 5684 23920 5685 23960
rect 5643 23911 5685 23920
rect 5547 23120 5589 23129
rect 5740 23120 5780 24835
rect 6123 24716 6165 24725
rect 6123 24676 6124 24716
rect 6164 24676 6165 24716
rect 6123 24667 6165 24676
rect 6124 24632 6164 24667
rect 6124 24581 6164 24592
rect 5835 24380 5877 24389
rect 5835 24340 5836 24380
rect 5876 24340 5877 24380
rect 5835 24331 5877 24340
rect 6123 24380 6165 24389
rect 6123 24340 6124 24380
rect 6164 24340 6165 24380
rect 6123 24331 6165 24340
rect 5547 23080 5548 23120
rect 5588 23080 5589 23120
rect 5547 23071 5589 23080
rect 5644 23080 5740 23120
rect 5644 22709 5684 23080
rect 5740 23071 5780 23080
rect 5836 22952 5876 24331
rect 6028 23801 6068 23886
rect 6027 23792 6069 23801
rect 6027 23752 6028 23792
rect 6068 23752 6069 23792
rect 6027 23743 6069 23752
rect 5931 23204 5973 23213
rect 5931 23164 5932 23204
rect 5972 23164 5973 23204
rect 5931 23155 5973 23164
rect 5932 23070 5972 23155
rect 5740 22912 5876 22952
rect 5451 22700 5493 22709
rect 5451 22660 5452 22700
rect 5492 22660 5493 22700
rect 5451 22651 5493 22660
rect 5643 22700 5685 22709
rect 5643 22660 5644 22700
rect 5684 22660 5685 22700
rect 5643 22651 5685 22660
rect 5355 22532 5397 22541
rect 5355 22492 5356 22532
rect 5396 22492 5397 22532
rect 5355 22483 5397 22492
rect 5452 22457 5492 22542
rect 5451 22448 5493 22457
rect 5451 22408 5452 22448
rect 5492 22408 5493 22448
rect 5451 22399 5493 22408
rect 4780 22147 4820 22156
rect 5260 22280 5300 22289
rect 5260 22121 5300 22240
rect 5452 22280 5492 22289
rect 5452 22196 5492 22240
rect 5644 22196 5684 22205
rect 5452 22156 5644 22196
rect 5644 22147 5684 22156
rect 5259 22112 5301 22121
rect 5259 22072 5260 22112
rect 5300 22072 5301 22112
rect 5259 22063 5301 22072
rect 4395 21524 4437 21533
rect 4395 21484 4396 21524
rect 4436 21484 4437 21524
rect 4395 21475 4437 21484
rect 3724 21400 3860 21440
rect 3724 21356 3764 21400
rect 4492 21356 4532 21568
rect 3436 20803 3476 20812
rect 3532 21316 3764 21356
rect 4300 21316 4532 21356
rect 4588 21904 4724 21944
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 3532 20852 3572 21316
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 3532 20803 3572 20812
rect 4012 20768 4052 20777
rect 4012 19853 4052 20728
rect 4107 20432 4149 20441
rect 4107 20392 4108 20432
rect 4148 20392 4149 20432
rect 4107 20383 4149 20392
rect 4108 20096 4148 20383
rect 4300 20273 4340 21316
rect 4588 20936 4628 21904
rect 4928 21895 5296 21904
rect 4683 21776 4725 21785
rect 4683 21736 4684 21776
rect 4724 21736 4725 21776
rect 4683 21727 4725 21736
rect 4684 21642 4724 21727
rect 5355 21692 5397 21701
rect 5355 21652 5356 21692
rect 5396 21652 5397 21692
rect 5355 21643 5397 21652
rect 4396 20896 4628 20936
rect 4299 20264 4341 20273
rect 4299 20224 4300 20264
rect 4340 20224 4341 20264
rect 4299 20215 4341 20224
rect 3531 19844 3573 19853
rect 3531 19804 3532 19844
rect 3572 19804 3573 19844
rect 3531 19795 3573 19804
rect 4011 19844 4053 19853
rect 4011 19804 4012 19844
rect 4052 19804 4053 19844
rect 4011 19795 4053 19804
rect 3339 18584 3381 18593
rect 3339 18544 3340 18584
rect 3380 18544 3381 18584
rect 3339 18535 3381 18544
rect 3340 18450 3380 18535
rect 3435 18080 3477 18089
rect 3435 18040 3436 18080
rect 3476 18040 3477 18080
rect 3435 18031 3477 18040
rect 3339 17996 3381 18005
rect 3244 17956 3340 17996
rect 3380 17956 3381 17996
rect 2859 17912 2901 17921
rect 2859 17872 2860 17912
rect 2900 17872 2901 17912
rect 2859 17863 2901 17872
rect 2763 17828 2805 17837
rect 2763 17788 2764 17828
rect 2804 17788 2805 17828
rect 2763 17779 2805 17788
rect 2860 17828 2900 17863
rect 2572 17452 2708 17492
rect 2380 17368 2612 17408
rect 2475 17072 2517 17081
rect 2475 17032 2476 17072
rect 2516 17032 2517 17072
rect 2475 17023 2517 17032
rect 2476 16938 2516 17023
rect 2284 16360 2420 16400
rect 2283 16232 2325 16241
rect 2283 16192 2284 16232
rect 2324 16192 2325 16232
rect 2283 16183 2325 16192
rect 2284 16098 2324 16183
rect 2188 14344 2324 14384
rect 2187 14216 2229 14225
rect 2187 14176 2188 14216
rect 2228 14176 2229 14216
rect 2187 14167 2229 14176
rect 2091 11276 2133 11285
rect 2091 11236 2092 11276
rect 2132 11236 2133 11276
rect 2091 11227 2133 11236
rect 1995 10940 2037 10949
rect 1995 10900 1996 10940
rect 2036 10900 2037 10940
rect 1995 10891 2037 10900
rect 1900 10732 2036 10772
rect 1268 10144 1652 10184
rect 1228 10135 1268 10144
rect 1803 9764 1845 9773
rect 1803 9724 1804 9764
rect 1844 9724 1845 9764
rect 1803 9715 1845 9724
rect 1611 9512 1653 9521
rect 1611 9472 1612 9512
rect 1652 9472 1653 9512
rect 1611 9463 1653 9472
rect 1612 9378 1652 9463
rect 363 8672 405 8681
rect 363 8632 364 8672
rect 404 8632 405 8672
rect 363 8623 405 8632
rect 1804 80 1844 9715
rect 1899 9428 1941 9437
rect 1899 9388 1900 9428
rect 1940 9388 1941 9428
rect 1899 9379 1941 9388
rect 1900 8672 1940 9379
rect 1900 8623 1940 8632
rect 1996 80 2036 10732
rect 2188 80 2228 14167
rect 2284 6320 2324 14344
rect 2380 8261 2420 16360
rect 2475 15140 2517 15149
rect 2475 15100 2476 15140
rect 2516 15100 2517 15140
rect 2475 15091 2517 15100
rect 2476 14720 2516 15091
rect 2572 14972 2612 17368
rect 2668 17249 2708 17452
rect 2667 17240 2709 17249
rect 2667 17200 2668 17240
rect 2708 17200 2709 17240
rect 2667 17191 2709 17200
rect 2667 17072 2709 17081
rect 2667 17032 2668 17072
rect 2708 17032 2709 17072
rect 2667 17023 2709 17032
rect 2668 16904 2708 17023
rect 2668 16855 2708 16864
rect 2764 16241 2804 17779
rect 2860 17777 2900 17788
rect 2955 17828 2997 17837
rect 2955 17788 2956 17828
rect 2996 17788 2997 17828
rect 2955 17779 2997 17788
rect 2956 17694 2996 17779
rect 3052 17744 3092 17956
rect 3339 17947 3381 17956
rect 3436 17744 3476 18031
rect 3052 17704 3188 17744
rect 3051 17576 3093 17585
rect 3051 17536 3052 17576
rect 3092 17536 3093 17576
rect 3051 17527 3093 17536
rect 2955 17408 2997 17417
rect 2955 17368 2956 17408
rect 2996 17368 2997 17408
rect 2955 17359 2997 17368
rect 2956 17072 2996 17359
rect 2956 17023 2996 17032
rect 2859 16904 2901 16913
rect 2859 16864 2860 16904
rect 2900 16864 2901 16904
rect 2859 16855 2901 16864
rect 2860 16770 2900 16855
rect 2763 16232 2805 16241
rect 2763 16192 2764 16232
rect 2804 16192 2805 16232
rect 2763 16183 2805 16192
rect 2859 15812 2901 15821
rect 2859 15772 2860 15812
rect 2900 15772 2901 15812
rect 2859 15763 2901 15772
rect 2860 15560 2900 15763
rect 3052 15728 3092 17527
rect 3052 15679 3092 15688
rect 2860 15149 2900 15520
rect 2859 15140 2901 15149
rect 2859 15100 2860 15140
rect 2900 15100 2901 15140
rect 2859 15091 2901 15100
rect 2668 14972 2708 14981
rect 2572 14932 2668 14972
rect 2668 14923 2708 14932
rect 3148 14888 3188 17704
rect 3436 17695 3476 17704
rect 3435 17576 3477 17585
rect 3435 17536 3436 17576
rect 3476 17536 3477 17576
rect 3435 17527 3477 17536
rect 3238 17156 3280 17165
rect 3238 17116 3239 17156
rect 3279 17116 3280 17156
rect 3238 17107 3280 17116
rect 3239 17072 3279 17107
rect 3239 17021 3279 17032
rect 3340 17072 3380 17081
rect 3340 16988 3380 17032
rect 3436 17072 3476 17527
rect 3532 17240 3572 19795
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 4108 18677 4148 20056
rect 4299 19928 4341 19937
rect 4299 19888 4300 19928
rect 4340 19888 4341 19928
rect 4299 19879 4341 19888
rect 4300 19794 4340 19879
rect 4396 19676 4436 20896
rect 4492 20773 4532 20782
rect 4492 19937 4532 20733
rect 4683 20684 4725 20693
rect 4683 20644 4684 20684
rect 4724 20644 4725 20684
rect 4683 20635 4725 20644
rect 4684 20550 4724 20635
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 4928 20383 5296 20392
rect 5356 20264 5396 21643
rect 5451 21608 5493 21617
rect 5451 21568 5452 21608
rect 5492 21568 5493 21608
rect 5451 21559 5493 21568
rect 5452 21474 5492 21559
rect 5547 21440 5589 21449
rect 5547 21400 5548 21440
rect 5588 21400 5589 21440
rect 5547 21391 5589 21400
rect 5452 20768 5492 20777
rect 5452 20609 5492 20728
rect 5451 20600 5493 20609
rect 5451 20560 5452 20600
rect 5492 20560 5493 20600
rect 5451 20551 5493 20560
rect 5451 20348 5493 20357
rect 5451 20308 5452 20348
rect 5492 20308 5493 20348
rect 5451 20299 5493 20308
rect 5164 20224 5396 20264
rect 4683 20180 4725 20189
rect 4683 20140 4684 20180
rect 4724 20140 4725 20180
rect 4683 20131 4725 20140
rect 4588 20096 4628 20105
rect 4491 19928 4533 19937
rect 4491 19888 4492 19928
rect 4532 19888 4533 19928
rect 4491 19879 4533 19888
rect 4300 19636 4436 19676
rect 4300 19349 4340 19636
rect 4492 19508 4532 19517
rect 4588 19508 4628 20056
rect 4684 20096 4724 20131
rect 4684 20045 4724 20056
rect 5164 20096 5204 20224
rect 5164 20047 5204 20056
rect 5068 20012 5108 20023
rect 5068 19937 5108 19972
rect 5067 19928 5109 19937
rect 5067 19888 5068 19928
rect 5108 19888 5109 19928
rect 5067 19879 5109 19888
rect 4532 19468 4628 19508
rect 4492 19459 4532 19468
rect 4299 19340 4341 19349
rect 4299 19300 4300 19340
rect 4340 19300 4341 19340
rect 4299 19291 4341 19300
rect 4300 19256 4340 19291
rect 4300 19206 4340 19216
rect 4779 19256 4821 19265
rect 4779 19216 4780 19256
rect 4820 19216 4821 19256
rect 4779 19207 4821 19216
rect 4780 19122 4820 19207
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 4107 18668 4149 18677
rect 4107 18628 4108 18668
rect 4148 18628 4149 18668
rect 4107 18619 4149 18628
rect 5067 18668 5109 18677
rect 5067 18628 5068 18668
rect 5108 18628 5109 18668
rect 5067 18619 5109 18628
rect 4203 18584 4245 18593
rect 4203 18544 4204 18584
rect 4244 18544 4245 18584
rect 4203 18535 4245 18544
rect 4588 18584 4628 18593
rect 4204 18425 4244 18535
rect 4203 18416 4245 18425
rect 4203 18376 4204 18416
rect 4244 18376 4245 18416
rect 4203 18367 4245 18376
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 3916 17749 3956 17758
rect 3819 17660 3861 17669
rect 3916 17660 3956 17709
rect 4108 17660 4148 17669
rect 3819 17620 3820 17660
rect 3860 17620 3956 17660
rect 4012 17620 4108 17660
rect 3819 17611 3861 17620
rect 3532 17191 3572 17200
rect 3915 17240 3957 17249
rect 3915 17200 3916 17240
rect 3956 17200 3957 17240
rect 3915 17191 3957 17200
rect 3724 17081 3764 17166
rect 3916 17106 3956 17191
rect 3628 17072 3668 17081
rect 3436 17023 3476 17032
rect 3532 17032 3628 17072
rect 3335 16948 3380 16988
rect 3243 16904 3285 16913
rect 3335 16904 3375 16948
rect 3243 16864 3244 16904
rect 3284 16864 3375 16904
rect 3435 16904 3477 16913
rect 3435 16864 3436 16904
rect 3476 16864 3477 16904
rect 3243 16855 3285 16864
rect 3435 16855 3477 16864
rect 3339 16736 3381 16745
rect 3339 16696 3340 16736
rect 3380 16696 3381 16736
rect 3339 16687 3381 16696
rect 3340 15149 3380 16687
rect 3436 15476 3476 16855
rect 3532 16409 3572 17032
rect 3628 17023 3668 17032
rect 3723 17072 3765 17081
rect 3723 17032 3724 17072
rect 3764 17032 3765 17072
rect 3723 17023 3765 17032
rect 4012 16913 4052 17620
rect 4108 17611 4148 17620
rect 4107 17324 4149 17333
rect 4107 17284 4108 17324
rect 4148 17284 4149 17324
rect 4107 17275 4149 17284
rect 4108 17072 4148 17275
rect 4204 17249 4244 18367
rect 4588 18248 4628 18544
rect 4971 18584 5013 18593
rect 4971 18544 4972 18584
rect 5012 18544 5013 18584
rect 4971 18535 5013 18544
rect 4972 18450 5012 18535
rect 5068 18534 5108 18619
rect 5164 18584 5204 18593
rect 5356 18584 5396 18595
rect 5204 18544 5300 18584
rect 5164 18535 5204 18544
rect 4780 18332 4820 18341
rect 4300 18208 4628 18248
rect 4684 18292 4780 18332
rect 4300 17333 4340 18208
rect 4395 17996 4437 18005
rect 4395 17956 4396 17996
rect 4436 17956 4437 17996
rect 4395 17947 4437 17956
rect 4396 17744 4436 17947
rect 4396 17695 4436 17704
rect 4588 17744 4628 17753
rect 4492 17576 4532 17585
rect 4299 17324 4341 17333
rect 4299 17284 4300 17324
rect 4340 17284 4341 17324
rect 4299 17275 4341 17284
rect 4203 17240 4245 17249
rect 4203 17200 4204 17240
rect 4244 17200 4245 17240
rect 4203 17191 4245 17200
rect 4492 17081 4532 17536
rect 4588 17165 4628 17704
rect 4684 17744 4724 18292
rect 4780 18283 4820 18292
rect 5163 17828 5205 17837
rect 5163 17788 5164 17828
rect 5204 17788 5205 17828
rect 5163 17779 5205 17788
rect 4684 17585 4724 17704
rect 4875 17744 4917 17753
rect 4875 17704 4876 17744
rect 4916 17704 4917 17744
rect 4875 17695 4917 17704
rect 5067 17744 5109 17753
rect 5067 17704 5068 17744
rect 5108 17704 5109 17744
rect 5067 17695 5109 17704
rect 5164 17744 5204 17779
rect 4683 17576 4725 17585
rect 4683 17536 4684 17576
rect 4724 17536 4725 17576
rect 4683 17527 4725 17536
rect 4876 17576 4916 17695
rect 5068 17610 5108 17695
rect 5164 17693 5204 17704
rect 5260 17576 5300 18544
rect 5356 18509 5396 18544
rect 5355 18500 5397 18509
rect 5355 18460 5356 18500
rect 5396 18460 5397 18500
rect 5355 18451 5397 18460
rect 5452 18173 5492 20299
rect 5451 18164 5493 18173
rect 5451 18124 5452 18164
rect 5492 18124 5493 18164
rect 5451 18115 5493 18124
rect 5356 17753 5396 17838
rect 5451 17828 5493 17837
rect 5451 17788 5452 17828
rect 5492 17788 5493 17828
rect 5451 17779 5493 17788
rect 5355 17744 5397 17753
rect 5355 17704 5356 17744
rect 5396 17704 5397 17744
rect 5355 17695 5397 17704
rect 5260 17536 5396 17576
rect 4876 17527 4916 17536
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 5356 17240 5396 17536
rect 5260 17200 5396 17240
rect 4587 17156 4629 17165
rect 4587 17116 4588 17156
rect 4628 17116 4629 17156
rect 4587 17107 4629 17116
rect 4491 17072 4533 17081
rect 4148 17032 4244 17072
rect 4011 16904 4053 16913
rect 4011 16864 4012 16904
rect 4052 16864 4053 16904
rect 4011 16855 4053 16864
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 3627 16484 3669 16493
rect 4108 16484 4148 17032
rect 4204 16829 4244 17032
rect 4491 17032 4492 17072
rect 4532 17032 4533 17072
rect 4491 17023 4533 17032
rect 4203 16820 4245 16829
rect 4203 16780 4204 16820
rect 4244 16780 4245 16820
rect 4203 16771 4245 16780
rect 4299 16652 4341 16661
rect 4299 16612 4300 16652
rect 4340 16612 4341 16652
rect 4299 16603 4341 16612
rect 3627 16444 3628 16484
rect 3668 16444 3669 16484
rect 3627 16435 3669 16444
rect 4012 16444 4148 16484
rect 3531 16400 3573 16409
rect 3531 16360 3532 16400
rect 3572 16360 3573 16400
rect 3531 16351 3573 16360
rect 3532 16232 3572 16241
rect 3532 15989 3572 16192
rect 3531 15980 3573 15989
rect 3531 15940 3532 15980
rect 3572 15940 3573 15980
rect 3531 15931 3573 15940
rect 3628 15728 3668 16435
rect 3915 16400 3957 16409
rect 3915 16360 3916 16400
rect 3956 16360 3957 16400
rect 3915 16351 3957 16360
rect 3723 16148 3765 16157
rect 3723 16108 3724 16148
rect 3764 16108 3765 16148
rect 3723 16099 3765 16108
rect 3724 16014 3764 16099
rect 3916 16064 3956 16351
rect 3916 16015 3956 16024
rect 4012 15989 4052 16444
rect 4203 16400 4245 16409
rect 4203 16360 4204 16400
rect 4244 16360 4245 16400
rect 4203 16351 4245 16360
rect 4107 16232 4149 16241
rect 4107 16192 4108 16232
rect 4148 16192 4149 16232
rect 4107 16183 4149 16192
rect 4204 16232 4244 16351
rect 4204 16183 4244 16192
rect 4108 16098 4148 16183
rect 4011 15980 4053 15989
rect 4011 15940 4012 15980
rect 4052 15940 4053 15980
rect 4011 15931 4053 15940
rect 3628 15679 3668 15688
rect 3436 15427 3476 15436
rect 3916 15560 3956 15569
rect 3916 15308 3956 15520
rect 4011 15560 4053 15569
rect 4011 15520 4012 15560
rect 4052 15520 4053 15560
rect 4011 15511 4053 15520
rect 4012 15426 4052 15511
rect 3916 15268 4148 15308
rect 3339 15140 3381 15149
rect 3339 15100 3340 15140
rect 3380 15100 3381 15140
rect 3339 15091 3381 15100
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 2764 14848 3188 14888
rect 3244 14932 3668 14972
rect 2764 14804 2804 14848
rect 3244 14804 3284 14932
rect 3628 14888 3668 14932
rect 3628 14839 3668 14848
rect 4011 14888 4053 14897
rect 4011 14848 4012 14888
rect 4052 14848 4053 14888
rect 4011 14839 4053 14848
rect 2476 14671 2516 14680
rect 2572 14764 2804 14804
rect 3148 14764 3284 14804
rect 2475 11108 2517 11117
rect 2475 11068 2476 11108
rect 2516 11068 2517 11108
rect 2475 11059 2517 11068
rect 2476 11024 2516 11059
rect 2476 10193 2516 10984
rect 2475 10184 2517 10193
rect 2475 10144 2476 10184
rect 2516 10144 2517 10184
rect 2475 10135 2517 10144
rect 2379 8252 2421 8261
rect 2379 8212 2380 8252
rect 2420 8212 2421 8252
rect 2379 8203 2421 8212
rect 2572 7841 2612 14764
rect 3052 14720 3092 14729
rect 2955 14384 2997 14393
rect 2955 14344 2956 14384
rect 2996 14344 2997 14384
rect 2955 14335 2997 14344
rect 2956 14048 2996 14335
rect 2956 13999 2996 14008
rect 3052 13460 3092 14680
rect 3148 14384 3188 14764
rect 3532 14729 3572 14814
rect 3340 14720 3380 14729
rect 3243 14636 3285 14645
rect 3243 14596 3244 14636
rect 3284 14596 3285 14636
rect 3243 14587 3285 14596
rect 3244 14502 3284 14587
rect 3148 14344 3284 14384
rect 3147 14216 3189 14225
rect 3147 14176 3148 14216
rect 3188 14176 3189 14216
rect 3147 14167 3189 14176
rect 3148 14082 3188 14167
rect 3148 13460 3188 13469
rect 3052 13420 3148 13460
rect 3148 13411 3188 13420
rect 2955 13292 2997 13301
rect 2955 13252 2956 13292
rect 2996 13252 2997 13292
rect 2955 13243 2997 13252
rect 2956 13208 2996 13243
rect 2859 12620 2901 12629
rect 2859 12580 2860 12620
rect 2900 12580 2901 12620
rect 2859 12571 2901 12580
rect 2667 12452 2709 12461
rect 2667 12412 2668 12452
rect 2708 12412 2709 12452
rect 2667 12403 2709 12412
rect 2668 11192 2708 12403
rect 2860 12209 2900 12571
rect 2956 12536 2996 13168
rect 3147 13040 3189 13049
rect 3147 13000 3148 13040
rect 3188 13000 3189 13040
rect 3147 12991 3189 13000
rect 3148 12906 3188 12991
rect 2859 12200 2901 12209
rect 2859 12160 2860 12200
rect 2900 12160 2901 12200
rect 2859 12151 2901 12160
rect 2956 11696 2996 12496
rect 3147 12284 3189 12293
rect 3147 12244 3148 12284
rect 3188 12244 3189 12284
rect 3147 12235 3189 12244
rect 3148 12150 3188 12235
rect 3147 11948 3189 11957
rect 3147 11908 3148 11948
rect 3188 11908 3189 11948
rect 3147 11899 3189 11908
rect 3051 11864 3093 11873
rect 3051 11824 3052 11864
rect 3092 11824 3093 11864
rect 3051 11815 3093 11824
rect 2859 11276 2901 11285
rect 2859 11236 2860 11276
rect 2900 11236 2901 11276
rect 2859 11227 2901 11236
rect 2668 11143 2708 11152
rect 2860 11024 2900 11227
rect 2956 11033 2996 11656
rect 2860 10975 2900 10984
rect 2955 11024 2997 11033
rect 2955 10984 2956 11024
rect 2996 10984 2997 11024
rect 2955 10975 2997 10984
rect 2668 10436 2708 10445
rect 2708 10396 2900 10436
rect 2668 10387 2708 10396
rect 2860 10184 2900 10396
rect 2860 10135 2900 10144
rect 3052 10184 3092 11815
rect 3148 11814 3188 11899
rect 3244 11705 3284 14344
rect 3340 12713 3380 14680
rect 3531 14720 3573 14729
rect 3531 14680 3532 14720
rect 3572 14680 3573 14720
rect 3531 14671 3573 14680
rect 3723 14720 3765 14729
rect 3723 14680 3724 14720
rect 3764 14680 3765 14720
rect 3723 14671 3765 14680
rect 3820 14720 3860 14729
rect 3435 14636 3477 14645
rect 3435 14596 3436 14636
rect 3476 14596 3477 14636
rect 3435 14587 3477 14596
rect 3436 14300 3476 14587
rect 3724 14586 3764 14671
rect 3820 14309 3860 14680
rect 4012 14720 4052 14839
rect 4012 14671 4052 14680
rect 4011 14552 4053 14561
rect 4011 14512 4012 14552
rect 4052 14512 4053 14552
rect 4011 14503 4053 14512
rect 3819 14300 3861 14309
rect 3436 14260 3668 14300
rect 3531 14048 3573 14057
rect 3531 14008 3532 14048
rect 3572 14008 3573 14048
rect 3531 13999 3573 14008
rect 3628 14048 3668 14260
rect 3819 14260 3820 14300
rect 3860 14260 3861 14300
rect 3819 14251 3861 14260
rect 3628 13999 3668 14008
rect 3724 14048 3764 14057
rect 3532 13914 3572 13999
rect 3724 13796 3764 14008
rect 3819 14048 3861 14057
rect 3819 14008 3820 14048
rect 3860 14008 3861 14048
rect 3819 13999 3861 14008
rect 4012 14048 4052 14503
rect 4108 14225 4148 15268
rect 4300 14897 4340 16603
rect 4588 16409 4628 17107
rect 5260 16484 5300 17200
rect 5356 17072 5396 17081
rect 5356 16661 5396 17032
rect 5355 16652 5397 16661
rect 5355 16612 5356 16652
rect 5396 16612 5397 16652
rect 5355 16603 5397 16612
rect 5260 16435 5300 16444
rect 4587 16400 4629 16409
rect 4587 16360 4588 16400
rect 4628 16360 4629 16400
rect 4587 16351 4629 16360
rect 4875 16400 4917 16409
rect 4875 16360 4876 16400
rect 4916 16360 4917 16400
rect 4875 16351 4917 16360
rect 4587 16232 4629 16241
rect 4587 16192 4588 16232
rect 4628 16192 4629 16232
rect 4587 16183 4629 16192
rect 4876 16232 4916 16351
rect 5452 16241 5492 17779
rect 5548 17669 5588 21391
rect 5644 20096 5684 20105
rect 5644 19853 5684 20056
rect 5740 19937 5780 22912
rect 6027 22868 6069 22877
rect 6027 22828 6028 22868
rect 6068 22828 6069 22868
rect 6027 22819 6069 22828
rect 5836 22285 5876 22294
rect 5836 21785 5876 22245
rect 5931 22028 5973 22037
rect 5931 21988 5932 22028
rect 5972 21988 5973 22028
rect 5931 21979 5973 21988
rect 5835 21776 5877 21785
rect 5835 21736 5836 21776
rect 5876 21736 5877 21776
rect 5835 21727 5877 21736
rect 5739 19928 5781 19937
rect 5739 19888 5740 19928
rect 5780 19888 5781 19928
rect 5739 19879 5781 19888
rect 5643 19844 5685 19853
rect 5643 19804 5644 19844
rect 5684 19804 5685 19844
rect 5643 19795 5685 19804
rect 5643 18668 5685 18677
rect 5643 18628 5644 18668
rect 5684 18628 5685 18668
rect 5643 18619 5685 18628
rect 5644 18584 5684 18619
rect 5644 18533 5684 18544
rect 5643 18416 5685 18425
rect 5643 18376 5644 18416
rect 5684 18376 5685 18416
rect 5643 18367 5685 18376
rect 5644 18282 5684 18367
rect 5547 17660 5589 17669
rect 5547 17620 5548 17660
rect 5588 17620 5589 17660
rect 5547 17611 5589 17620
rect 4876 16183 4916 16192
rect 5451 16232 5493 16241
rect 5451 16192 5452 16232
rect 5492 16192 5493 16232
rect 5451 16183 5493 16192
rect 5548 16232 5588 16241
rect 4588 16098 4628 16183
rect 4972 16148 5012 16157
rect 4972 16064 5012 16108
rect 4684 16024 5012 16064
rect 4491 15980 4533 15989
rect 4491 15940 4492 15980
rect 4532 15940 4533 15980
rect 4491 15931 4533 15940
rect 4492 15560 4532 15931
rect 4492 15511 4532 15520
rect 4396 15476 4436 15485
rect 4396 15317 4436 15436
rect 4395 15308 4437 15317
rect 4395 15268 4396 15308
rect 4436 15268 4437 15308
rect 4395 15259 4437 15268
rect 4299 14888 4341 14897
rect 4299 14848 4300 14888
rect 4340 14848 4341 14888
rect 4299 14839 4341 14848
rect 4396 14561 4436 15259
rect 4395 14552 4437 14561
rect 4395 14512 4396 14552
rect 4436 14512 4437 14552
rect 4395 14503 4437 14512
rect 4587 14468 4629 14477
rect 4587 14428 4588 14468
rect 4628 14428 4629 14468
rect 4587 14419 4629 14428
rect 4588 14225 4628 14419
rect 4107 14216 4149 14225
rect 4107 14176 4108 14216
rect 4148 14176 4149 14216
rect 4107 14167 4149 14176
rect 4587 14216 4629 14225
rect 4587 14176 4588 14216
rect 4628 14176 4629 14216
rect 4587 14167 4629 14176
rect 3820 13914 3860 13999
rect 4012 13973 4052 14008
rect 4396 14048 4436 14057
rect 4684 14048 4724 16024
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 5548 15653 5588 16192
rect 5547 15644 5589 15653
rect 5547 15604 5548 15644
rect 5588 15604 5589 15644
rect 5547 15595 5589 15604
rect 5644 15644 5684 15653
rect 4972 15560 5012 15569
rect 4972 15401 5012 15520
rect 5452 15546 5492 15555
rect 4971 15392 5013 15401
rect 4971 15352 4972 15392
rect 5012 15352 5013 15392
rect 4971 15343 5013 15352
rect 5452 14972 5492 15506
rect 5644 15485 5684 15604
rect 5643 15476 5685 15485
rect 5643 15436 5644 15476
rect 5684 15436 5685 15476
rect 5740 15476 5780 19879
rect 5932 18752 5972 21979
rect 6028 19928 6068 22819
rect 6124 21533 6164 24331
rect 6220 23801 6260 29623
rect 6315 29168 6357 29177
rect 6315 29128 6316 29168
rect 6356 29128 6357 29168
rect 6315 29119 6357 29128
rect 6316 28328 6356 29119
rect 6316 28279 6356 28288
rect 6412 28076 6452 29800
rect 6508 29791 6548 29800
rect 6603 29840 6645 29849
rect 6603 29800 6604 29840
rect 6644 29800 6645 29840
rect 6603 29791 6645 29800
rect 6700 29177 6740 30295
rect 6892 29924 6932 30892
rect 6988 30680 7028 30689
rect 6988 30269 7028 30640
rect 7084 30680 7124 30689
rect 6987 30260 7029 30269
rect 6987 30220 6988 30260
rect 7028 30220 7029 30260
rect 6987 30211 7029 30220
rect 7084 30101 7124 30640
rect 7180 30680 7220 30689
rect 7180 30185 7220 30640
rect 7275 30680 7317 30689
rect 7275 30640 7276 30680
rect 7316 30640 7317 30680
rect 7275 30631 7317 30640
rect 7276 30546 7316 30631
rect 7372 30605 7412 31312
rect 7371 30596 7413 30605
rect 7371 30556 7372 30596
rect 7412 30556 7413 30596
rect 7371 30547 7413 30556
rect 7179 30176 7221 30185
rect 7179 30136 7180 30176
rect 7220 30136 7221 30176
rect 7179 30127 7221 30136
rect 7083 30092 7125 30101
rect 7083 30052 7084 30092
rect 7124 30052 7125 30092
rect 7083 30043 7125 30052
rect 6892 29884 7124 29924
rect 6892 29252 6932 29261
rect 6699 29168 6741 29177
rect 6699 29128 6700 29168
rect 6740 29128 6741 29168
rect 6892 29168 6932 29212
rect 6987 29168 7029 29177
rect 6892 29128 6988 29168
rect 7028 29128 7029 29168
rect 6699 29119 6741 29128
rect 6987 29119 7029 29128
rect 6700 29034 6740 29119
rect 7084 28580 7124 29884
rect 7276 29840 7316 29849
rect 7276 29429 7316 29800
rect 7275 29420 7317 29429
rect 7275 29380 7276 29420
rect 7316 29380 7317 29420
rect 7275 29371 7317 29380
rect 7468 29177 7508 31900
rect 7179 29168 7221 29177
rect 7179 29128 7180 29168
rect 7220 29128 7221 29168
rect 7179 29119 7221 29128
rect 7276 29168 7316 29177
rect 7180 29034 7220 29119
rect 7276 29000 7316 29128
rect 7467 29168 7509 29177
rect 7467 29128 7468 29168
rect 7508 29128 7509 29168
rect 7467 29119 7509 29128
rect 7276 28960 7412 29000
rect 7084 28540 7316 28580
rect 6891 28496 6933 28505
rect 6891 28456 6892 28496
rect 6932 28456 6933 28496
rect 6891 28447 6933 28456
rect 6796 28328 6836 28337
rect 6508 28244 6548 28253
rect 6796 28244 6836 28288
rect 6548 28204 6836 28244
rect 6892 28328 6932 28447
rect 7276 28337 7316 28540
rect 6508 28195 6548 28204
rect 6412 28036 6740 28076
rect 6507 27740 6549 27749
rect 6507 27700 6508 27740
rect 6548 27700 6549 27740
rect 6507 27691 6549 27700
rect 6316 27656 6356 27665
rect 6316 27077 6356 27616
rect 6412 27656 6452 27665
rect 6315 27068 6357 27077
rect 6315 27028 6316 27068
rect 6356 27028 6357 27068
rect 6315 27019 6357 27028
rect 6412 25733 6452 27616
rect 6508 27606 6548 27691
rect 6604 27656 6644 27665
rect 6604 27413 6644 27616
rect 6603 27404 6645 27413
rect 6603 27364 6604 27404
rect 6644 27364 6645 27404
rect 6603 27355 6645 27364
rect 6507 27320 6549 27329
rect 6507 27280 6508 27320
rect 6548 27280 6549 27320
rect 6507 27271 6549 27280
rect 6411 25724 6453 25733
rect 6411 25684 6412 25724
rect 6452 25684 6453 25724
rect 6411 25675 6453 25684
rect 6508 25220 6548 27271
rect 6603 27236 6645 27245
rect 6603 27196 6604 27236
rect 6644 27196 6645 27236
rect 6603 27187 6645 27196
rect 6412 25180 6548 25220
rect 6315 25052 6357 25061
rect 6315 25012 6316 25052
rect 6356 25012 6357 25052
rect 6315 25003 6357 25012
rect 6219 23792 6261 23801
rect 6219 23752 6220 23792
rect 6260 23752 6261 23792
rect 6219 23743 6261 23752
rect 6316 22280 6356 25003
rect 6316 22231 6356 22240
rect 6219 21608 6261 21617
rect 6219 21568 6220 21608
rect 6260 21568 6261 21608
rect 6219 21559 6261 21568
rect 6123 21524 6165 21533
rect 6123 21484 6124 21524
rect 6164 21484 6165 21524
rect 6123 21475 6165 21484
rect 6220 20348 6260 21559
rect 6412 20693 6452 25180
rect 6604 23297 6644 27187
rect 6700 26480 6740 28036
rect 6796 27665 6836 27750
rect 6795 27656 6837 27665
rect 6795 27616 6796 27656
rect 6836 27616 6837 27656
rect 6795 27607 6837 27616
rect 6892 26489 6932 28288
rect 6987 28328 7029 28337
rect 6987 28288 6988 28328
rect 7028 28288 7029 28328
rect 6987 28279 7029 28288
rect 7275 28328 7317 28337
rect 7275 28288 7276 28328
rect 7316 28288 7317 28328
rect 7275 28279 7317 28288
rect 7372 28328 7412 28960
rect 6891 26480 6933 26489
rect 6700 26440 6836 26480
rect 6700 26144 6740 26153
rect 6700 24641 6740 26104
rect 6796 25136 6836 26440
rect 6891 26440 6892 26480
rect 6932 26440 6933 26480
rect 6891 26431 6933 26440
rect 6892 25892 6932 25901
rect 6892 25304 6932 25852
rect 6988 25481 7028 28279
rect 7179 28244 7221 28253
rect 7179 28204 7180 28244
rect 7220 28204 7221 28244
rect 7179 28195 7221 28204
rect 7084 26144 7124 26153
rect 7084 25985 7124 26104
rect 7083 25976 7125 25985
rect 7083 25936 7084 25976
rect 7124 25936 7125 25976
rect 7083 25927 7125 25936
rect 6987 25472 7029 25481
rect 6987 25432 6988 25472
rect 7028 25432 7029 25472
rect 6987 25423 7029 25432
rect 6988 25304 7028 25313
rect 6892 25264 6988 25304
rect 6988 25255 7028 25264
rect 7083 25304 7125 25313
rect 7083 25264 7084 25304
rect 7124 25264 7125 25304
rect 7083 25255 7125 25264
rect 7084 25170 7124 25255
rect 6796 25096 7028 25136
rect 6699 24632 6741 24641
rect 6699 24592 6700 24632
rect 6740 24592 6741 24632
rect 6699 24583 6741 24592
rect 6891 23960 6933 23969
rect 6891 23920 6892 23960
rect 6932 23920 6933 23960
rect 6891 23911 6933 23920
rect 6603 23288 6645 23297
rect 6603 23248 6604 23288
rect 6644 23248 6645 23288
rect 6603 23239 6645 23248
rect 6795 23288 6837 23297
rect 6795 23248 6796 23288
rect 6836 23248 6837 23288
rect 6795 23239 6837 23248
rect 6507 23204 6549 23213
rect 6507 23164 6508 23204
rect 6548 23164 6549 23204
rect 6507 23155 6549 23164
rect 6508 23120 6548 23155
rect 6508 23069 6548 23080
rect 6796 23120 6836 23239
rect 6796 23071 6836 23080
rect 6892 23120 6932 23911
rect 6892 22961 6932 23080
rect 6891 22952 6933 22961
rect 6891 22912 6892 22952
rect 6932 22912 6933 22952
rect 6891 22903 6933 22912
rect 6507 22700 6549 22709
rect 6507 22660 6508 22700
rect 6548 22660 6549 22700
rect 6507 22651 6549 22660
rect 6508 21617 6548 22651
rect 6603 22280 6645 22289
rect 6796 22280 6836 22289
rect 6603 22240 6604 22280
rect 6644 22240 6796 22280
rect 6603 22231 6645 22240
rect 6796 22231 6836 22240
rect 6892 22280 6932 22291
rect 6507 21608 6549 21617
rect 6507 21568 6508 21608
rect 6548 21568 6549 21608
rect 6507 21559 6549 21568
rect 6411 20684 6453 20693
rect 6411 20644 6412 20684
rect 6452 20644 6453 20684
rect 6411 20635 6453 20644
rect 6220 20308 6452 20348
rect 6123 20264 6165 20273
rect 6123 20224 6124 20264
rect 6164 20224 6165 20264
rect 6123 20215 6165 20224
rect 6124 20091 6164 20215
rect 6124 20042 6164 20051
rect 6316 20180 6356 20189
rect 6028 19888 6164 19928
rect 6124 19685 6164 19888
rect 6123 19676 6165 19685
rect 6123 19636 6124 19676
rect 6164 19636 6165 19676
rect 6123 19627 6165 19636
rect 6027 19340 6069 19349
rect 6027 19300 6028 19340
rect 6068 19300 6069 19340
rect 6027 19291 6069 19300
rect 6028 19256 6068 19291
rect 6028 19097 6068 19216
rect 6027 19088 6069 19097
rect 6027 19048 6028 19088
rect 6068 19048 6069 19088
rect 6027 19039 6069 19048
rect 6124 18752 6164 19627
rect 6219 19508 6261 19517
rect 6219 19468 6220 19508
rect 6260 19468 6261 19508
rect 6219 19459 6261 19468
rect 6220 19374 6260 19459
rect 6316 18836 6356 20140
rect 6412 19769 6452 20308
rect 6411 19760 6453 19769
rect 6411 19720 6412 19760
rect 6452 19720 6453 19760
rect 6411 19711 6453 19720
rect 6604 18920 6644 22231
rect 6892 22205 6932 22240
rect 6891 22196 6933 22205
rect 6891 22156 6892 22196
rect 6932 22156 6933 22196
rect 6891 22147 6933 22156
rect 6795 22112 6837 22121
rect 6795 22072 6796 22112
rect 6836 22072 6837 22112
rect 6795 22063 6837 22072
rect 6699 21608 6741 21617
rect 6699 21568 6700 21608
rect 6740 21568 6741 21608
rect 6699 21559 6741 21568
rect 6700 20768 6740 21559
rect 6796 21020 6836 22063
rect 6891 21776 6933 21785
rect 6891 21736 6892 21776
rect 6932 21736 6933 21776
rect 6891 21727 6933 21736
rect 6892 21642 6932 21727
rect 6891 21524 6933 21533
rect 6891 21484 6892 21524
rect 6932 21484 6933 21524
rect 6891 21475 6933 21484
rect 6892 21272 6932 21475
rect 6988 21449 7028 25096
rect 7083 23120 7125 23129
rect 7083 23080 7084 23120
rect 7124 23080 7125 23120
rect 7083 23071 7125 23080
rect 6987 21440 7029 21449
rect 6987 21400 6988 21440
rect 7028 21400 7029 21440
rect 7084 21440 7124 23071
rect 7180 23045 7220 28195
rect 7276 28194 7316 28279
rect 7275 27656 7317 27665
rect 7275 27616 7276 27656
rect 7316 27616 7317 27656
rect 7275 27607 7317 27616
rect 7276 26816 7316 27607
rect 7372 26825 7412 28288
rect 7468 26909 7508 29119
rect 7564 28505 7604 32824
rect 7660 32789 7700 33823
rect 7756 33704 7796 34075
rect 7659 32780 7701 32789
rect 7659 32740 7660 32780
rect 7700 32740 7701 32780
rect 7659 32731 7701 32740
rect 7756 32612 7796 33664
rect 7660 32572 7796 32612
rect 7660 31940 7700 32572
rect 7755 32192 7797 32201
rect 7755 32152 7756 32192
rect 7796 32152 7797 32192
rect 7755 32143 7797 32152
rect 7852 32192 7892 34915
rect 8044 34376 8084 34385
rect 7948 34208 7988 34217
rect 7948 33041 7988 34168
rect 8044 34133 8084 34336
rect 8043 34124 8085 34133
rect 8043 34084 8044 34124
rect 8084 34084 8085 34124
rect 8043 34075 8085 34084
rect 7947 33032 7989 33041
rect 7947 32992 7948 33032
rect 7988 32992 7989 33032
rect 7947 32983 7989 32992
rect 8043 32948 8085 32957
rect 8043 32908 8044 32948
rect 8084 32908 8085 32948
rect 8043 32899 8085 32908
rect 7948 32864 7988 32875
rect 7948 32789 7988 32824
rect 8044 32814 8084 32899
rect 7947 32780 7989 32789
rect 7947 32740 7948 32780
rect 7988 32740 7989 32780
rect 7947 32731 7989 32740
rect 7852 32143 7892 32152
rect 7756 32058 7796 32143
rect 7660 31900 7892 31940
rect 7659 31184 7701 31193
rect 7659 31144 7660 31184
rect 7700 31144 7701 31184
rect 7659 31135 7701 31144
rect 7660 30680 7700 31135
rect 7852 30857 7892 31900
rect 7851 30848 7893 30857
rect 7851 30808 7852 30848
rect 7892 30808 7893 30848
rect 7851 30799 7893 30808
rect 7851 30680 7893 30689
rect 7660 30631 7700 30640
rect 7756 30661 7852 30680
rect 7796 30640 7852 30661
rect 7892 30640 7893 30680
rect 7851 30631 7893 30640
rect 7756 30612 7796 30621
rect 7948 30512 7988 32731
rect 8043 32360 8085 32369
rect 8043 32320 8044 32360
rect 8084 32320 8085 32360
rect 8043 32311 8085 32320
rect 8044 32226 8084 32311
rect 8043 31352 8085 31361
rect 8043 31312 8044 31352
rect 8084 31312 8085 31352
rect 8043 31303 8085 31312
rect 7756 30472 7988 30512
rect 7659 29168 7701 29177
rect 7659 29128 7660 29168
rect 7700 29128 7701 29168
rect 7659 29119 7701 29128
rect 7756 29168 7796 30472
rect 8044 30269 8084 31303
rect 8139 31268 8181 31277
rect 8139 31228 8140 31268
rect 8180 31228 8181 31268
rect 8139 31219 8181 31228
rect 8140 31025 8180 31219
rect 8139 31016 8181 31025
rect 8139 30976 8140 31016
rect 8180 30976 8181 31016
rect 8139 30967 8181 30976
rect 8140 30680 8180 30967
rect 8140 30631 8180 30640
rect 8236 30596 8276 34999
rect 8523 34964 8565 34973
rect 8523 34924 8524 34964
rect 8564 34924 8565 34964
rect 8523 34915 8565 34924
rect 8524 34830 8564 34915
rect 8523 34628 8565 34637
rect 8523 34588 8524 34628
rect 8564 34588 8565 34628
rect 8523 34579 8565 34588
rect 8332 34460 8372 34469
rect 8524 34460 8564 34579
rect 8372 34420 8564 34460
rect 8332 34411 8372 34420
rect 8524 34376 8564 34420
rect 8524 34327 8564 34336
rect 8331 33032 8373 33041
rect 8331 32992 8332 33032
rect 8372 32992 8373 33032
rect 8331 32983 8373 32992
rect 8043 30260 8085 30269
rect 8043 30220 8044 30260
rect 8084 30220 8085 30260
rect 8043 30211 8085 30220
rect 7851 29840 7893 29849
rect 7851 29800 7852 29840
rect 7892 29800 7893 29840
rect 7851 29791 7893 29800
rect 7660 29034 7700 29119
rect 7563 28496 7605 28505
rect 7563 28456 7564 28496
rect 7604 28456 7605 28496
rect 7563 28447 7605 28456
rect 7756 27245 7796 29128
rect 7852 28328 7892 29791
rect 7852 27404 7892 28288
rect 8044 27665 8084 30211
rect 8236 29765 8276 30556
rect 8332 30521 8372 32983
rect 8524 32864 8564 32875
rect 8524 32789 8564 32824
rect 8523 32780 8565 32789
rect 8523 32740 8524 32780
rect 8564 32740 8565 32780
rect 8523 32731 8565 32740
rect 8427 32444 8469 32453
rect 8427 32404 8428 32444
rect 8468 32404 8469 32444
rect 8427 32395 8469 32404
rect 8428 32192 8468 32395
rect 8428 32143 8468 32152
rect 8523 31352 8565 31361
rect 8523 31312 8524 31352
rect 8564 31312 8565 31352
rect 8523 31303 8565 31312
rect 8524 31218 8564 31303
rect 8620 31025 8660 35251
rect 9004 35048 9044 35680
rect 9100 35225 9140 39535
rect 9484 37820 9524 39712
rect 9676 38585 9716 39880
rect 9963 39752 10005 39761
rect 9963 39712 9964 39752
rect 10004 39712 10005 39752
rect 9963 39703 10005 39712
rect 9867 39668 9909 39677
rect 9867 39628 9868 39668
rect 9908 39628 9909 39668
rect 9867 39619 9909 39628
rect 9868 39534 9908 39619
rect 9964 39618 10004 39703
rect 9675 38576 9717 38585
rect 9675 38536 9676 38576
rect 9716 38536 9717 38576
rect 9675 38527 9717 38536
rect 9675 38240 9717 38249
rect 9675 38200 9676 38240
rect 9716 38200 9717 38240
rect 9675 38191 9717 38200
rect 9868 38240 9908 38249
rect 9676 38106 9716 38191
rect 9772 37988 9812 37997
rect 9772 37820 9812 37948
rect 9292 37780 9524 37820
rect 9676 37780 9812 37820
rect 9195 37400 9237 37409
rect 9195 37360 9196 37400
rect 9236 37360 9237 37400
rect 9195 37351 9237 37360
rect 9196 36065 9236 37351
rect 9195 36056 9237 36065
rect 9195 36016 9196 36056
rect 9236 36016 9237 36056
rect 9195 36007 9237 36016
rect 9099 35216 9141 35225
rect 9099 35176 9100 35216
rect 9140 35176 9141 35216
rect 9099 35167 9141 35176
rect 9195 35132 9237 35141
rect 9195 35092 9196 35132
rect 9236 35092 9237 35132
rect 9195 35083 9237 35092
rect 8908 35008 9004 35048
rect 8811 33704 8853 33713
rect 8811 33664 8812 33704
rect 8852 33664 8853 33704
rect 8811 33655 8853 33664
rect 8812 32117 8852 33655
rect 8908 32780 8948 35008
rect 9004 34999 9044 35008
rect 9196 34133 9236 35083
rect 9195 34124 9237 34133
rect 9195 34084 9196 34124
rect 9236 34084 9237 34124
rect 9195 34075 9237 34084
rect 9003 33704 9045 33713
rect 9003 33664 9004 33704
rect 9044 33664 9045 33704
rect 9003 33655 9045 33664
rect 9004 33570 9044 33655
rect 9196 33452 9236 33461
rect 9196 32948 9236 33412
rect 9052 32908 9236 32948
rect 9052 32906 9092 32908
rect 9052 32857 9092 32866
rect 8908 32740 9044 32780
rect 8811 32108 8853 32117
rect 8811 32068 8812 32108
rect 8852 32068 8853 32108
rect 8811 32059 8853 32068
rect 8811 31520 8853 31529
rect 8811 31480 8812 31520
rect 8852 31480 8853 31520
rect 8811 31471 8853 31480
rect 8715 31184 8757 31193
rect 8715 31144 8716 31184
rect 8756 31144 8757 31184
rect 8715 31135 8757 31144
rect 8716 31050 8756 31135
rect 8619 31016 8661 31025
rect 8619 30976 8620 31016
rect 8660 30976 8661 31016
rect 8619 30967 8661 30976
rect 8716 30680 8756 30689
rect 8331 30512 8373 30521
rect 8331 30472 8332 30512
rect 8372 30472 8373 30512
rect 8331 30463 8373 30472
rect 8235 29756 8277 29765
rect 8235 29716 8236 29756
rect 8276 29716 8277 29756
rect 8235 29707 8277 29716
rect 8236 29345 8276 29707
rect 8235 29336 8277 29345
rect 8235 29296 8236 29336
rect 8276 29296 8277 29336
rect 8235 29287 8277 29296
rect 8235 29168 8277 29177
rect 8332 29168 8372 30463
rect 8523 30176 8565 30185
rect 8523 30136 8524 30176
rect 8564 30136 8565 30176
rect 8523 30127 8565 30136
rect 8524 29840 8564 30127
rect 8619 30092 8661 30101
rect 8619 30052 8620 30092
rect 8660 30052 8661 30092
rect 8619 30043 8661 30052
rect 8524 29791 8564 29800
rect 8235 29128 8236 29168
rect 8276 29128 8372 29168
rect 8235 29119 8277 29128
rect 8236 29034 8276 29119
rect 8332 28333 8372 28342
rect 8236 27824 8276 27833
rect 8332 27824 8372 28293
rect 8276 27784 8372 27824
rect 8524 28160 8564 28169
rect 8236 27775 8276 27784
rect 8043 27656 8085 27665
rect 8428 27656 8468 27665
rect 8043 27616 8044 27656
rect 8084 27616 8180 27656
rect 8043 27607 8085 27616
rect 8044 27522 8084 27607
rect 7852 27364 8084 27404
rect 7755 27236 7797 27245
rect 7755 27196 7756 27236
rect 7796 27196 7797 27236
rect 7755 27187 7797 27196
rect 7947 27152 7989 27161
rect 7947 27112 7948 27152
rect 7988 27112 7989 27152
rect 7947 27103 7989 27112
rect 7467 26900 7509 26909
rect 7467 26860 7468 26900
rect 7508 26860 7509 26900
rect 7467 26851 7509 26860
rect 7276 26767 7316 26776
rect 7371 26816 7413 26825
rect 7371 26776 7372 26816
rect 7412 26776 7413 26816
rect 7371 26767 7413 26776
rect 7756 26816 7796 26825
rect 7468 26732 7508 26741
rect 7756 26732 7796 26776
rect 7508 26692 7796 26732
rect 7852 26816 7892 26825
rect 7468 26683 7508 26692
rect 7275 26648 7317 26657
rect 7275 26608 7276 26648
rect 7316 26608 7317 26648
rect 7275 26599 7317 26608
rect 7276 25220 7316 26599
rect 7852 26489 7892 26776
rect 7851 26480 7893 26489
rect 7851 26440 7852 26480
rect 7892 26440 7893 26480
rect 7851 26431 7893 26440
rect 7468 25304 7508 25313
rect 7468 25220 7508 25264
rect 7564 25304 7604 25315
rect 7564 25229 7604 25264
rect 7755 25304 7797 25313
rect 7852 25304 7892 26431
rect 7755 25264 7756 25304
rect 7796 25264 7892 25304
rect 7755 25255 7797 25264
rect 7276 25180 7508 25220
rect 7563 25220 7605 25229
rect 7563 25180 7564 25220
rect 7604 25180 7605 25220
rect 7276 23969 7316 25180
rect 7563 25171 7605 25180
rect 7563 24800 7605 24809
rect 7563 24760 7564 24800
rect 7604 24760 7605 24800
rect 7563 24751 7605 24760
rect 7564 24666 7604 24751
rect 7756 24641 7796 25255
rect 7948 24800 7988 27103
rect 8044 25304 8084 27364
rect 8140 26144 8180 27616
rect 8428 27497 8468 27616
rect 8427 27488 8469 27497
rect 8427 27448 8428 27488
rect 8468 27448 8469 27488
rect 8427 27439 8469 27448
rect 8235 27236 8277 27245
rect 8235 27196 8236 27236
rect 8276 27196 8277 27236
rect 8235 27187 8277 27196
rect 8236 26900 8276 27187
rect 8524 26909 8564 28120
rect 8236 26851 8276 26860
rect 8523 26900 8565 26909
rect 8523 26860 8524 26900
rect 8564 26860 8565 26900
rect 8523 26851 8565 26860
rect 8331 26816 8373 26825
rect 8331 26776 8332 26816
rect 8372 26776 8468 26816
rect 8331 26767 8373 26776
rect 8332 26682 8372 26767
rect 8331 26144 8373 26153
rect 8140 26104 8332 26144
rect 8372 26104 8373 26144
rect 8331 26095 8373 26104
rect 8332 26010 8372 26095
rect 8331 25808 8373 25817
rect 8331 25768 8332 25808
rect 8372 25768 8373 25808
rect 8331 25759 8373 25768
rect 8084 25264 8180 25304
rect 8044 25255 8084 25264
rect 7948 24760 8084 24800
rect 7371 24632 7413 24641
rect 7371 24592 7372 24632
rect 7412 24592 7413 24632
rect 7371 24583 7413 24592
rect 7755 24632 7797 24641
rect 7755 24592 7756 24632
rect 7796 24592 7797 24632
rect 7755 24583 7797 24592
rect 7852 24632 7892 24641
rect 7372 24498 7412 24583
rect 7852 23969 7892 24592
rect 7947 24632 7989 24641
rect 7947 24592 7948 24632
rect 7988 24592 7989 24632
rect 7947 24583 7989 24592
rect 7948 24498 7988 24583
rect 7947 24212 7989 24221
rect 7947 24172 7948 24212
rect 7988 24172 7989 24212
rect 7947 24163 7989 24172
rect 7275 23960 7317 23969
rect 7275 23920 7276 23960
rect 7316 23920 7317 23960
rect 7275 23911 7317 23920
rect 7467 23960 7509 23969
rect 7467 23920 7468 23960
rect 7508 23920 7509 23960
rect 7467 23911 7509 23920
rect 7851 23960 7893 23969
rect 7851 23920 7852 23960
rect 7892 23920 7893 23960
rect 7851 23911 7893 23920
rect 7468 23826 7508 23911
rect 7276 23792 7316 23801
rect 7276 23717 7316 23752
rect 7948 23792 7988 24163
rect 7275 23708 7317 23717
rect 7275 23668 7276 23708
rect 7316 23668 7317 23708
rect 7275 23659 7317 23668
rect 7276 23657 7316 23659
rect 7948 23381 7988 23752
rect 7947 23372 7989 23381
rect 7276 23332 7508 23372
rect 7179 23036 7221 23045
rect 7179 22996 7180 23036
rect 7220 22996 7221 23036
rect 7179 22987 7221 22996
rect 7180 22868 7220 22877
rect 7180 22289 7220 22828
rect 7276 22457 7316 23332
rect 7468 23120 7508 23332
rect 7947 23332 7948 23372
rect 7988 23332 7989 23372
rect 7947 23323 7989 23332
rect 7563 23204 7605 23213
rect 7563 23164 7564 23204
rect 7604 23164 7605 23204
rect 7563 23155 7605 23164
rect 7468 23071 7508 23080
rect 7564 23070 7604 23155
rect 7948 23129 7988 23214
rect 7660 23120 7700 23129
rect 7467 22952 7509 22961
rect 7467 22912 7468 22952
rect 7508 22912 7509 22952
rect 7467 22903 7509 22912
rect 7468 22709 7508 22903
rect 7467 22700 7509 22709
rect 7467 22660 7468 22700
rect 7508 22660 7509 22700
rect 7467 22651 7509 22660
rect 7275 22448 7317 22457
rect 7275 22408 7276 22448
rect 7316 22408 7317 22448
rect 7275 22399 7317 22408
rect 7371 22364 7413 22373
rect 7371 22324 7372 22364
rect 7412 22324 7413 22364
rect 7371 22315 7413 22324
rect 7372 22299 7412 22315
rect 7179 22280 7221 22289
rect 7179 22240 7180 22280
rect 7220 22240 7221 22280
rect 7179 22231 7221 22240
rect 7276 22280 7316 22289
rect 7276 22037 7316 22240
rect 7275 22028 7317 22037
rect 7275 21988 7276 22028
rect 7316 21988 7317 22028
rect 7275 21979 7317 21988
rect 7179 21860 7221 21869
rect 7179 21820 7180 21860
rect 7220 21820 7221 21860
rect 7179 21811 7221 21820
rect 7180 21608 7220 21811
rect 7180 21559 7220 21568
rect 7276 21524 7316 21979
rect 7372 21869 7412 22259
rect 7660 22112 7700 23080
rect 7756 23120 7796 23129
rect 7756 22952 7796 23080
rect 7947 23120 7989 23129
rect 7947 23080 7948 23120
rect 7988 23080 7989 23120
rect 7947 23071 7989 23080
rect 7948 22952 7988 22961
rect 7756 22912 7948 22952
rect 7948 22903 7988 22912
rect 8044 22784 8084 24760
rect 8140 24464 8180 25264
rect 8332 24632 8372 25759
rect 8428 25229 8468 26776
rect 8523 26312 8565 26321
rect 8523 26272 8524 26312
rect 8564 26272 8565 26312
rect 8523 26263 8565 26272
rect 8524 26178 8564 26263
rect 8524 25309 8564 25318
rect 8427 25220 8469 25229
rect 8427 25180 8428 25220
rect 8468 25180 8469 25220
rect 8427 25171 8469 25180
rect 8332 24583 8372 24592
rect 8428 24548 8468 25171
rect 8524 24809 8564 25269
rect 8523 24800 8565 24809
rect 8523 24760 8524 24800
rect 8564 24760 8565 24800
rect 8523 24751 8565 24760
rect 8468 24508 8564 24548
rect 8428 24499 8468 24508
rect 8140 24424 8372 24464
rect 7660 22063 7700 22072
rect 7756 22744 8084 22784
rect 8140 23120 8180 23129
rect 7659 21944 7701 21953
rect 7659 21904 7660 21944
rect 7700 21904 7701 21944
rect 7659 21895 7701 21904
rect 7371 21860 7413 21869
rect 7371 21820 7372 21860
rect 7412 21820 7413 21860
rect 7371 21811 7413 21820
rect 7563 21860 7605 21869
rect 7563 21820 7564 21860
rect 7604 21820 7605 21860
rect 7563 21811 7605 21820
rect 7468 21617 7508 21702
rect 7564 21692 7604 21811
rect 7564 21643 7604 21652
rect 7467 21608 7509 21617
rect 7467 21568 7468 21608
rect 7508 21568 7509 21608
rect 7467 21559 7509 21568
rect 7276 21484 7412 21524
rect 7084 21400 7316 21440
rect 6987 21391 7029 21400
rect 6892 21232 7124 21272
rect 6892 21020 6932 21029
rect 6796 20980 6892 21020
rect 6892 20971 6932 20980
rect 6700 19349 6740 20728
rect 7084 20768 7124 21232
rect 7084 20719 7124 20728
rect 6892 20600 6932 20609
rect 6932 20560 7220 20600
rect 6892 20551 6932 20560
rect 7180 20096 7220 20560
rect 7276 20180 7316 21400
rect 7372 20189 7412 21484
rect 7467 21440 7509 21449
rect 7467 21400 7468 21440
rect 7508 21400 7509 21440
rect 7467 21391 7509 21400
rect 7276 20131 7316 20140
rect 7371 20180 7413 20189
rect 7371 20140 7372 20180
rect 7412 20140 7413 20180
rect 7371 20131 7413 20140
rect 7180 20047 7220 20056
rect 6699 19340 6741 19349
rect 6699 19300 6700 19340
rect 6740 19300 6741 19340
rect 6699 19291 6741 19300
rect 6796 19256 6836 19267
rect 6796 19181 6836 19216
rect 6795 19172 6837 19181
rect 6795 19132 6796 19172
rect 6836 19132 6837 19172
rect 6795 19123 6837 19132
rect 7275 19088 7317 19097
rect 7275 19048 7276 19088
rect 7316 19048 7317 19088
rect 7275 19039 7317 19048
rect 6604 18880 6740 18920
rect 6316 18796 6644 18836
rect 5932 18712 6068 18752
rect 5835 18668 5877 18677
rect 5835 18628 5836 18668
rect 5876 18628 5877 18668
rect 5835 18619 5877 18628
rect 5836 18584 5876 18619
rect 5836 18533 5876 18544
rect 5932 18584 5972 18595
rect 6028 18584 6068 18712
rect 6124 18703 6164 18712
rect 6219 18752 6261 18761
rect 6219 18712 6220 18752
rect 6260 18712 6261 18752
rect 6219 18703 6261 18712
rect 6028 18544 6164 18584
rect 5932 18509 5972 18544
rect 5931 18500 5973 18509
rect 5931 18460 5932 18500
rect 5972 18460 5973 18500
rect 5931 18451 5973 18460
rect 5835 18164 5877 18173
rect 5835 18124 5836 18164
rect 5876 18124 5877 18164
rect 5835 18115 5877 18124
rect 5836 17921 5876 18115
rect 5835 17912 5877 17921
rect 5835 17872 5836 17912
rect 5876 17872 5877 17912
rect 5835 17863 5877 17872
rect 5836 17072 5876 17863
rect 6027 17576 6069 17585
rect 6027 17536 6028 17576
rect 6068 17536 6069 17576
rect 6027 17527 6069 17536
rect 5836 17023 5876 17032
rect 6028 15905 6068 17527
rect 6027 15896 6069 15905
rect 6027 15856 6028 15896
rect 6068 15856 6069 15896
rect 6027 15847 6069 15856
rect 5835 15476 5877 15485
rect 5740 15436 5836 15476
rect 5876 15436 5877 15476
rect 5643 15427 5685 15436
rect 5835 15427 5877 15436
rect 5931 15056 5973 15065
rect 5931 15016 5932 15056
rect 5972 15016 5973 15056
rect 5931 15007 5973 15016
rect 5452 14923 5492 14932
rect 5259 14720 5301 14729
rect 5259 14680 5260 14720
rect 5300 14680 5301 14720
rect 5259 14671 5301 14680
rect 5644 14720 5684 14729
rect 5260 14561 5300 14671
rect 5259 14552 5301 14561
rect 5259 14512 5260 14552
rect 5300 14512 5301 14552
rect 5259 14503 5301 14512
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 5163 14216 5205 14225
rect 5163 14176 5164 14216
rect 5204 14176 5205 14216
rect 5163 14167 5205 14176
rect 5356 14216 5396 14225
rect 5396 14176 5588 14216
rect 5356 14167 5396 14176
rect 4876 14048 4916 14057
rect 4436 14008 4532 14048
rect 4396 13999 4436 14008
rect 4011 13964 4053 13973
rect 4011 13924 4012 13964
rect 4052 13924 4053 13964
rect 4011 13915 4053 13924
rect 4108 13964 4148 13975
rect 4108 13889 4148 13924
rect 4299 13964 4341 13973
rect 4299 13924 4300 13964
rect 4340 13924 4341 13964
rect 4299 13915 4341 13924
rect 4107 13880 4149 13889
rect 4107 13840 4108 13880
rect 4148 13840 4149 13880
rect 4107 13831 4149 13840
rect 4204 13880 4244 13889
rect 3532 13756 3764 13796
rect 3532 13208 3572 13756
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 3628 13376 3668 13385
rect 3668 13336 3764 13376
rect 3628 13327 3668 13336
rect 3532 13168 3668 13208
rect 3339 12704 3381 12713
rect 3339 12664 3340 12704
rect 3380 12664 3381 12704
rect 3339 12655 3381 12664
rect 3532 12545 3572 12630
rect 3628 12620 3668 13168
rect 3628 12571 3668 12580
rect 3339 12536 3381 12545
rect 3339 12496 3340 12536
rect 3380 12496 3381 12536
rect 3339 12487 3381 12496
rect 3436 12536 3476 12545
rect 3340 12402 3380 12487
rect 3436 12377 3476 12496
rect 3531 12536 3573 12545
rect 3531 12496 3532 12536
rect 3572 12496 3573 12536
rect 3531 12487 3573 12496
rect 3435 12368 3477 12377
rect 3724 12368 3764 13336
rect 4011 13292 4053 13301
rect 4011 13252 4012 13292
rect 4052 13252 4053 13292
rect 4011 13243 4053 13252
rect 3915 13208 3957 13217
rect 3915 13168 3916 13208
rect 3956 13168 3957 13208
rect 3915 13159 3957 13168
rect 4012 13208 4052 13243
rect 3916 13074 3956 13159
rect 4012 13157 4052 13168
rect 4107 13040 4149 13049
rect 4107 13000 4108 13040
rect 4148 13000 4149 13040
rect 4107 12991 4149 13000
rect 3915 12620 3957 12629
rect 3915 12580 3916 12620
rect 3956 12580 3957 12620
rect 3915 12571 3957 12580
rect 3819 12536 3861 12545
rect 3819 12496 3820 12536
rect 3860 12496 3861 12536
rect 3819 12487 3861 12496
rect 3916 12536 3956 12571
rect 3820 12402 3860 12487
rect 3916 12485 3956 12496
rect 4011 12536 4053 12545
rect 4011 12496 4012 12536
rect 4052 12496 4053 12536
rect 4011 12487 4053 12496
rect 4108 12536 4148 12991
rect 4108 12487 4148 12496
rect 4012 12402 4052 12487
rect 3435 12328 3436 12368
rect 3476 12328 3477 12368
rect 3435 12319 3477 12328
rect 3532 12328 3764 12368
rect 3339 12284 3381 12293
rect 3339 12244 3340 12284
rect 3380 12244 3381 12284
rect 3339 12235 3381 12244
rect 3243 11696 3285 11705
rect 3243 11656 3244 11696
rect 3284 11656 3285 11696
rect 3243 11647 3285 11656
rect 3340 11696 3380 12235
rect 3436 11873 3476 11958
rect 3435 11864 3477 11873
rect 3435 11824 3436 11864
rect 3476 11824 3477 11864
rect 3435 11815 3477 11824
rect 3532 11696 3572 12328
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 3724 11873 3764 11958
rect 3915 11948 3957 11957
rect 3915 11908 3916 11948
rect 3956 11908 3957 11948
rect 3915 11899 3957 11908
rect 3723 11864 3765 11873
rect 3723 11824 3724 11864
rect 3764 11824 3765 11864
rect 3723 11815 3765 11824
rect 3628 11696 3668 11705
rect 3380 11656 3476 11696
rect 3532 11656 3628 11696
rect 3340 11647 3380 11656
rect 3339 11528 3381 11537
rect 3339 11488 3340 11528
rect 3380 11488 3381 11528
rect 3436 11528 3476 11656
rect 3628 11647 3668 11656
rect 3724 11696 3764 11705
rect 3724 11528 3764 11656
rect 3916 11696 3956 11899
rect 3916 11647 3956 11656
rect 4107 11696 4149 11705
rect 4107 11656 4108 11696
rect 4148 11656 4149 11696
rect 4107 11647 4149 11656
rect 4204 11696 4244 13840
rect 4300 13830 4340 13915
rect 4300 13208 4340 13217
rect 4300 12713 4340 13168
rect 4299 12704 4341 12713
rect 4299 12664 4300 12704
rect 4340 12664 4341 12704
rect 4299 12655 4341 12664
rect 4300 12452 4340 12655
rect 4395 12452 4437 12461
rect 4300 12412 4396 12452
rect 4436 12412 4437 12452
rect 4395 12403 4437 12412
rect 4299 12116 4341 12125
rect 4299 12076 4300 12116
rect 4340 12076 4341 12116
rect 4299 12067 4341 12076
rect 4300 11864 4340 12067
rect 4300 11815 4340 11824
rect 4204 11647 4244 11656
rect 4396 11696 4436 12403
rect 4492 11789 4532 14008
rect 4588 14008 4724 14048
rect 4780 14008 4876 14048
rect 4588 13217 4628 14008
rect 4684 13880 4724 13889
rect 4684 13721 4724 13840
rect 4683 13712 4725 13721
rect 4683 13672 4684 13712
rect 4724 13672 4725 13712
rect 4683 13663 4725 13672
rect 4684 13376 4724 13663
rect 4587 13208 4629 13217
rect 4587 13168 4588 13208
rect 4628 13168 4629 13208
rect 4587 13159 4629 13168
rect 4684 12629 4724 13336
rect 4683 12620 4725 12629
rect 4683 12580 4684 12620
rect 4724 12580 4725 12620
rect 4683 12571 4725 12580
rect 4587 12368 4629 12377
rect 4587 12328 4588 12368
rect 4628 12328 4629 12368
rect 4587 12319 4629 12328
rect 4588 12234 4628 12319
rect 4684 11864 4724 12571
rect 4780 11873 4820 14008
rect 4876 13999 4916 14008
rect 4972 14048 5012 14057
rect 4972 13805 5012 14008
rect 5164 14048 5204 14167
rect 5251 14132 5293 14141
rect 5251 14092 5252 14132
rect 5292 14092 5300 14132
rect 5251 14083 5300 14092
rect 5164 13999 5204 14008
rect 5260 14048 5300 14083
rect 5260 13999 5300 14008
rect 5417 14033 5457 14042
rect 4971 13796 5013 13805
rect 4971 13756 4972 13796
rect 5012 13756 5013 13796
rect 4971 13747 5013 13756
rect 5163 13628 5205 13637
rect 5163 13588 5164 13628
rect 5204 13588 5205 13628
rect 5417 13628 5457 13993
rect 5417 13588 5492 13628
rect 5163 13579 5205 13588
rect 5164 13208 5204 13579
rect 5164 13159 5204 13168
rect 5260 13208 5300 13217
rect 5300 13168 5396 13208
rect 5260 13159 5300 13168
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 4875 12620 4917 12629
rect 4875 12580 4876 12620
rect 4916 12580 4917 12620
rect 4875 12571 4917 12580
rect 5259 12620 5301 12629
rect 5259 12580 5260 12620
rect 5300 12580 5301 12620
rect 5259 12571 5301 12580
rect 4876 12486 4916 12571
rect 4972 12536 5012 12547
rect 4972 12461 5012 12496
rect 5260 12536 5300 12571
rect 4971 12452 5013 12461
rect 4971 12412 4972 12452
rect 5012 12412 5013 12452
rect 4971 12403 5013 12412
rect 5260 12293 5300 12496
rect 5259 12284 5301 12293
rect 5259 12244 5260 12284
rect 5300 12244 5301 12284
rect 5259 12235 5301 12244
rect 4491 11780 4533 11789
rect 4491 11740 4492 11780
rect 4532 11740 4533 11780
rect 4491 11731 4533 11740
rect 4684 11705 4724 11824
rect 4779 11864 4821 11873
rect 4779 11824 4780 11864
rect 4820 11824 4821 11864
rect 4779 11815 4821 11824
rect 4971 11864 5013 11873
rect 4971 11824 4972 11864
rect 5012 11824 5013 11864
rect 4971 11815 5013 11824
rect 4396 11647 4436 11656
rect 4683 11696 4725 11705
rect 4683 11656 4684 11696
rect 4724 11656 4725 11696
rect 4683 11647 4725 11656
rect 4972 11696 5012 11815
rect 4972 11647 5012 11656
rect 4108 11562 4148 11647
rect 3436 11488 3764 11528
rect 4491 11528 4533 11537
rect 4491 11488 4492 11528
rect 4532 11488 4533 11528
rect 3339 11479 3381 11488
rect 4491 11479 4533 11488
rect 3148 10184 3188 10193
rect 3052 10144 3148 10184
rect 2763 10100 2805 10109
rect 2763 10060 2764 10100
rect 2804 10060 2805 10100
rect 2763 10051 2805 10060
rect 2955 10100 2997 10109
rect 2955 10060 2956 10100
rect 2996 10060 2997 10100
rect 2955 10051 2997 10060
rect 2764 9512 2804 10051
rect 2956 9966 2996 10051
rect 3052 9680 3092 10144
rect 3148 10135 3188 10144
rect 3052 9631 3092 9640
rect 2860 9521 2900 9606
rect 2859 9512 2901 9521
rect 2764 9472 2860 9512
rect 2900 9472 2901 9512
rect 2859 9463 2901 9472
rect 3243 9512 3285 9521
rect 3243 9472 3244 9512
rect 3284 9472 3285 9512
rect 3243 9463 3285 9472
rect 2859 9344 2901 9353
rect 2859 9304 2860 9344
rect 2900 9304 2901 9344
rect 2859 9295 2901 9304
rect 2571 7832 2613 7841
rect 2571 7792 2572 7832
rect 2612 7792 2613 7832
rect 2571 7783 2613 7792
rect 2860 7748 2900 9295
rect 3052 9260 3092 9269
rect 2956 9220 3052 9260
rect 2956 8429 2996 9220
rect 3052 9211 3092 9220
rect 3148 8672 3188 8700
rect 3244 8672 3284 9463
rect 3340 9092 3380 11479
rect 3435 11360 3477 11369
rect 4492 11360 4532 11479
rect 3435 11320 3436 11360
rect 3476 11320 3477 11360
rect 3435 11311 3477 11320
rect 4396 11320 4532 11360
rect 3436 10436 3476 11311
rect 3723 11276 3765 11285
rect 3723 11236 3724 11276
rect 3764 11236 3765 11276
rect 3723 11227 3765 11236
rect 3531 11108 3573 11117
rect 3531 11068 3532 11108
rect 3572 11068 3573 11108
rect 3531 11059 3573 11068
rect 3436 10387 3476 10396
rect 3435 10184 3477 10193
rect 3435 10144 3436 10184
rect 3476 10144 3477 10184
rect 3435 10135 3477 10144
rect 3436 10050 3476 10135
rect 3532 9932 3572 11059
rect 3724 10865 3764 11227
rect 4203 11192 4245 11201
rect 4203 11152 4204 11192
rect 4244 11152 4245 11192
rect 4203 11143 4245 11152
rect 4107 11024 4149 11033
rect 4107 10984 4108 11024
rect 4148 10984 4149 11024
rect 4107 10975 4149 10984
rect 4108 10890 4148 10975
rect 3723 10856 3765 10865
rect 3723 10816 3724 10856
rect 3764 10816 3765 10856
rect 3723 10807 3765 10816
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 3819 10352 3861 10361
rect 3819 10312 3820 10352
rect 3860 10312 3861 10352
rect 3819 10303 3861 10312
rect 3724 10268 3764 10277
rect 3628 10184 3668 10195
rect 3628 10109 3668 10144
rect 3627 10100 3669 10109
rect 3627 10060 3628 10100
rect 3668 10060 3669 10100
rect 3627 10051 3669 10060
rect 3436 9892 3572 9932
rect 3436 9521 3476 9892
rect 3724 9680 3764 10228
rect 3820 10218 3860 10303
rect 3916 10268 3956 10277
rect 3916 10025 3956 10228
rect 4012 10184 4052 10193
rect 4204 10184 4244 11143
rect 4299 10772 4341 10781
rect 4299 10732 4300 10772
rect 4340 10732 4341 10772
rect 4299 10723 4341 10732
rect 4300 10638 4340 10723
rect 3915 10016 3957 10025
rect 3915 9976 3916 10016
rect 3956 9976 3957 10016
rect 3915 9967 3957 9976
rect 4012 9764 4052 10144
rect 3532 9640 3764 9680
rect 3916 9724 4052 9764
rect 4108 10144 4204 10184
rect 3435 9512 3477 9521
rect 3435 9472 3436 9512
rect 3476 9472 3477 9512
rect 3435 9463 3477 9472
rect 3436 9269 3476 9463
rect 3532 9344 3572 9640
rect 3916 9605 3956 9724
rect 3915 9596 3957 9605
rect 3915 9556 3916 9596
rect 3956 9556 3957 9596
rect 3915 9547 3957 9556
rect 3627 9512 3669 9521
rect 3716 9512 3756 9520
rect 3627 9472 3628 9512
rect 3668 9511 3756 9512
rect 3668 9472 3716 9511
rect 3627 9463 3669 9472
rect 3716 9462 3756 9471
rect 4012 9512 4052 9521
rect 4108 9512 4148 10144
rect 4204 10135 4244 10144
rect 4396 10184 4436 11320
rect 4684 11192 4724 11647
rect 4928 11360 5296 11369
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 4684 11143 4724 11152
rect 5356 11033 5396 13168
rect 5452 12377 5492 13588
rect 5548 12545 5588 14176
rect 5644 13973 5684 14680
rect 5836 14720 5876 14729
rect 5740 14552 5780 14561
rect 5740 14057 5780 14512
rect 5836 14393 5876 14680
rect 5932 14720 5972 15007
rect 6028 14729 6068 15847
rect 5932 14671 5972 14680
rect 6027 14720 6069 14729
rect 6027 14680 6028 14720
rect 6068 14680 6069 14720
rect 6027 14671 6069 14680
rect 6124 14552 6164 18544
rect 6220 18173 6260 18703
rect 6316 18584 6356 18593
rect 6219 18164 6261 18173
rect 6219 18124 6220 18164
rect 6260 18124 6261 18164
rect 6219 18115 6261 18124
rect 6316 17837 6356 18544
rect 6411 18584 6453 18593
rect 6501 18584 6541 18592
rect 6411 18544 6412 18584
rect 6452 18583 6541 18584
rect 6452 18544 6501 18583
rect 6411 18535 6453 18544
rect 6501 18534 6541 18543
rect 6604 18416 6644 18796
rect 6700 18761 6740 18880
rect 6699 18752 6741 18761
rect 6699 18712 6700 18752
rect 6740 18712 6741 18752
rect 6699 18703 6741 18712
rect 6795 18584 6837 18593
rect 6795 18544 6796 18584
rect 6836 18544 6837 18584
rect 6795 18535 6837 18544
rect 6987 18584 7029 18593
rect 6987 18544 6988 18584
rect 7028 18544 7029 18584
rect 6987 18535 7029 18544
rect 6796 18416 6836 18535
rect 6508 18376 6644 18416
rect 6700 18376 6836 18416
rect 6411 18332 6453 18341
rect 6411 18292 6412 18332
rect 6452 18292 6453 18332
rect 6411 18283 6453 18292
rect 6412 18198 6452 18283
rect 6411 17996 6453 18005
rect 6411 17956 6412 17996
rect 6452 17956 6453 17996
rect 6411 17947 6453 17956
rect 6315 17828 6357 17837
rect 6315 17788 6316 17828
rect 6356 17788 6357 17828
rect 6315 17779 6357 17788
rect 5932 14512 6164 14552
rect 5835 14384 5877 14393
rect 5835 14344 5836 14384
rect 5876 14344 5877 14384
rect 5835 14335 5877 14344
rect 5836 14216 5876 14225
rect 5739 14048 5781 14057
rect 5739 14008 5740 14048
rect 5780 14008 5781 14048
rect 5739 13999 5781 14008
rect 5643 13964 5685 13973
rect 5643 13924 5644 13964
rect 5684 13924 5685 13964
rect 5643 13915 5685 13924
rect 5836 13889 5876 14176
rect 5835 13880 5877 13889
rect 5835 13840 5836 13880
rect 5876 13840 5877 13880
rect 5835 13831 5877 13840
rect 5643 13208 5685 13217
rect 5643 13168 5644 13208
rect 5684 13168 5685 13208
rect 5643 13159 5685 13168
rect 5740 13208 5780 13217
rect 5780 13168 5876 13208
rect 5740 13159 5780 13168
rect 5644 13074 5684 13159
rect 5643 12872 5685 12881
rect 5643 12832 5644 12872
rect 5684 12832 5685 12872
rect 5643 12823 5685 12832
rect 5644 12713 5684 12823
rect 5643 12704 5685 12713
rect 5643 12664 5644 12704
rect 5684 12664 5685 12704
rect 5643 12655 5685 12664
rect 5547 12536 5589 12545
rect 5547 12496 5548 12536
rect 5588 12496 5589 12536
rect 5547 12487 5589 12496
rect 5644 12536 5684 12655
rect 5644 12487 5684 12496
rect 5739 12536 5781 12545
rect 5739 12496 5740 12536
rect 5780 12496 5781 12536
rect 5739 12487 5781 12496
rect 5740 12402 5780 12487
rect 5451 12368 5493 12377
rect 5451 12328 5452 12368
rect 5492 12328 5493 12368
rect 5451 12319 5493 12328
rect 5451 11192 5493 11201
rect 5451 11152 5452 11192
rect 5492 11152 5493 11192
rect 5451 11143 5493 11152
rect 5163 11024 5205 11033
rect 5163 10984 5164 11024
rect 5204 10984 5205 11024
rect 5163 10975 5205 10984
rect 5355 11024 5397 11033
rect 5355 10984 5356 11024
rect 5396 10984 5397 11024
rect 5355 10975 5397 10984
rect 5452 11024 5492 11143
rect 5644 11024 5684 11033
rect 5452 10975 5492 10984
rect 5548 10984 5644 11024
rect 5164 10890 5204 10975
rect 4779 10772 4821 10781
rect 4779 10732 4780 10772
rect 4820 10732 4821 10772
rect 4779 10723 4821 10732
rect 4588 10352 4628 10361
rect 4396 10135 4436 10144
rect 4492 10312 4588 10352
rect 4300 10100 4340 10109
rect 4300 9680 4340 10060
rect 4052 9472 4148 9512
rect 4012 9463 4052 9472
rect 3628 9344 3668 9353
rect 3532 9304 3579 9344
rect 3435 9260 3477 9269
rect 3435 9220 3436 9260
rect 3476 9220 3477 9260
rect 3435 9211 3477 9220
rect 3340 9052 3476 9092
rect 3340 8840 3380 8849
rect 3340 8681 3380 8800
rect 3188 8632 3284 8672
rect 3148 8623 3188 8632
rect 3051 8588 3093 8597
rect 3051 8548 3052 8588
rect 3092 8548 3093 8588
rect 3051 8539 3093 8548
rect 2955 8420 2997 8429
rect 2955 8380 2956 8420
rect 2996 8380 2997 8420
rect 2955 8371 2997 8380
rect 2955 8000 2997 8009
rect 2955 7960 2956 8000
rect 2996 7960 2997 8000
rect 2955 7951 2997 7960
rect 3052 8000 3092 8539
rect 3244 8504 3284 8632
rect 3339 8672 3381 8681
rect 3339 8632 3340 8672
rect 3380 8632 3381 8672
rect 3339 8623 3381 8632
rect 3244 8464 3380 8504
rect 3147 8420 3189 8429
rect 3147 8380 3148 8420
rect 3188 8380 3189 8420
rect 3147 8371 3189 8380
rect 3052 7951 3092 7960
rect 3148 8000 3188 8371
rect 3243 8336 3285 8345
rect 3243 8296 3244 8336
rect 3284 8296 3285 8336
rect 3243 8287 3285 8296
rect 3148 7951 3188 7960
rect 3244 8000 3284 8287
rect 3244 7951 3284 7960
rect 2956 7866 2996 7951
rect 2860 7708 3284 7748
rect 2284 6280 2420 6320
rect 2380 80 2420 6280
rect 3147 3716 3189 3725
rect 3147 3676 3148 3716
rect 3188 3676 3189 3716
rect 3147 3667 3189 3676
rect 2955 1280 2997 1289
rect 2955 1240 2956 1280
rect 2996 1240 2997 1280
rect 2955 1231 2997 1240
rect 2571 944 2613 953
rect 2571 904 2572 944
rect 2612 904 2613 944
rect 2571 895 2613 904
rect 2572 80 2612 895
rect 2763 608 2805 617
rect 2763 568 2764 608
rect 2804 568 2805 608
rect 2763 559 2805 568
rect 2764 80 2804 559
rect 2956 80 2996 1231
rect 3148 80 3188 3667
rect 3244 1196 3284 7708
rect 3340 3221 3380 8464
rect 3436 8000 3476 9052
rect 3539 8840 3579 9304
rect 3628 9269 3668 9304
rect 3628 9260 3676 9269
rect 3628 9220 3635 9260
rect 3675 9220 3676 9260
rect 3634 9211 3676 9220
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3627 8924 3669 8933
rect 3627 8884 3628 8924
rect 3668 8884 3669 8924
rect 3627 8875 3669 8884
rect 3915 8924 3957 8933
rect 3915 8884 3916 8924
rect 3956 8884 3957 8924
rect 3915 8875 3957 8884
rect 3532 8800 3579 8840
rect 3532 8177 3572 8800
rect 3628 8345 3668 8875
rect 3723 8840 3765 8849
rect 3826 8840 3868 8849
rect 3723 8800 3724 8840
rect 3764 8800 3765 8840
rect 3723 8791 3765 8800
rect 3820 8800 3827 8840
rect 3867 8800 3868 8840
rect 3820 8791 3868 8800
rect 3627 8336 3669 8345
rect 3627 8296 3628 8336
rect 3668 8296 3669 8336
rect 3627 8287 3669 8296
rect 3531 8168 3573 8177
rect 3531 8128 3532 8168
rect 3572 8128 3573 8168
rect 3531 8119 3573 8128
rect 3628 8168 3668 8177
rect 3724 8168 3764 8791
rect 3668 8128 3764 8168
rect 3628 8119 3668 8128
rect 3820 8084 3860 8791
rect 3916 8790 3956 8875
rect 4108 8840 4148 9472
rect 4012 8800 4148 8840
rect 4204 9640 4340 9680
rect 3916 8672 3956 8683
rect 4012 8681 4052 8800
rect 3916 8597 3956 8632
rect 4011 8672 4053 8681
rect 4011 8632 4012 8672
rect 4052 8632 4053 8672
rect 4011 8623 4053 8632
rect 4108 8672 4148 8681
rect 3915 8588 3957 8597
rect 3915 8548 3916 8588
rect 3956 8548 3957 8588
rect 3915 8539 3957 8548
rect 3916 8177 3956 8262
rect 3915 8168 3957 8177
rect 3915 8128 3916 8168
rect 3956 8128 3957 8168
rect 3915 8119 3957 8128
rect 3724 8044 3860 8084
rect 3436 7951 3476 7960
rect 3531 8000 3573 8009
rect 3531 7960 3532 8000
rect 3572 7960 3573 8000
rect 3531 7951 3573 7960
rect 3724 8000 3764 8044
rect 3724 7951 3764 7960
rect 3916 8000 3956 8009
rect 4012 8000 4052 8623
rect 4108 8345 4148 8632
rect 4204 8672 4244 9640
rect 4300 9512 4340 9521
rect 4300 9353 4340 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4299 9344 4341 9353
rect 4299 9304 4300 9344
rect 4340 9304 4341 9344
rect 4299 9295 4341 9304
rect 4396 9008 4436 9463
rect 4492 9269 4532 10312
rect 4588 10303 4628 10312
rect 4588 10184 4628 10193
rect 4491 9260 4533 9269
rect 4491 9220 4492 9260
rect 4532 9220 4533 9260
rect 4491 9211 4533 9220
rect 4204 8623 4244 8632
rect 4300 8968 4436 9008
rect 4491 9008 4533 9017
rect 4491 8968 4492 9008
rect 4532 8968 4533 9008
rect 4203 8504 4245 8513
rect 4203 8464 4204 8504
rect 4244 8464 4245 8504
rect 4203 8455 4245 8464
rect 4107 8336 4149 8345
rect 4107 8296 4108 8336
rect 4148 8296 4149 8336
rect 4107 8287 4149 8296
rect 4107 8168 4149 8177
rect 4107 8128 4108 8168
rect 4148 8128 4149 8168
rect 4107 8119 4149 8128
rect 3956 7960 4052 8000
rect 4108 8000 4148 8119
rect 3916 7951 3956 7960
rect 4108 7951 4148 7960
rect 4204 8000 4244 8455
rect 4204 7951 4244 7960
rect 3532 7866 3572 7951
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 4203 7580 4245 7589
rect 4203 7540 4204 7580
rect 4244 7540 4245 7580
rect 4203 7531 4245 7540
rect 4204 7160 4244 7531
rect 4204 7111 4244 7120
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 3339 3212 3381 3221
rect 3339 3172 3340 3212
rect 3380 3172 3381 3212
rect 3339 3163 3381 3172
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4300 2540 4340 8968
rect 4491 8959 4533 8968
rect 4492 8756 4532 8959
rect 4492 8707 4532 8716
rect 4395 8672 4437 8681
rect 4395 8632 4396 8672
rect 4436 8632 4437 8672
rect 4395 8623 4437 8632
rect 4396 8538 4436 8623
rect 4491 8420 4533 8429
rect 4491 8380 4492 8420
rect 4532 8380 4533 8420
rect 4491 8371 4533 8380
rect 4492 7664 4532 8371
rect 4588 7832 4628 10144
rect 4780 10184 4820 10723
rect 5356 10613 5396 10975
rect 5452 10856 5492 10865
rect 5548 10856 5588 10984
rect 5644 10975 5684 10984
rect 5739 11024 5781 11033
rect 5739 10984 5740 11024
rect 5780 10984 5781 11024
rect 5739 10975 5781 10984
rect 5836 11024 5876 13168
rect 5932 12713 5972 14512
rect 6027 14384 6069 14393
rect 6027 14344 6028 14384
rect 6068 14344 6069 14384
rect 6027 14335 6069 14344
rect 6028 14048 6068 14335
rect 6412 14309 6452 17947
rect 6123 14300 6165 14309
rect 6123 14260 6124 14300
rect 6164 14260 6165 14300
rect 6123 14251 6165 14260
rect 6411 14300 6453 14309
rect 6411 14260 6412 14300
rect 6452 14260 6453 14300
rect 6411 14251 6453 14260
rect 6124 14057 6164 14251
rect 6023 14008 6028 14033
rect 6023 13993 6068 14008
rect 6123 14048 6165 14057
rect 6123 14008 6124 14048
rect 6164 14008 6165 14048
rect 6123 13999 6165 14008
rect 6412 14048 6452 14057
rect 6023 13880 6063 13993
rect 6315 13964 6357 13973
rect 6315 13924 6316 13964
rect 6356 13924 6357 13964
rect 6315 13915 6357 13924
rect 6023 13840 6068 13880
rect 6028 13637 6068 13840
rect 6316 13830 6356 13915
rect 6412 13805 6452 14008
rect 6411 13796 6453 13805
rect 6411 13756 6412 13796
rect 6452 13756 6453 13796
rect 6411 13747 6453 13756
rect 6027 13628 6069 13637
rect 6027 13588 6028 13628
rect 6068 13588 6069 13628
rect 6027 13579 6069 13588
rect 6123 13544 6165 13553
rect 6123 13504 6124 13544
rect 6164 13504 6165 13544
rect 6123 13495 6165 13504
rect 6124 12881 6164 13495
rect 6220 13208 6260 13217
rect 6123 12872 6165 12881
rect 6123 12832 6124 12872
rect 6164 12832 6165 12872
rect 6123 12823 6165 12832
rect 5931 12704 5973 12713
rect 5931 12664 5932 12704
rect 5972 12664 5973 12704
rect 5931 12655 5973 12664
rect 5932 12536 5972 12545
rect 6124 12536 6164 12823
rect 5972 12496 6068 12536
rect 5932 12487 5972 12496
rect 5931 12368 5973 12377
rect 5931 12328 5932 12368
rect 5972 12328 5973 12368
rect 5931 12319 5973 12328
rect 5932 12234 5972 12319
rect 6028 12284 6068 12496
rect 6124 12487 6164 12496
rect 6124 12284 6164 12293
rect 6028 12244 6124 12284
rect 6124 12235 6164 12244
rect 6220 12116 6260 13168
rect 6412 12881 6452 13747
rect 6508 13217 6548 18376
rect 6603 18164 6645 18173
rect 6603 18124 6604 18164
rect 6644 18124 6645 18164
rect 6603 18115 6645 18124
rect 6604 17744 6644 18115
rect 6604 17585 6644 17704
rect 6603 17576 6645 17585
rect 6603 17536 6604 17576
rect 6644 17536 6645 17576
rect 6603 17527 6645 17536
rect 6700 16064 6740 18376
rect 6891 17744 6933 17753
rect 6796 17704 6892 17744
rect 6932 17704 6933 17744
rect 6796 17660 6836 17704
rect 6891 17695 6933 17704
rect 6796 17611 6836 17620
rect 6988 17576 7028 18535
rect 7084 17753 7124 17838
rect 7083 17744 7125 17753
rect 7083 17704 7084 17744
rect 7124 17704 7125 17744
rect 7083 17695 7125 17704
rect 7180 17744 7220 17753
rect 7180 17585 7220 17704
rect 6892 17536 7028 17576
rect 7179 17576 7221 17585
rect 7179 17536 7180 17576
rect 7220 17536 7221 17576
rect 6892 16745 6932 17536
rect 7179 17527 7221 17536
rect 7276 17408 7316 19039
rect 7084 17368 7316 17408
rect 7084 17072 7124 17368
rect 7372 17324 7412 20131
rect 7468 17417 7508 21391
rect 7563 21356 7605 21365
rect 7563 21316 7564 21356
rect 7604 21316 7605 21356
rect 7563 21307 7605 21316
rect 7564 19097 7604 21307
rect 7563 19088 7605 19097
rect 7563 19048 7564 19088
rect 7604 19048 7605 19088
rect 7563 19039 7605 19048
rect 7563 18752 7605 18761
rect 7563 18712 7564 18752
rect 7604 18712 7605 18752
rect 7563 18703 7605 18712
rect 7564 18248 7604 18703
rect 7660 18425 7700 21895
rect 7659 18416 7701 18425
rect 7659 18376 7660 18416
rect 7700 18376 7701 18416
rect 7659 18367 7701 18376
rect 7564 18208 7700 18248
rect 7564 17744 7604 17753
rect 7564 17585 7604 17704
rect 7660 17744 7700 18208
rect 7756 17921 7796 22744
rect 8140 22448 8180 23080
rect 7948 22408 8180 22448
rect 8236 23120 8276 23129
rect 7851 22280 7893 22289
rect 7851 22240 7852 22280
rect 7892 22240 7893 22280
rect 7851 22231 7893 22240
rect 7948 22280 7988 22408
rect 7852 22146 7892 22231
rect 7948 21785 7988 22240
rect 8140 22280 8180 22289
rect 8140 22121 8180 22240
rect 8139 22112 8181 22121
rect 8139 22072 8140 22112
rect 8180 22072 8181 22112
rect 8139 22063 8181 22072
rect 7947 21776 7989 21785
rect 7947 21736 7948 21776
rect 7988 21736 7989 21776
rect 7947 21727 7989 21736
rect 8044 21617 8084 21702
rect 8043 21608 8085 21617
rect 8043 21568 8044 21608
rect 8084 21568 8085 21608
rect 8043 21559 8085 21568
rect 7852 21440 7892 21449
rect 8236 21440 8276 23080
rect 8332 21953 8372 24424
rect 8524 23129 8564 24508
rect 8620 24389 8660 30043
rect 8716 29849 8756 30640
rect 8715 29840 8757 29849
rect 8715 29800 8716 29840
rect 8756 29800 8757 29840
rect 8715 29791 8757 29800
rect 8716 29672 8756 29681
rect 8716 29163 8756 29632
rect 8716 29114 8756 29123
rect 8715 27404 8757 27413
rect 8715 27364 8716 27404
rect 8756 27364 8757 27404
rect 8715 27355 8757 27364
rect 8716 26144 8756 27355
rect 8812 26816 8852 31471
rect 9004 31445 9044 32740
rect 9196 32696 9236 32705
rect 9196 31445 9236 32656
rect 9003 31436 9045 31445
rect 9003 31396 9004 31436
rect 9044 31396 9045 31436
rect 9003 31387 9045 31396
rect 9195 31436 9237 31445
rect 9195 31396 9196 31436
rect 9236 31396 9237 31436
rect 9195 31387 9237 31396
rect 8908 31352 8948 31361
rect 8908 30269 8948 31312
rect 9195 31184 9237 31193
rect 9195 31144 9196 31184
rect 9236 31144 9237 31184
rect 9195 31135 9237 31144
rect 9196 30675 9236 31135
rect 9196 30626 9236 30635
rect 8907 30260 8949 30269
rect 8907 30220 8908 30260
rect 8948 30220 8949 30260
rect 8907 30211 8949 30220
rect 8908 30017 8948 30211
rect 8907 30008 8949 30017
rect 8907 29968 8908 30008
rect 8948 29968 8949 30008
rect 8907 29959 8949 29968
rect 9099 29840 9141 29849
rect 9099 29800 9100 29840
rect 9140 29800 9141 29840
rect 9099 29791 9141 29800
rect 9100 29706 9140 29791
rect 8908 29252 8948 29261
rect 8908 28589 8948 29212
rect 9292 29000 9332 37780
rect 9388 37409 9428 37494
rect 9387 37400 9429 37409
rect 9387 37360 9388 37400
rect 9428 37360 9429 37400
rect 9387 37351 9429 37360
rect 9580 37400 9620 37409
rect 9388 37232 9428 37241
rect 9428 37192 9524 37232
rect 9388 37183 9428 37192
rect 9387 36560 9429 36569
rect 9387 36520 9388 36560
rect 9428 36520 9429 36560
rect 9387 36511 9429 36520
rect 9388 35888 9428 36511
rect 9388 35839 9428 35848
rect 9388 35216 9428 35225
rect 9388 34469 9428 35176
rect 9484 35132 9524 37192
rect 9580 36896 9620 37360
rect 9676 37400 9716 37780
rect 9676 37351 9716 37360
rect 9580 36847 9620 36856
rect 9771 36728 9813 36737
rect 9771 36688 9772 36728
rect 9812 36688 9813 36728
rect 9771 36679 9813 36688
rect 9868 36728 9908 38200
rect 10060 37820 10100 39880
rect 10156 39761 10196 41476
rect 10252 41348 10292 41357
rect 10292 41308 10388 41348
rect 10252 41299 10292 41308
rect 10155 39752 10197 39761
rect 10155 39712 10156 39752
rect 10196 39712 10197 39752
rect 10155 39703 10197 39712
rect 10155 39080 10197 39089
rect 10155 39040 10156 39080
rect 10196 39040 10197 39080
rect 10155 39031 10197 39040
rect 10156 38240 10196 39031
rect 10251 38996 10293 39005
rect 10251 38956 10252 38996
rect 10292 38956 10293 38996
rect 10251 38947 10293 38956
rect 10252 38912 10292 38947
rect 10252 38585 10292 38872
rect 10251 38576 10293 38585
rect 10251 38536 10252 38576
rect 10292 38536 10293 38576
rect 10251 38527 10293 38536
rect 10156 38191 10196 38200
rect 10251 38240 10293 38249
rect 10251 38200 10252 38240
rect 10292 38200 10293 38240
rect 10251 38191 10293 38200
rect 10252 37820 10292 38191
rect 9772 36594 9812 36679
rect 9868 36569 9908 36688
rect 9964 37780 10100 37820
rect 10156 37780 10292 37820
rect 9867 36560 9909 36569
rect 9867 36520 9868 36560
rect 9908 36520 9909 36560
rect 9867 36511 9909 36520
rect 9675 35888 9717 35897
rect 9675 35848 9676 35888
rect 9716 35848 9717 35888
rect 9675 35839 9717 35848
rect 9676 35754 9716 35839
rect 9771 35804 9813 35813
rect 9771 35764 9772 35804
rect 9812 35764 9813 35804
rect 9771 35755 9813 35764
rect 9772 35670 9812 35755
rect 9771 35300 9813 35309
rect 9771 35260 9772 35300
rect 9812 35260 9813 35300
rect 9771 35251 9813 35260
rect 9676 35216 9716 35225
rect 9484 35092 9620 35132
rect 9387 34460 9429 34469
rect 9387 34420 9388 34460
rect 9428 34420 9429 34460
rect 9387 34411 9429 34420
rect 9580 34385 9620 35092
rect 9676 35057 9716 35176
rect 9772 35166 9812 35251
rect 9867 35216 9909 35225
rect 9867 35176 9868 35216
rect 9908 35176 9909 35216
rect 9867 35167 9909 35176
rect 9868 35057 9908 35167
rect 9675 35048 9717 35057
rect 9675 35008 9676 35048
rect 9716 35008 9717 35048
rect 9675 34999 9717 35008
rect 9867 35048 9909 35057
rect 9867 35008 9868 35048
rect 9908 35008 9909 35048
rect 9867 34999 9909 35008
rect 9675 34796 9717 34805
rect 9675 34756 9676 34796
rect 9716 34756 9717 34796
rect 9675 34747 9717 34756
rect 9579 34376 9621 34385
rect 9579 34336 9580 34376
rect 9620 34336 9621 34376
rect 9579 34327 9621 34336
rect 9387 34292 9429 34301
rect 9387 34252 9388 34292
rect 9428 34252 9429 34292
rect 9387 34243 9429 34252
rect 9388 30932 9428 34243
rect 9483 34124 9525 34133
rect 9483 34084 9484 34124
rect 9524 34084 9525 34124
rect 9483 34075 9525 34084
rect 9484 33704 9524 34075
rect 9484 33655 9524 33664
rect 9580 33704 9620 34327
rect 9580 33655 9620 33664
rect 9676 33368 9716 34747
rect 9771 34544 9813 34553
rect 9771 34504 9772 34544
rect 9812 34504 9813 34544
rect 9771 34495 9813 34504
rect 9772 34376 9812 34495
rect 9772 34327 9812 34336
rect 9771 34040 9813 34049
rect 9771 34000 9772 34040
rect 9812 34000 9813 34040
rect 9771 33991 9813 34000
rect 9580 33328 9716 33368
rect 9772 33872 9812 33991
rect 9868 33956 9908 34999
rect 9964 34805 10004 37780
rect 10156 37568 10196 37780
rect 10156 37519 10196 37528
rect 10060 37232 10100 37241
rect 10060 36569 10100 37192
rect 10348 36737 10388 41308
rect 10444 39752 10484 45088
rect 10444 39703 10484 39712
rect 10443 38744 10485 38753
rect 10443 38704 10444 38744
rect 10484 38704 10485 38744
rect 10443 38695 10485 38704
rect 10444 38610 10484 38695
rect 10540 37400 10580 45172
rect 10636 40424 10676 45256
rect 10732 45053 10772 46348
rect 10923 46348 10924 46388
rect 10964 46348 10965 46388
rect 10923 46339 10965 46348
rect 10827 45800 10869 45809
rect 10827 45760 10828 45800
rect 10868 45760 10869 45800
rect 10827 45751 10869 45760
rect 10828 45666 10868 45751
rect 10924 45473 10964 46339
rect 11019 45632 11061 45641
rect 11019 45592 11020 45632
rect 11060 45592 11061 45632
rect 11019 45583 11061 45592
rect 11020 45498 11060 45583
rect 10923 45464 10965 45473
rect 10923 45424 10924 45464
rect 10964 45424 10965 45464
rect 10923 45415 10965 45424
rect 10731 45044 10773 45053
rect 10731 45004 10732 45044
rect 10772 45004 10773 45044
rect 10731 44995 10773 45004
rect 10924 43709 10964 45415
rect 10923 43700 10965 43709
rect 10923 43660 10924 43700
rect 10964 43660 10965 43700
rect 10923 43651 10965 43660
rect 10731 42776 10773 42785
rect 10731 42736 10732 42776
rect 10772 42736 10773 42776
rect 10731 42727 10773 42736
rect 10732 42642 10772 42727
rect 10731 41936 10773 41945
rect 10731 41896 10732 41936
rect 10772 41896 10773 41936
rect 10731 41887 10773 41896
rect 10732 41802 10772 41887
rect 11116 41021 11156 46600
rect 11211 46472 11253 46481
rect 11211 46432 11212 46472
rect 11252 46432 11253 46472
rect 11211 46423 11253 46432
rect 11212 46338 11252 46423
rect 11212 45800 11252 45809
rect 11212 45305 11252 45760
rect 11211 45296 11253 45305
rect 11211 45256 11212 45296
rect 11252 45256 11253 45296
rect 11211 45247 11253 45256
rect 11403 45212 11445 45221
rect 11403 45172 11404 45212
rect 11444 45172 11445 45212
rect 11403 45163 11445 45172
rect 11404 44960 11444 45163
rect 11404 44911 11444 44920
rect 11307 43448 11349 43457
rect 11307 43408 11308 43448
rect 11348 43408 11349 43448
rect 11307 43399 11349 43408
rect 11308 43314 11348 43399
rect 11212 41941 11252 41950
rect 11115 41012 11157 41021
rect 11115 40972 11116 41012
rect 11156 40972 11157 41012
rect 11115 40963 11157 40972
rect 11212 40685 11252 41901
rect 11404 41768 11444 41777
rect 11211 40676 11253 40685
rect 11211 40636 11212 40676
rect 11252 40636 11253 40676
rect 11211 40627 11253 40636
rect 10732 40424 10772 40433
rect 10636 40384 10732 40424
rect 10732 38417 10772 40384
rect 11404 39929 11444 41728
rect 11500 41693 11540 47776
rect 11595 46556 11637 46565
rect 11595 46516 11596 46556
rect 11636 46516 11637 46556
rect 11595 46507 11637 46516
rect 11596 45725 11636 46507
rect 11692 46477 11732 46486
rect 11595 45716 11637 45725
rect 11595 45676 11596 45716
rect 11636 45676 11637 45716
rect 11595 45667 11637 45676
rect 11692 45641 11732 46437
rect 11884 46472 11924 48439
rect 11980 46649 12020 52891
rect 11979 46640 12021 46649
rect 11979 46600 11980 46640
rect 12020 46600 12021 46640
rect 11979 46591 12021 46600
rect 12076 46481 12116 53983
rect 12172 50345 12212 57931
rect 12268 52520 12308 58612
rect 12363 57056 12405 57065
rect 12363 57016 12364 57056
rect 12404 57016 12405 57056
rect 12363 57007 12405 57016
rect 12364 53117 12404 57007
rect 12459 56384 12501 56393
rect 12459 56344 12460 56384
rect 12500 56344 12501 56384
rect 12459 56335 12501 56344
rect 12460 55637 12500 56335
rect 12459 55628 12501 55637
rect 12459 55588 12460 55628
rect 12500 55588 12501 55628
rect 12459 55579 12501 55588
rect 12460 54032 12500 55579
rect 12460 53705 12500 53992
rect 12459 53696 12501 53705
rect 12459 53656 12460 53696
rect 12500 53656 12501 53696
rect 12459 53647 12501 53656
rect 12556 53528 12596 59284
rect 12652 54041 12692 60367
rect 12844 60341 12884 76831
rect 13132 76754 13172 76806
rect 13228 76754 13268 79024
rect 13324 76973 13364 80536
rect 13419 80240 13461 80249
rect 13419 80200 13420 80240
rect 13460 80200 13461 80240
rect 13419 80191 13461 80200
rect 13420 79736 13460 80191
rect 13420 79409 13460 79696
rect 13419 79400 13461 79409
rect 13419 79360 13420 79400
rect 13460 79360 13461 79400
rect 13419 79351 13461 79360
rect 13516 77468 13556 81880
rect 13803 81332 13845 81341
rect 13803 81292 13804 81332
rect 13844 81292 13845 81332
rect 13803 81283 13845 81292
rect 13707 79568 13749 79577
rect 13707 79528 13708 79568
rect 13748 79528 13749 79568
rect 13707 79519 13749 79528
rect 13708 79064 13748 79519
rect 13420 77428 13556 77468
rect 13612 78980 13652 78989
rect 13323 76964 13365 76973
rect 13323 76924 13324 76964
rect 13364 76924 13365 76964
rect 13323 76915 13365 76924
rect 13132 76726 13268 76754
rect 13036 76712 13076 76721
rect 12940 76672 13036 76712
rect 13127 76714 13268 76726
rect 13127 76712 13173 76714
rect 13127 76672 13132 76712
rect 13172 76672 13173 76712
rect 12940 75872 12980 76672
rect 13036 76663 13076 76672
rect 13131 76663 13173 76672
rect 13131 76544 13171 76663
rect 13420 76544 13460 77428
rect 13612 76880 13652 78940
rect 13708 76889 13748 79024
rect 13516 76840 13652 76880
rect 13707 76880 13749 76889
rect 13707 76840 13708 76880
rect 13748 76840 13749 76880
rect 13516 76721 13556 76840
rect 13707 76831 13749 76840
rect 13515 76712 13557 76721
rect 13515 76672 13516 76712
rect 13556 76672 13557 76712
rect 13515 76663 13557 76672
rect 13612 76712 13652 76721
rect 13708 76712 13748 76831
rect 13652 76672 13748 76712
rect 13612 76663 13652 76672
rect 13131 76504 13172 76544
rect 13420 76504 13556 76544
rect 13132 75872 13172 76504
rect 13419 76292 13461 76301
rect 13419 76252 13420 76292
rect 13460 76252 13461 76292
rect 13419 76243 13461 76252
rect 13323 76208 13365 76217
rect 13323 76168 13324 76208
rect 13364 76168 13365 76208
rect 13323 76159 13365 76168
rect 13324 76040 13364 76159
rect 13324 75991 13364 76000
rect 13132 75832 13364 75872
rect 12940 75823 12980 75832
rect 12939 75536 12981 75545
rect 12939 75496 12940 75536
rect 12980 75496 12981 75536
rect 12939 75487 12981 75496
rect 12940 74108 12980 75487
rect 13035 75200 13077 75209
rect 13035 75160 13036 75200
rect 13076 75160 13077 75200
rect 13035 75151 13077 75160
rect 13036 75066 13076 75151
rect 13131 74444 13173 74453
rect 13131 74404 13132 74444
rect 13172 74404 13173 74444
rect 13131 74395 13173 74404
rect 13228 74444 13268 74453
rect 13132 74310 13172 74395
rect 12940 74068 13076 74108
rect 12939 73940 12981 73949
rect 12939 73900 12940 73940
rect 12980 73900 12981 73940
rect 12939 73891 12981 73900
rect 12940 73702 12980 73891
rect 12940 73653 12980 73662
rect 13036 73604 13076 74068
rect 13228 73865 13268 74404
rect 13227 73856 13269 73865
rect 13227 73816 13228 73856
rect 13268 73816 13269 73856
rect 13227 73807 13269 73816
rect 12940 73564 13076 73604
rect 13131 73604 13173 73613
rect 13131 73564 13132 73604
rect 13172 73564 13173 73604
rect 12940 67649 12980 73564
rect 13131 73555 13173 73564
rect 13132 73470 13172 73555
rect 13035 73436 13077 73445
rect 13035 73396 13036 73436
rect 13076 73396 13077 73436
rect 13035 73387 13077 73396
rect 13036 73016 13076 73387
rect 13132 73016 13172 73044
rect 13036 72976 13132 73016
rect 13036 71513 13076 72976
rect 13132 72967 13172 72976
rect 13227 72260 13269 72269
rect 13227 72220 13228 72260
rect 13268 72220 13269 72260
rect 13227 72211 13269 72220
rect 13131 72176 13173 72185
rect 13131 72136 13132 72176
rect 13172 72136 13173 72176
rect 13131 72127 13173 72136
rect 13228 72176 13268 72211
rect 13035 71504 13077 71513
rect 13035 71464 13036 71504
rect 13076 71464 13077 71504
rect 13035 71455 13077 71464
rect 13036 71370 13076 71455
rect 13132 70832 13172 72127
rect 13228 72125 13268 72136
rect 13227 72008 13269 72017
rect 13227 71968 13228 72008
rect 13268 71968 13269 72008
rect 13227 71959 13269 71968
rect 13036 70792 13172 70832
rect 12939 67640 12981 67649
rect 12939 67600 12940 67640
rect 12980 67600 12981 67640
rect 12939 67591 12981 67600
rect 13036 67640 13076 70792
rect 13228 70664 13268 71959
rect 13228 70615 13268 70624
rect 13324 69236 13364 75832
rect 13420 74117 13460 76243
rect 13419 74108 13461 74117
rect 13419 74068 13420 74108
rect 13460 74068 13461 74108
rect 13419 74059 13461 74068
rect 13419 73940 13461 73949
rect 13419 73900 13420 73940
rect 13460 73900 13461 73940
rect 13419 73891 13461 73900
rect 13420 73688 13460 73891
rect 13420 73639 13460 73648
rect 13419 72008 13461 72017
rect 13419 71968 13420 72008
rect 13460 71968 13461 72008
rect 13419 71959 13461 71968
rect 13420 71874 13460 71959
rect 13516 71756 13556 76504
rect 13611 76124 13653 76133
rect 13611 76084 13612 76124
rect 13652 76084 13653 76124
rect 13611 76075 13653 76084
rect 13612 73100 13652 76075
rect 13708 74528 13748 74537
rect 13708 73445 13748 74488
rect 13804 74201 13844 81283
rect 13900 75209 13940 82795
rect 14283 82256 14325 82265
rect 14283 82216 14284 82256
rect 14324 82216 14325 82256
rect 14283 82207 14325 82216
rect 14284 82122 14324 82207
rect 14092 82004 14132 82013
rect 14092 79745 14132 81964
rect 15340 81929 15380 83476
rect 15723 83096 15765 83105
rect 15723 83056 15724 83096
rect 15764 83056 15765 83096
rect 15723 83047 15765 83056
rect 15724 82256 15764 83047
rect 15724 82207 15764 82216
rect 15532 82004 15572 82013
rect 15436 81964 15532 82004
rect 15339 81920 15381 81929
rect 15339 81880 15340 81920
rect 15380 81880 15381 81920
rect 15339 81871 15381 81880
rect 14476 80576 14516 80585
rect 14516 80536 14612 80576
rect 14476 80527 14516 80536
rect 14283 79820 14325 79829
rect 14283 79780 14284 79820
rect 14324 79780 14325 79820
rect 14283 79771 14325 79780
rect 14091 79736 14133 79745
rect 14091 79696 14092 79736
rect 14132 79696 14133 79736
rect 14091 79687 14133 79696
rect 14187 79316 14229 79325
rect 14187 79276 14188 79316
rect 14228 79276 14229 79316
rect 14187 79267 14229 79276
rect 14188 79064 14228 79267
rect 14092 79024 14188 79064
rect 14092 78233 14132 79024
rect 14188 79015 14228 79024
rect 14091 78224 14133 78233
rect 14091 78184 14092 78224
rect 14132 78184 14133 78224
rect 14091 78175 14133 78184
rect 14092 76721 14132 78175
rect 14284 77552 14324 79771
rect 14572 79736 14612 80536
rect 14668 80324 14708 80333
rect 14708 80284 14804 80324
rect 14668 80275 14708 80284
rect 14668 79736 14708 79745
rect 14572 79696 14668 79736
rect 14572 79409 14612 79696
rect 14668 79687 14708 79696
rect 14571 79400 14613 79409
rect 14571 79360 14572 79400
rect 14612 79360 14613 79400
rect 14571 79351 14613 79360
rect 14572 78149 14612 79351
rect 14764 79064 14804 80284
rect 14860 79568 14900 79577
rect 14900 79528 14996 79568
rect 14860 79519 14900 79528
rect 14716 79054 14804 79064
rect 14756 79024 14804 79054
rect 14860 79148 14900 79157
rect 14716 79005 14756 79014
rect 14379 78140 14421 78149
rect 14379 78100 14380 78140
rect 14420 78100 14421 78140
rect 14379 78091 14421 78100
rect 14571 78140 14613 78149
rect 14763 78140 14805 78149
rect 14571 78100 14572 78140
rect 14612 78100 14613 78140
rect 14571 78091 14613 78100
rect 14668 78100 14764 78140
rect 14804 78100 14805 78140
rect 14284 77503 14324 77512
rect 14091 76712 14133 76721
rect 14091 76672 14092 76712
rect 14132 76672 14133 76712
rect 14091 76663 14133 76672
rect 14092 76578 14132 76663
rect 14380 76040 14420 78091
rect 14476 77300 14516 77309
rect 14516 77260 14612 77300
rect 14476 77251 14516 77260
rect 14572 76726 14612 77260
rect 14572 76677 14612 76686
rect 14572 76040 14612 76049
rect 14380 76000 14572 76040
rect 14091 75620 14133 75629
rect 14091 75580 14092 75620
rect 14132 75580 14133 75620
rect 14091 75571 14133 75580
rect 13899 75200 13941 75209
rect 13899 75160 13900 75200
rect 13940 75160 13941 75200
rect 13899 75151 13941 75160
rect 13803 74192 13845 74201
rect 13803 74152 13804 74192
rect 13844 74152 13845 74192
rect 13803 74143 13845 74152
rect 13707 73436 13749 73445
rect 13707 73396 13708 73436
rect 13748 73396 13749 73436
rect 13707 73387 13749 73396
rect 13803 73100 13845 73109
rect 13612 73060 13748 73100
rect 13612 73002 13652 73011
rect 13612 72773 13652 72962
rect 13611 72764 13653 72773
rect 13611 72724 13612 72764
rect 13652 72724 13653 72764
rect 13611 72715 13653 72724
rect 13708 72101 13748 73060
rect 13803 73060 13804 73100
rect 13844 73060 13845 73100
rect 13803 73051 13845 73060
rect 13804 72966 13844 73051
rect 13900 72185 13940 75151
rect 14092 74957 14132 75571
rect 14572 75293 14612 76000
rect 14283 75284 14325 75293
rect 14283 75244 14284 75284
rect 14324 75244 14325 75284
rect 14283 75235 14325 75244
rect 14571 75284 14613 75293
rect 14571 75244 14572 75284
rect 14612 75244 14613 75284
rect 14571 75235 14613 75244
rect 14284 75200 14324 75235
rect 14284 75149 14324 75160
rect 14476 75032 14516 75041
rect 14284 74992 14476 75032
rect 14091 74948 14133 74957
rect 14091 74908 14092 74948
rect 14132 74908 14133 74948
rect 14091 74899 14133 74908
rect 13899 72176 13941 72185
rect 13899 72136 13900 72176
rect 13940 72136 13941 72176
rect 13899 72127 13941 72136
rect 13707 72092 13749 72101
rect 13707 72052 13708 72092
rect 13748 72052 13749 72092
rect 13707 72043 13749 72052
rect 13900 72042 13940 72127
rect 13995 72008 14037 72017
rect 13995 71968 13996 72008
rect 14036 71968 14037 72008
rect 13995 71959 14037 71968
rect 13899 71840 13941 71849
rect 13899 71800 13900 71840
rect 13940 71800 13941 71840
rect 13899 71791 13941 71800
rect 13516 71716 13844 71756
rect 13707 71588 13749 71597
rect 13707 71548 13708 71588
rect 13748 71548 13749 71588
rect 13707 71539 13749 71548
rect 13516 71490 13556 71499
rect 13420 70916 13460 70925
rect 13516 70916 13556 71450
rect 13708 70925 13748 71539
rect 13460 70876 13556 70916
rect 13707 70916 13749 70925
rect 13707 70876 13708 70916
rect 13748 70876 13749 70916
rect 13420 70867 13460 70876
rect 13707 70867 13749 70876
rect 13515 69992 13557 70001
rect 13515 69952 13516 69992
rect 13556 69952 13557 69992
rect 13515 69943 13557 69952
rect 13516 69858 13556 69943
rect 13228 69196 13364 69236
rect 13131 69152 13173 69161
rect 13131 69112 13132 69152
rect 13172 69112 13173 69152
rect 13131 69103 13173 69112
rect 13132 69018 13172 69103
rect 13228 68648 13268 69196
rect 13612 69152 13652 69161
rect 13324 69068 13364 69077
rect 13612 69068 13652 69112
rect 13707 69152 13749 69161
rect 13707 69112 13708 69152
rect 13748 69112 13749 69152
rect 13707 69103 13749 69112
rect 13364 69028 13652 69068
rect 13324 69019 13364 69028
rect 13036 67472 13076 67600
rect 12940 67432 13076 67472
rect 13132 68608 13268 68648
rect 12940 66800 12980 67432
rect 13036 66977 13076 67062
rect 13035 66968 13077 66977
rect 13035 66928 13036 66968
rect 13076 66928 13077 66968
rect 13035 66919 13077 66928
rect 12940 66760 13076 66800
rect 13036 66473 13076 66760
rect 13035 66464 13077 66473
rect 13035 66424 13036 66464
rect 13076 66424 13077 66464
rect 13035 66415 13077 66424
rect 12939 65540 12981 65549
rect 12939 65500 12940 65540
rect 12980 65500 12981 65540
rect 12939 65491 12981 65500
rect 12843 60332 12885 60341
rect 12843 60292 12844 60332
rect 12884 60292 12885 60332
rect 12843 60283 12885 60292
rect 12940 60173 12980 65491
rect 13036 61265 13076 66415
rect 13035 61256 13077 61265
rect 13035 61216 13036 61256
rect 13076 61216 13077 61256
rect 13035 61207 13077 61216
rect 13132 60248 13172 68608
rect 13419 67640 13461 67649
rect 13419 67600 13420 67640
rect 13460 67600 13461 67640
rect 13419 67591 13461 67600
rect 13420 67506 13460 67591
rect 13228 67052 13268 67061
rect 13268 67012 13556 67052
rect 13228 67003 13268 67012
rect 13516 66988 13556 67012
rect 13516 66939 13556 66948
rect 13612 66968 13652 66977
rect 13708 66968 13748 69103
rect 13652 66928 13748 66968
rect 13612 66884 13652 66928
rect 13324 66844 13652 66884
rect 13324 63953 13364 66844
rect 13804 66800 13844 71716
rect 13900 70664 13940 71791
rect 13996 71504 14036 71959
rect 14092 71672 14132 74899
rect 14284 74528 14324 74992
rect 14476 74983 14516 74992
rect 14236 74518 14324 74528
rect 14276 74488 14324 74518
rect 14380 74612 14420 74621
rect 14236 74469 14276 74478
rect 14380 74369 14420 74572
rect 14379 74360 14421 74369
rect 14379 74320 14380 74360
rect 14420 74320 14421 74360
rect 14379 74311 14421 74320
rect 14668 74192 14708 78100
rect 14763 78091 14805 78100
rect 14860 76628 14900 79108
rect 14956 78224 14996 79528
rect 15436 79484 15476 81964
rect 15532 81955 15572 81964
rect 15724 79988 15764 79997
rect 15820 79988 15860 85936
rect 15915 83516 15957 83525
rect 15915 83476 15916 83516
rect 15956 83476 15957 83516
rect 15915 83467 15957 83476
rect 15916 83382 15956 83467
rect 15764 79948 15860 79988
rect 15916 79988 15956 79997
rect 16012 79988 16052 85936
rect 15956 79948 16052 79988
rect 15724 79939 15764 79948
rect 15916 79939 15956 79948
rect 15531 79820 15573 79829
rect 15531 79780 15532 79820
rect 15572 79780 15573 79820
rect 15531 79771 15573 79780
rect 15915 79820 15957 79829
rect 15915 79780 15916 79820
rect 15956 79780 15957 79820
rect 15915 79771 15957 79780
rect 16108 79820 16148 79829
rect 15532 79686 15572 79771
rect 15244 79444 15476 79484
rect 15244 78905 15284 79444
rect 15339 79316 15381 79325
rect 15339 79276 15340 79316
rect 15380 79276 15381 79316
rect 15339 79267 15381 79276
rect 15340 79064 15380 79267
rect 15243 78896 15285 78905
rect 15243 78856 15244 78896
rect 15284 78856 15285 78896
rect 15243 78847 15285 78856
rect 14956 78175 14996 78184
rect 15052 78224 15092 78233
rect 15092 78184 15188 78224
rect 15052 78175 15092 78184
rect 15051 78056 15093 78065
rect 15051 78016 15052 78056
rect 15092 78016 15093 78056
rect 15051 78007 15093 78016
rect 15052 77552 15092 78007
rect 15052 77503 15092 77512
rect 15052 76712 15092 76721
rect 14860 76588 14996 76628
rect 14764 76544 14804 76553
rect 14804 76504 14900 76544
rect 14764 76495 14804 76504
rect 14763 76208 14805 76217
rect 14763 76168 14764 76208
rect 14804 76168 14805 76208
rect 14763 76159 14805 76168
rect 14764 76074 14804 76159
rect 14860 74780 14900 76504
rect 14380 74152 14708 74192
rect 14764 74740 14900 74780
rect 14187 74024 14229 74033
rect 14187 73984 14188 74024
rect 14228 73984 14229 74024
rect 14187 73975 14229 73984
rect 14188 71849 14228 73975
rect 14283 73856 14325 73865
rect 14283 73816 14284 73856
rect 14324 73816 14325 73856
rect 14283 73807 14325 73816
rect 14284 73613 14324 73807
rect 14283 73604 14325 73613
rect 14283 73564 14284 73604
rect 14324 73564 14325 73604
rect 14283 73555 14325 73564
rect 14187 71840 14229 71849
rect 14187 71800 14188 71840
rect 14228 71800 14229 71840
rect 14187 71791 14229 71800
rect 14092 71632 14228 71672
rect 13996 71455 14036 71464
rect 14092 71504 14132 71513
rect 14092 71345 14132 71464
rect 14091 71336 14133 71345
rect 14091 71296 14092 71336
rect 14132 71296 14133 71336
rect 14091 71287 14133 71296
rect 14188 71168 14228 71632
rect 14092 71128 14228 71168
rect 13940 70624 14036 70664
rect 13900 70615 13940 70624
rect 13899 69992 13941 70001
rect 13899 69952 13900 69992
rect 13940 69952 13941 69992
rect 13899 69943 13941 69952
rect 13516 66760 13844 66800
rect 13323 63944 13365 63953
rect 13323 63904 13324 63944
rect 13364 63904 13365 63944
rect 13323 63895 13365 63904
rect 13419 63608 13461 63617
rect 13419 63568 13420 63608
rect 13460 63568 13461 63608
rect 13419 63559 13461 63568
rect 13323 61760 13365 61769
rect 13323 61720 13324 61760
rect 13364 61720 13365 61760
rect 13323 61711 13365 61720
rect 13324 60920 13364 61711
rect 13324 60509 13364 60880
rect 13323 60500 13365 60509
rect 13323 60460 13324 60500
rect 13364 60460 13365 60500
rect 13323 60451 13365 60460
rect 13132 60208 13364 60248
rect 12939 60164 12981 60173
rect 12939 60124 12940 60164
rect 12980 60124 12981 60164
rect 12939 60115 12981 60124
rect 13324 60089 13364 60208
rect 12747 60080 12789 60089
rect 12747 60040 12748 60080
rect 12788 60040 12789 60080
rect 12747 60031 12789 60040
rect 13228 60080 13268 60089
rect 12748 59946 12788 60031
rect 12843 59996 12885 60005
rect 12843 59956 12844 59996
rect 12884 59956 12885 59996
rect 12843 59947 12885 59956
rect 12940 59996 12980 60005
rect 13228 59996 13268 60040
rect 13323 60080 13365 60089
rect 13323 60040 13324 60080
rect 13364 60040 13365 60080
rect 13323 60031 13365 60040
rect 12980 59956 13268 59996
rect 12940 59947 12980 59956
rect 12747 58568 12789 58577
rect 12747 58528 12748 58568
rect 12788 58528 12789 58568
rect 12747 58519 12789 58528
rect 12748 58434 12788 58519
rect 12747 58064 12789 58073
rect 12747 58024 12748 58064
rect 12788 58024 12789 58064
rect 12747 58015 12789 58024
rect 12748 54788 12788 58015
rect 12844 54872 12884 59947
rect 13324 59946 13364 60031
rect 12939 59828 12981 59837
rect 12939 59788 12940 59828
rect 12980 59788 12981 59828
rect 12939 59779 12981 59788
rect 12940 55460 12980 59779
rect 13420 58829 13460 63559
rect 13419 58820 13461 58829
rect 13419 58780 13420 58820
rect 13460 58780 13461 58820
rect 13419 58771 13461 58780
rect 13419 58652 13461 58661
rect 13419 58612 13420 58652
rect 13460 58612 13461 58652
rect 13419 58603 13461 58612
rect 13276 58577 13316 58586
rect 13316 58537 13364 58568
rect 13276 58528 13364 58537
rect 13324 58064 13364 58528
rect 13420 58484 13460 58603
rect 13420 58435 13460 58444
rect 13324 58015 13364 58024
rect 13131 57896 13173 57905
rect 13131 57856 13132 57896
rect 13172 57856 13173 57896
rect 13131 57847 13173 57856
rect 13132 57762 13172 57847
rect 13516 57317 13556 66760
rect 13611 66632 13653 66641
rect 13611 66592 13612 66632
rect 13652 66592 13653 66632
rect 13611 66583 13653 66592
rect 13612 66137 13652 66583
rect 13611 66128 13653 66137
rect 13611 66088 13612 66128
rect 13652 66088 13653 66128
rect 13611 66079 13653 66088
rect 13900 66128 13940 69943
rect 13996 69413 14036 70624
rect 14092 70589 14132 71128
rect 14187 70916 14229 70925
rect 14187 70876 14188 70916
rect 14228 70876 14229 70916
rect 14187 70867 14229 70876
rect 14091 70580 14133 70589
rect 14091 70540 14092 70580
rect 14132 70540 14133 70580
rect 14091 70531 14133 70540
rect 13995 69404 14037 69413
rect 13995 69364 13996 69404
rect 14036 69364 14037 69404
rect 13995 69355 14037 69364
rect 14092 69152 14132 69161
rect 13996 69112 14092 69152
rect 13996 66968 14036 69112
rect 14092 69103 14132 69112
rect 14188 69152 14228 70867
rect 14284 69236 14324 73555
rect 14380 70001 14420 74152
rect 14667 73688 14709 73697
rect 14667 73648 14668 73688
rect 14708 73648 14709 73688
rect 14667 73639 14709 73648
rect 14668 73554 14708 73639
rect 14764 71597 14804 74740
rect 14956 74621 14996 76588
rect 15052 76217 15092 76672
rect 15148 76712 15188 78184
rect 15244 78149 15284 78847
rect 15243 78140 15285 78149
rect 15243 78100 15244 78140
rect 15284 78100 15285 78140
rect 15243 78091 15285 78100
rect 15148 76637 15188 76672
rect 15147 76628 15189 76637
rect 15147 76588 15148 76628
rect 15188 76588 15189 76628
rect 15147 76579 15189 76588
rect 15340 76385 15380 79024
rect 15436 78224 15476 78233
rect 15436 77972 15476 78184
rect 15532 78224 15572 78233
rect 15572 78184 15668 78224
rect 15532 78175 15572 78184
rect 15436 77932 15572 77972
rect 15435 77384 15477 77393
rect 15435 77344 15436 77384
rect 15476 77344 15477 77384
rect 15435 77335 15477 77344
rect 15339 76376 15381 76385
rect 15339 76336 15340 76376
rect 15380 76336 15381 76376
rect 15339 76327 15381 76336
rect 15051 76208 15093 76217
rect 15051 76168 15052 76208
rect 15092 76168 15093 76208
rect 15051 76159 15093 76168
rect 15243 76040 15285 76049
rect 15243 76000 15244 76040
rect 15284 76000 15285 76040
rect 15243 75991 15285 76000
rect 15244 75956 15284 75991
rect 15244 75905 15284 75916
rect 15340 75704 15380 76327
rect 15436 76208 15476 77335
rect 15436 76159 15476 76168
rect 15532 76712 15572 77932
rect 15628 76889 15668 78184
rect 15723 77300 15765 77309
rect 15723 77260 15724 77300
rect 15764 77260 15765 77300
rect 15723 77251 15765 77260
rect 15627 76880 15669 76889
rect 15627 76840 15628 76880
rect 15668 76840 15669 76880
rect 15627 76831 15669 76840
rect 15628 76796 15668 76831
rect 15628 76745 15668 76756
rect 15052 75664 15380 75704
rect 14955 74612 14997 74621
rect 14955 74572 14956 74612
rect 14996 74572 14997 74612
rect 14955 74563 14997 74572
rect 14859 73940 14901 73949
rect 14859 73900 14860 73940
rect 14900 73900 14901 73940
rect 14859 73891 14901 73900
rect 14860 73806 14900 73891
rect 14956 73688 14996 74563
rect 15052 74192 15092 75664
rect 15339 75536 15381 75545
rect 15339 75496 15340 75536
rect 15380 75496 15381 75536
rect 15339 75487 15381 75496
rect 15340 75200 15380 75487
rect 15340 75151 15380 75160
rect 15244 74528 15284 74537
rect 15052 74152 15188 74192
rect 15051 74024 15093 74033
rect 15051 73984 15052 74024
rect 15092 73984 15093 74024
rect 15051 73975 15093 73984
rect 14860 73648 14996 73688
rect 15052 73688 15092 73975
rect 14763 71588 14805 71597
rect 14763 71548 14764 71588
rect 14804 71548 14805 71588
rect 14763 71539 14805 71548
rect 14475 71504 14517 71513
rect 14475 71464 14476 71504
rect 14516 71464 14517 71504
rect 14475 71455 14517 71464
rect 14476 71370 14516 71455
rect 14572 71420 14612 71429
rect 14860 71420 14900 73648
rect 15052 73639 15092 73648
rect 15148 73520 15188 74152
rect 15244 73949 15284 74488
rect 15339 74528 15381 74537
rect 15532 74528 15572 76672
rect 15724 76208 15764 77251
rect 15628 76168 15764 76208
rect 15628 76040 15668 76168
rect 15628 75545 15668 76000
rect 15723 75956 15765 75965
rect 15723 75916 15724 75956
rect 15764 75916 15765 75956
rect 15723 75907 15765 75916
rect 15627 75536 15669 75545
rect 15627 75496 15628 75536
rect 15668 75496 15669 75536
rect 15627 75487 15669 75496
rect 15627 75284 15669 75293
rect 15627 75244 15628 75284
rect 15668 75244 15669 75284
rect 15627 75235 15669 75244
rect 15628 74705 15668 75235
rect 15627 74696 15669 74705
rect 15627 74656 15628 74696
rect 15668 74656 15669 74696
rect 15627 74647 15669 74656
rect 15339 74488 15340 74528
rect 15380 74488 15572 74528
rect 15339 74479 15381 74488
rect 15340 74394 15380 74479
rect 15628 74444 15668 74647
rect 15724 74528 15764 75907
rect 15724 74479 15764 74488
rect 15532 74404 15668 74444
rect 15820 74444 15860 74455
rect 15243 73940 15285 73949
rect 15243 73900 15244 73940
rect 15284 73900 15285 73940
rect 15243 73891 15285 73900
rect 15339 73688 15381 73697
rect 15339 73648 15340 73688
rect 15380 73648 15381 73688
rect 15339 73639 15381 73648
rect 14956 73480 15188 73520
rect 14956 73016 14996 73480
rect 14996 72976 15092 73016
rect 14956 72967 14996 72976
rect 14955 72176 14997 72185
rect 14955 72136 14956 72176
rect 14996 72136 14997 72176
rect 14955 72127 14997 72136
rect 14612 71380 14900 71420
rect 14379 69992 14421 70001
rect 14379 69952 14380 69992
rect 14420 69952 14421 69992
rect 14379 69943 14421 69952
rect 14284 69196 14516 69236
rect 14228 69112 14324 69152
rect 14188 69103 14228 69112
rect 14187 68984 14229 68993
rect 14187 68944 14188 68984
rect 14228 68944 14229 68984
rect 14187 68935 14229 68944
rect 14092 68480 14132 68489
rect 14092 68321 14132 68440
rect 14091 68312 14133 68321
rect 14091 68272 14092 68312
rect 14132 68272 14133 68312
rect 14091 68263 14133 68272
rect 14091 67136 14133 67145
rect 14091 67096 14092 67136
rect 14132 67096 14133 67136
rect 14091 67087 14133 67096
rect 13996 66389 14036 66928
rect 14092 66884 14132 67087
rect 14188 67052 14228 68935
rect 14284 67313 14324 69112
rect 14283 67304 14325 67313
rect 14283 67264 14284 67304
rect 14324 67264 14325 67304
rect 14283 67255 14325 67264
rect 14476 67145 14516 69196
rect 14572 68069 14612 71380
rect 14859 71084 14901 71093
rect 14859 71044 14860 71084
rect 14900 71044 14901 71084
rect 14859 71035 14901 71044
rect 14860 70925 14900 71035
rect 14859 70916 14901 70925
rect 14859 70876 14860 70916
rect 14900 70876 14901 70916
rect 14859 70867 14901 70876
rect 14860 70589 14900 70867
rect 14859 70580 14901 70589
rect 14859 70540 14860 70580
rect 14900 70540 14901 70580
rect 14859 70531 14901 70540
rect 14763 70496 14805 70505
rect 14763 70456 14764 70496
rect 14804 70456 14805 70496
rect 14763 70447 14805 70456
rect 14764 69992 14804 70447
rect 14668 69152 14708 69163
rect 14668 69077 14708 69112
rect 14667 69068 14709 69077
rect 14667 69028 14668 69068
rect 14708 69028 14709 69068
rect 14667 69019 14709 69028
rect 14764 68489 14804 69952
rect 14956 69917 14996 72127
rect 15052 71849 15092 72976
rect 15147 72932 15189 72941
rect 15147 72892 15148 72932
rect 15188 72892 15189 72932
rect 15147 72883 15189 72892
rect 15148 72353 15188 72883
rect 15147 72344 15189 72353
rect 15147 72304 15148 72344
rect 15188 72304 15189 72344
rect 15147 72295 15189 72304
rect 15243 72260 15285 72269
rect 15243 72220 15244 72260
rect 15284 72220 15285 72260
rect 15243 72211 15285 72220
rect 15147 72176 15189 72185
rect 15147 72136 15148 72176
rect 15188 72136 15189 72176
rect 15147 72127 15189 72136
rect 15051 71840 15093 71849
rect 15051 71800 15052 71840
rect 15092 71800 15093 71840
rect 15051 71791 15093 71800
rect 15051 71588 15093 71597
rect 15051 71548 15052 71588
rect 15092 71548 15093 71588
rect 15051 71539 15093 71548
rect 15052 71504 15092 71539
rect 14955 69908 14997 69917
rect 14955 69868 14956 69908
rect 14996 69868 14997 69908
rect 14955 69859 14997 69868
rect 14955 69740 14997 69749
rect 14955 69700 14956 69740
rect 14996 69700 14997 69740
rect 14955 69691 14997 69700
rect 14956 69606 14996 69691
rect 14763 68480 14805 68489
rect 14763 68440 14764 68480
rect 14804 68440 14805 68480
rect 14763 68431 14805 68440
rect 14571 68060 14613 68069
rect 14571 68020 14572 68060
rect 14612 68020 14613 68060
rect 14571 68011 14613 68020
rect 15052 67733 15092 71464
rect 15148 71345 15188 72127
rect 15147 71336 15189 71345
rect 15147 71296 15148 71336
rect 15188 71296 15189 71336
rect 15147 71287 15189 71296
rect 15148 70664 15188 71287
rect 15148 70505 15188 70624
rect 15147 70496 15189 70505
rect 15147 70456 15148 70496
rect 15188 70456 15189 70496
rect 15147 70447 15189 70456
rect 15147 69740 15189 69749
rect 15147 69700 15148 69740
rect 15188 69700 15189 69740
rect 15147 69691 15189 69700
rect 15148 69166 15188 69691
rect 15148 69117 15188 69126
rect 15244 69068 15284 72211
rect 15340 72185 15380 73639
rect 15339 72176 15381 72185
rect 15339 72136 15340 72176
rect 15380 72136 15381 72176
rect 15339 72127 15381 72136
rect 15532 72017 15572 74404
rect 15820 74369 15860 74404
rect 15819 74360 15861 74369
rect 15819 74320 15820 74360
rect 15860 74320 15861 74360
rect 15819 74311 15861 74320
rect 15819 74192 15861 74201
rect 15819 74152 15820 74192
rect 15860 74152 15861 74192
rect 15819 74143 15861 74152
rect 15627 73016 15669 73025
rect 15627 72976 15628 73016
rect 15668 72976 15669 73016
rect 15627 72967 15669 72976
rect 15340 72008 15380 72017
rect 15340 71849 15380 71968
rect 15531 72008 15573 72017
rect 15531 71968 15532 72008
rect 15572 71968 15573 72008
rect 15531 71959 15573 71968
rect 15339 71840 15381 71849
rect 15339 71800 15340 71840
rect 15380 71800 15381 71840
rect 15339 71791 15381 71800
rect 15531 71504 15573 71513
rect 15531 71459 15532 71504
rect 15572 71459 15573 71504
rect 15531 71455 15573 71459
rect 15532 71369 15572 71455
rect 15628 70664 15668 72967
rect 15723 71672 15765 71681
rect 15723 71632 15724 71672
rect 15764 71632 15765 71672
rect 15723 71623 15765 71632
rect 15724 71538 15764 71623
rect 15532 70624 15668 70664
rect 15339 70496 15381 70505
rect 15339 70456 15340 70496
rect 15380 70456 15381 70496
rect 15339 70447 15381 70456
rect 15340 70362 15380 70447
rect 15435 69992 15477 70001
rect 15435 69952 15436 69992
rect 15476 69952 15477 69992
rect 15435 69943 15477 69952
rect 15340 69068 15380 69077
rect 15244 69028 15340 69068
rect 15340 69019 15380 69028
rect 15147 68984 15189 68993
rect 15147 68944 15148 68984
rect 15188 68944 15189 68984
rect 15147 68935 15189 68944
rect 15051 67724 15093 67733
rect 15051 67684 15052 67724
rect 15092 67684 15093 67724
rect 15051 67675 15093 67684
rect 14571 67640 14613 67649
rect 14571 67600 14572 67640
rect 14612 67600 14613 67640
rect 14571 67591 14613 67600
rect 14668 67640 14708 67649
rect 14763 67640 14805 67649
rect 14708 67600 14764 67640
rect 14804 67600 14805 67640
rect 14668 67591 14708 67600
rect 14763 67591 14805 67600
rect 14572 67472 14612 67591
rect 14572 67432 14708 67472
rect 14475 67136 14517 67145
rect 14475 67096 14476 67136
rect 14516 67096 14517 67136
rect 14475 67087 14517 67096
rect 14188 67012 14324 67052
rect 13995 66380 14037 66389
rect 13995 66340 13996 66380
rect 14036 66340 14037 66380
rect 13995 66331 14037 66340
rect 13996 66128 14036 66137
rect 13900 66088 13996 66128
rect 13612 64616 13652 66079
rect 13804 65960 13844 65969
rect 13708 65920 13804 65960
rect 13708 65456 13748 65920
rect 13804 65911 13844 65920
rect 13900 65549 13940 66088
rect 13996 66079 14036 66088
rect 13899 65540 13941 65549
rect 13899 65500 13900 65540
rect 13940 65500 13941 65540
rect 13899 65491 13941 65500
rect 13708 65407 13748 65416
rect 13803 65456 13845 65465
rect 13803 65416 13804 65456
rect 13844 65416 13845 65456
rect 13803 65407 13845 65416
rect 13804 65288 13844 65407
rect 13612 64205 13652 64576
rect 13708 65248 13844 65288
rect 13708 64280 13748 65248
rect 13995 64616 14037 64625
rect 13995 64576 13996 64616
rect 14036 64576 14037 64616
rect 13995 64567 14037 64576
rect 13996 64482 14036 64567
rect 13804 64448 13844 64457
rect 13844 64408 13940 64448
rect 13804 64399 13844 64408
rect 13708 64240 13844 64280
rect 13611 64196 13653 64205
rect 13611 64156 13612 64196
rect 13652 64156 13653 64196
rect 13611 64147 13653 64156
rect 13612 63020 13652 64147
rect 13804 63776 13844 64240
rect 13900 63944 13940 64408
rect 13996 63953 14036 64038
rect 13900 63895 13940 63904
rect 13995 63944 14037 63953
rect 13995 63904 13996 63944
rect 14036 63904 14037 63944
rect 13995 63895 14037 63904
rect 13804 63736 14036 63776
rect 13803 63104 13845 63113
rect 13803 63064 13804 63104
rect 13844 63064 13845 63104
rect 13803 63055 13845 63064
rect 13707 63020 13749 63029
rect 13612 62980 13708 63020
rect 13748 62980 13749 63020
rect 13707 62971 13749 62980
rect 13611 62852 13653 62861
rect 13611 62812 13612 62852
rect 13652 62812 13653 62852
rect 13611 62803 13653 62812
rect 13612 58568 13652 62803
rect 13708 61592 13748 62971
rect 13804 62970 13844 63055
rect 13900 62432 13940 62441
rect 13900 61844 13940 62392
rect 13900 61795 13940 61804
rect 13996 62432 14036 63736
rect 13708 61543 13748 61552
rect 13899 61256 13941 61265
rect 13899 61216 13900 61256
rect 13940 61216 13941 61256
rect 13899 61207 13941 61216
rect 13803 60332 13845 60341
rect 13803 60292 13804 60332
rect 13844 60292 13845 60332
rect 13803 60283 13845 60292
rect 13804 60164 13844 60283
rect 13804 60115 13844 60124
rect 13708 60080 13748 60089
rect 13708 59921 13748 60040
rect 13707 59912 13749 59921
rect 13707 59872 13708 59912
rect 13748 59872 13749 59912
rect 13707 59863 13749 59872
rect 13803 59744 13845 59753
rect 13803 59704 13804 59744
rect 13844 59704 13845 59744
rect 13803 59695 13845 59704
rect 13707 59660 13749 59669
rect 13707 59620 13708 59660
rect 13748 59620 13749 59660
rect 13707 59611 13749 59620
rect 13708 58745 13748 59611
rect 13804 59249 13844 59695
rect 13803 59240 13845 59249
rect 13803 59200 13804 59240
rect 13844 59200 13845 59240
rect 13803 59191 13845 59200
rect 13707 58736 13749 58745
rect 13707 58696 13708 58736
rect 13748 58696 13749 58736
rect 13707 58687 13749 58696
rect 13708 58568 13748 58577
rect 13612 58528 13708 58568
rect 13515 57308 13557 57317
rect 13515 57268 13516 57308
rect 13556 57268 13557 57308
rect 13515 57259 13557 57268
rect 13227 57140 13269 57149
rect 13227 57100 13228 57140
rect 13268 57100 13269 57140
rect 13227 57091 13269 57100
rect 13228 57056 13268 57091
rect 13228 57005 13268 57016
rect 13419 56972 13461 56981
rect 13419 56932 13420 56972
rect 13460 56932 13461 56972
rect 13419 56923 13461 56932
rect 13420 56838 13460 56923
rect 13612 56729 13652 58528
rect 13708 58519 13748 58528
rect 13803 58484 13845 58493
rect 13803 58444 13804 58484
rect 13844 58444 13845 58484
rect 13803 58435 13845 58444
rect 13804 57812 13844 58435
rect 13900 57896 13940 61207
rect 13996 59669 14036 62392
rect 14092 62264 14132 66844
rect 14187 66380 14229 66389
rect 14187 66340 14188 66380
rect 14228 66340 14229 66380
rect 14187 66331 14229 66340
rect 14188 65456 14228 66331
rect 14188 62348 14228 65416
rect 14284 65456 14324 67012
rect 14572 66968 14612 66979
rect 14572 66893 14612 66928
rect 14571 66884 14613 66893
rect 14571 66844 14572 66884
rect 14612 66844 14613 66884
rect 14571 66835 14613 66844
rect 14284 64373 14324 65416
rect 14283 64364 14325 64373
rect 14283 64324 14284 64364
rect 14324 64324 14325 64364
rect 14283 64315 14325 64324
rect 14284 62516 14324 64315
rect 14668 64280 14708 67432
rect 14764 66977 14804 67591
rect 14860 67472 14900 67481
rect 14900 67432 15092 67472
rect 14860 67423 14900 67432
rect 14763 66968 14805 66977
rect 14763 66928 14764 66968
rect 14804 66928 14805 66968
rect 14763 66919 14805 66928
rect 15052 66963 15092 67432
rect 15052 66914 15092 66923
rect 15148 66893 15188 68935
rect 15339 68480 15381 68489
rect 15339 68440 15340 68480
rect 15380 68440 15381 68480
rect 15339 68431 15381 68440
rect 15340 68321 15380 68431
rect 15339 68312 15381 68321
rect 15339 68272 15340 68312
rect 15380 68272 15381 68312
rect 15339 68263 15381 68272
rect 15436 68060 15476 69943
rect 15532 68732 15572 70624
rect 15627 70496 15669 70505
rect 15627 70456 15628 70496
rect 15668 70456 15669 70496
rect 15627 70447 15669 70456
rect 15628 69992 15668 70447
rect 15628 69943 15668 69952
rect 15723 69992 15765 70001
rect 15723 69952 15724 69992
rect 15764 69952 15765 69992
rect 15723 69943 15765 69952
rect 15724 69858 15764 69943
rect 15532 68692 15764 68732
rect 15532 68237 15572 68322
rect 15531 68228 15573 68237
rect 15531 68188 15532 68228
rect 15572 68188 15573 68228
rect 15531 68179 15573 68188
rect 15436 68020 15572 68060
rect 15243 67136 15285 67145
rect 15243 67096 15244 67136
rect 15284 67096 15285 67136
rect 15243 67087 15285 67096
rect 15244 67002 15284 67087
rect 14955 66884 14997 66893
rect 14955 66844 14956 66884
rect 14996 66844 14997 66884
rect 14955 66835 14997 66844
rect 15147 66884 15189 66893
rect 15147 66844 15148 66884
rect 15188 66844 15189 66884
rect 15147 66835 15189 66844
rect 14764 65456 14804 65465
rect 14804 65416 14900 65456
rect 14764 65407 14804 65416
rect 14860 64280 14900 65416
rect 14572 64240 14708 64280
rect 14764 64240 14900 64280
rect 14379 63860 14421 63869
rect 14379 63820 14380 63860
rect 14420 63820 14421 63860
rect 14379 63811 14421 63820
rect 14476 63860 14516 63869
rect 14380 63726 14420 63811
rect 14476 63281 14516 63820
rect 14475 63272 14517 63281
rect 14475 63232 14476 63272
rect 14516 63232 14517 63272
rect 14475 63223 14517 63232
rect 14284 62476 14516 62516
rect 14380 62348 14420 62357
rect 14188 62308 14380 62348
rect 14092 62224 14228 62264
rect 14091 61760 14133 61769
rect 14091 61720 14092 61760
rect 14132 61720 14133 61760
rect 14091 61711 14133 61720
rect 14092 61601 14132 61711
rect 14091 61592 14133 61601
rect 14091 61552 14092 61592
rect 14132 61552 14133 61592
rect 14091 61543 14133 61552
rect 13995 59660 14037 59669
rect 13995 59620 13996 59660
rect 14036 59620 14037 59660
rect 13995 59611 14037 59620
rect 14092 59492 14132 61543
rect 13996 59452 14132 59492
rect 13996 59408 14036 59452
rect 13996 59359 14036 59368
rect 13996 57896 14036 57905
rect 13900 57856 13996 57896
rect 13996 57847 14036 57856
rect 13804 57772 13940 57812
rect 13900 57728 13940 57772
rect 13900 57688 14036 57728
rect 13708 57056 13748 57067
rect 13708 56981 13748 57016
rect 13804 57056 13844 57065
rect 13707 56972 13749 56981
rect 13707 56932 13708 56972
rect 13748 56932 13749 56972
rect 13707 56923 13749 56932
rect 13611 56720 13653 56729
rect 13611 56680 13612 56720
rect 13652 56680 13653 56720
rect 13804 56720 13844 57016
rect 13899 56720 13941 56729
rect 13804 56680 13900 56720
rect 13940 56680 13941 56720
rect 13611 56671 13653 56680
rect 13899 56671 13941 56680
rect 13420 56468 13460 56477
rect 13460 56428 13844 56468
rect 13420 56419 13460 56428
rect 13227 56384 13269 56393
rect 13227 56344 13228 56384
rect 13268 56344 13269 56384
rect 13227 56335 13269 56344
rect 13804 56384 13844 56428
rect 13804 56335 13844 56344
rect 13900 56384 13940 56671
rect 13900 56335 13940 56344
rect 13228 56250 13268 56335
rect 13996 56216 14036 57688
rect 14188 57308 14228 62224
rect 14380 60668 14420 62308
rect 14476 62348 14516 62476
rect 14476 60752 14516 62308
rect 14572 61769 14612 64240
rect 14667 63944 14709 63953
rect 14667 63904 14668 63944
rect 14708 63904 14709 63944
rect 14667 63895 14709 63904
rect 14571 61760 14613 61769
rect 14571 61720 14572 61760
rect 14612 61720 14613 61760
rect 14571 61711 14613 61720
rect 14572 61592 14612 61601
rect 14572 61433 14612 61552
rect 14571 61424 14613 61433
rect 14571 61384 14572 61424
rect 14612 61384 14613 61424
rect 14571 61375 14613 61384
rect 14571 61256 14613 61265
rect 14571 61216 14572 61256
rect 14612 61216 14613 61256
rect 14571 61207 14613 61216
rect 14572 60920 14612 61207
rect 14572 60871 14612 60880
rect 14476 60712 14612 60752
rect 14380 60628 14516 60668
rect 14283 60500 14325 60509
rect 14283 60460 14284 60500
rect 14324 60460 14325 60500
rect 14283 60451 14325 60460
rect 14284 60080 14324 60451
rect 14284 59753 14324 60040
rect 14283 59744 14325 59753
rect 14283 59704 14284 59744
rect 14324 59704 14325 59744
rect 14283 59695 14325 59704
rect 13900 56176 14036 56216
rect 14092 57268 14228 57308
rect 13707 56132 13749 56141
rect 13707 56092 13708 56132
rect 13748 56092 13749 56132
rect 13707 56083 13749 56092
rect 13228 55544 13268 55553
rect 12940 55420 13076 55460
rect 12940 54872 12980 54881
rect 12844 54832 12940 54872
rect 12748 54748 12884 54788
rect 12651 54032 12693 54041
rect 12651 53992 12652 54032
rect 12692 53992 12693 54032
rect 12651 53983 12693 53992
rect 12460 53488 12596 53528
rect 12652 53864 12692 53873
rect 12460 53285 12500 53488
rect 12652 53369 12692 53824
rect 12747 53528 12789 53537
rect 12747 53488 12748 53528
rect 12788 53488 12789 53528
rect 12747 53479 12789 53488
rect 12748 53394 12788 53479
rect 12556 53360 12596 53369
rect 12459 53276 12501 53285
rect 12459 53236 12460 53276
rect 12500 53236 12501 53276
rect 12459 53227 12501 53236
rect 12363 53108 12405 53117
rect 12363 53068 12364 53108
rect 12404 53068 12405 53108
rect 12363 53059 12405 53068
rect 12364 52949 12404 53059
rect 12363 52940 12405 52949
rect 12363 52900 12364 52940
rect 12404 52900 12405 52940
rect 12363 52891 12405 52900
rect 12556 52697 12596 53320
rect 12651 53360 12693 53369
rect 12651 53320 12652 53360
rect 12692 53320 12693 53360
rect 12651 53311 12693 53320
rect 12555 52688 12597 52697
rect 12555 52648 12556 52688
rect 12596 52648 12597 52688
rect 12555 52639 12597 52648
rect 12748 52613 12788 52644
rect 12747 52604 12789 52613
rect 12747 52564 12748 52604
rect 12788 52564 12789 52604
rect 12747 52555 12789 52564
rect 12460 52520 12500 52529
rect 12268 52480 12460 52520
rect 12460 52471 12500 52480
rect 12556 52520 12596 52529
rect 12556 52436 12596 52480
rect 12748 52520 12788 52555
rect 12748 52436 12788 52480
rect 12556 52396 12788 52436
rect 12267 52352 12309 52361
rect 12267 52312 12268 52352
rect 12308 52312 12309 52352
rect 12267 52303 12309 52312
rect 12268 52218 12308 52303
rect 12459 52100 12501 52109
rect 12748 52100 12788 52396
rect 12459 52060 12460 52100
rect 12500 52060 12501 52100
rect 12459 52051 12501 52060
rect 12652 52060 12788 52100
rect 12267 51176 12309 51185
rect 12267 51136 12268 51176
rect 12308 51136 12309 51176
rect 12267 51127 12309 51136
rect 12171 50336 12213 50345
rect 12171 50296 12172 50336
rect 12212 50296 12213 50336
rect 12171 50287 12213 50296
rect 12171 48320 12213 48329
rect 12171 48280 12172 48320
rect 12212 48280 12213 48320
rect 12171 48271 12213 48280
rect 12172 47321 12212 48271
rect 12171 47312 12213 47321
rect 12171 47272 12172 47312
rect 12212 47272 12213 47312
rect 12171 47263 12213 47272
rect 12172 47178 12212 47263
rect 12268 46640 12308 51127
rect 12363 50336 12405 50345
rect 12363 50296 12364 50336
rect 12404 50296 12405 50336
rect 12363 50287 12405 50296
rect 12460 50336 12500 52051
rect 12555 51848 12597 51857
rect 12555 51808 12556 51848
rect 12596 51808 12597 51848
rect 12555 51799 12597 51808
rect 12364 48077 12404 50287
rect 12460 48329 12500 50296
rect 12556 51008 12596 51799
rect 12652 51260 12692 52060
rect 12747 51848 12789 51857
rect 12747 51808 12748 51848
rect 12788 51808 12789 51848
rect 12747 51799 12789 51808
rect 12748 51714 12788 51799
rect 12748 51260 12788 51269
rect 12652 51220 12748 51260
rect 12748 51211 12788 51220
rect 12844 51008 12884 54748
rect 12940 54368 12980 54832
rect 13036 54452 13076 55420
rect 13228 54881 13268 55504
rect 13227 54872 13269 54881
rect 13227 54832 13228 54872
rect 13268 54832 13269 54872
rect 13227 54823 13269 54832
rect 13036 54412 13268 54452
rect 12940 54328 13172 54368
rect 12939 54200 12981 54209
rect 12939 54160 12940 54200
rect 12980 54160 12981 54200
rect 12939 54151 12981 54160
rect 12940 54051 12980 54151
rect 12940 54002 12980 54011
rect 13036 54032 13076 54041
rect 13036 53948 13076 53992
rect 12940 53908 13076 53948
rect 12940 53201 12980 53908
rect 13132 53864 13172 54328
rect 13036 53824 13172 53864
rect 12939 53192 12981 53201
rect 12939 53152 12940 53192
rect 12980 53152 12981 53192
rect 12939 53143 12981 53152
rect 12939 52940 12981 52949
rect 12939 52900 12940 52940
rect 12980 52900 12981 52940
rect 12939 52891 12981 52900
rect 12940 52688 12980 52891
rect 13036 52865 13076 53824
rect 13228 53537 13268 54412
rect 13420 54032 13460 54041
rect 13420 53696 13460 53992
rect 13516 54032 13556 54041
rect 13516 53873 13556 53992
rect 13515 53864 13557 53873
rect 13515 53824 13516 53864
rect 13556 53824 13557 53864
rect 13515 53815 13557 53824
rect 13420 53656 13556 53696
rect 13227 53528 13269 53537
rect 13227 53488 13228 53528
rect 13268 53488 13269 53528
rect 13227 53479 13269 53488
rect 13419 53528 13461 53537
rect 13419 53488 13420 53528
rect 13460 53488 13461 53528
rect 13419 53479 13461 53488
rect 13131 53360 13173 53369
rect 13131 53320 13132 53360
rect 13172 53320 13173 53360
rect 13131 53311 13173 53320
rect 13228 53360 13268 53371
rect 13132 53226 13172 53311
rect 13228 53285 13268 53320
rect 13227 53276 13269 53285
rect 13227 53236 13228 53276
rect 13268 53236 13269 53276
rect 13227 53227 13269 53236
rect 13131 53024 13173 53033
rect 13131 52984 13132 53024
rect 13172 52984 13173 53024
rect 13131 52975 13173 52984
rect 13035 52856 13077 52865
rect 13035 52816 13036 52856
rect 13076 52816 13077 52856
rect 13035 52807 13077 52816
rect 12940 52639 12980 52648
rect 12940 52520 12980 52529
rect 12940 52193 12980 52480
rect 13036 52520 13076 52531
rect 13036 52445 13076 52480
rect 13035 52436 13077 52445
rect 13035 52396 13036 52436
rect 13076 52396 13077 52436
rect 13035 52387 13077 52396
rect 12939 52184 12981 52193
rect 12939 52144 12940 52184
rect 12980 52144 12981 52184
rect 12939 52135 12981 52144
rect 12940 52016 12980 52135
rect 12940 51967 12980 51976
rect 13035 52016 13077 52025
rect 13035 51976 13036 52016
rect 13076 51976 13077 52016
rect 13035 51967 13077 51976
rect 13036 51764 13076 51967
rect 12459 48320 12501 48329
rect 12459 48280 12460 48320
rect 12500 48280 12501 48320
rect 12459 48271 12501 48280
rect 12556 48152 12596 50968
rect 12748 50968 12884 51008
rect 12940 51724 13076 51764
rect 12651 50420 12693 50429
rect 12651 50380 12652 50420
rect 12692 50380 12693 50420
rect 12651 50371 12693 50380
rect 12652 50286 12692 50371
rect 12748 49496 12788 50968
rect 12844 50084 12884 50093
rect 12844 49589 12884 50044
rect 12940 49673 12980 51724
rect 13035 51596 13077 51605
rect 13035 51556 13036 51596
rect 13076 51556 13077 51596
rect 13035 51547 13077 51556
rect 13036 50924 13076 51547
rect 13132 50924 13172 52975
rect 13227 52940 13269 52949
rect 13227 52900 13228 52940
rect 13268 52900 13269 52940
rect 13227 52891 13269 52900
rect 13228 52520 13268 52891
rect 13228 52471 13268 52480
rect 13324 52520 13364 52529
rect 13324 52361 13364 52480
rect 13323 52352 13365 52361
rect 13323 52312 13324 52352
rect 13364 52312 13365 52352
rect 13323 52303 13365 52312
rect 13324 51596 13364 51605
rect 13228 51556 13324 51596
rect 13228 51022 13268 51556
rect 13324 51547 13364 51556
rect 13420 51101 13460 53479
rect 13516 53444 13556 53656
rect 13611 53444 13653 53453
rect 13516 53404 13612 53444
rect 13652 53404 13653 53444
rect 13611 53395 13653 53404
rect 13612 53360 13652 53395
rect 13612 53309 13652 53320
rect 13708 53360 13748 56083
rect 13803 54032 13845 54041
rect 13803 53992 13804 54032
rect 13844 53992 13845 54032
rect 13803 53983 13845 53992
rect 13708 53311 13748 53320
rect 13712 52604 13754 52613
rect 13712 52564 13713 52604
rect 13753 52564 13754 52604
rect 13712 52555 13754 52564
rect 13516 52520 13556 52529
rect 13516 52193 13556 52480
rect 13611 52520 13653 52529
rect 13611 52480 13612 52520
rect 13652 52480 13653 52520
rect 13611 52471 13653 52480
rect 13713 52520 13753 52555
rect 13612 52386 13652 52471
rect 13713 52469 13753 52480
rect 13708 52352 13748 52361
rect 13515 52184 13557 52193
rect 13515 52144 13516 52184
rect 13556 52144 13557 52184
rect 13515 52135 13557 52144
rect 13515 52016 13557 52025
rect 13515 51976 13516 52016
rect 13556 51976 13557 52016
rect 13515 51967 13557 51976
rect 13516 51848 13556 51967
rect 13516 51799 13556 51808
rect 13708 51260 13748 52312
rect 13804 51521 13844 53983
rect 13803 51512 13845 51521
rect 13803 51472 13804 51512
rect 13844 51472 13845 51512
rect 13803 51463 13845 51472
rect 13612 51220 13748 51260
rect 13419 51092 13461 51101
rect 13419 51052 13420 51092
rect 13460 51052 13461 51092
rect 13419 51043 13461 51052
rect 13228 50973 13268 50982
rect 13132 50884 13556 50924
rect 13036 50875 13076 50884
rect 13227 50588 13269 50597
rect 13227 50548 13228 50588
rect 13268 50548 13269 50588
rect 13227 50539 13269 50548
rect 13036 50336 13076 50345
rect 13036 50261 13076 50296
rect 13035 50252 13077 50261
rect 13035 50212 13036 50252
rect 13076 50212 13077 50252
rect 13035 50203 13077 50212
rect 12939 49664 12981 49673
rect 12939 49624 12940 49664
rect 12980 49624 12981 49664
rect 12939 49615 12981 49624
rect 12843 49580 12885 49589
rect 12843 49540 12844 49580
rect 12884 49540 12885 49580
rect 12843 49531 12885 49540
rect 12940 49505 12980 49510
rect 12652 49456 12788 49496
rect 12939 49501 12981 49505
rect 12939 49456 12940 49501
rect 12980 49456 12981 49501
rect 12652 49160 12692 49456
rect 12939 49447 12981 49456
rect 12940 49366 12980 49447
rect 12748 49328 12788 49337
rect 12788 49288 12884 49328
rect 12748 49279 12788 49288
rect 12652 49120 12788 49160
rect 12460 48112 12596 48152
rect 12363 48068 12405 48077
rect 12363 48028 12364 48068
rect 12404 48028 12405 48068
rect 12363 48019 12405 48028
rect 12460 47993 12500 48112
rect 12459 47984 12501 47993
rect 12459 47944 12460 47984
rect 12500 47944 12501 47984
rect 12459 47935 12501 47944
rect 12556 47984 12596 47993
rect 12364 47480 12404 47489
rect 12556 47480 12596 47944
rect 12404 47440 12596 47480
rect 12652 47984 12692 47993
rect 12364 47431 12404 47440
rect 12556 47312 12596 47321
rect 12556 46901 12596 47272
rect 12555 46892 12597 46901
rect 12555 46852 12556 46892
rect 12596 46852 12597 46892
rect 12555 46843 12597 46852
rect 12172 46600 12308 46640
rect 12075 46472 12117 46481
rect 11884 46432 12020 46472
rect 11884 46304 11924 46313
rect 11691 45632 11733 45641
rect 11691 45592 11692 45632
rect 11732 45592 11733 45632
rect 11691 45583 11733 45592
rect 11787 44288 11829 44297
rect 11787 44248 11788 44288
rect 11828 44248 11829 44288
rect 11787 44239 11829 44248
rect 11788 44154 11828 44239
rect 11692 44036 11732 44045
rect 11595 43532 11637 43541
rect 11595 43492 11596 43532
rect 11636 43492 11637 43532
rect 11595 43483 11637 43492
rect 11499 41684 11541 41693
rect 11499 41644 11500 41684
rect 11540 41644 11541 41684
rect 11499 41635 11541 41644
rect 11596 41516 11636 43483
rect 11692 43205 11732 43996
rect 11691 43196 11733 43205
rect 11691 43156 11692 43196
rect 11732 43156 11733 43196
rect 11691 43147 11733 43156
rect 11787 41600 11829 41609
rect 11787 41560 11788 41600
rect 11828 41560 11829 41600
rect 11787 41551 11829 41560
rect 11500 41476 11636 41516
rect 11403 39920 11445 39929
rect 11403 39880 11404 39920
rect 11444 39880 11445 39920
rect 11403 39871 11445 39880
rect 11116 39836 11156 39845
rect 10924 39738 10964 39747
rect 10827 38492 10869 38501
rect 10827 38452 10828 38492
rect 10868 38452 10869 38492
rect 10827 38443 10869 38452
rect 10731 38408 10773 38417
rect 10731 38368 10732 38408
rect 10772 38368 10773 38408
rect 10731 38359 10773 38368
rect 10635 38156 10677 38165
rect 10635 38116 10636 38156
rect 10676 38116 10677 38156
rect 10635 38107 10677 38116
rect 10732 38156 10772 38165
rect 10636 38022 10676 38107
rect 10732 37997 10772 38116
rect 10731 37988 10773 37997
rect 10731 37948 10732 37988
rect 10772 37948 10773 37988
rect 10731 37939 10773 37948
rect 10636 37400 10676 37409
rect 10444 37360 10636 37400
rect 10347 36728 10389 36737
rect 10347 36688 10348 36728
rect 10388 36688 10389 36728
rect 10347 36679 10389 36688
rect 10059 36560 10101 36569
rect 10059 36520 10060 36560
rect 10100 36520 10101 36560
rect 10059 36511 10101 36520
rect 10060 36426 10100 36511
rect 10060 36056 10100 36065
rect 10060 35897 10100 36016
rect 10059 35888 10101 35897
rect 10059 35848 10060 35888
rect 10100 35848 10101 35888
rect 10059 35839 10101 35848
rect 10347 35720 10389 35729
rect 10347 35680 10348 35720
rect 10388 35680 10389 35720
rect 10347 35671 10389 35680
rect 10155 35552 10197 35561
rect 10155 35512 10156 35552
rect 10196 35512 10197 35552
rect 10155 35503 10197 35512
rect 10060 34964 10100 34973
rect 9963 34796 10005 34805
rect 9963 34756 9964 34796
rect 10004 34756 10005 34796
rect 9963 34747 10005 34756
rect 9964 34544 10004 34555
rect 9964 34469 10004 34504
rect 9963 34460 10005 34469
rect 9963 34420 9964 34460
rect 10004 34420 10005 34460
rect 9963 34411 10005 34420
rect 10060 34049 10100 34924
rect 10156 34133 10196 35503
rect 10251 35216 10293 35225
rect 10251 35176 10252 35216
rect 10292 35176 10293 35216
rect 10251 35167 10293 35176
rect 10348 35216 10388 35671
rect 10444 35216 10484 37360
rect 10636 37351 10676 37360
rect 10731 36896 10773 36905
rect 10731 36856 10732 36896
rect 10772 36856 10773 36896
rect 10731 36847 10773 36856
rect 10636 36728 10676 36737
rect 10539 35972 10581 35981
rect 10539 35932 10540 35972
rect 10580 35932 10581 35972
rect 10539 35923 10581 35932
rect 10540 35888 10580 35923
rect 10540 35837 10580 35848
rect 10540 35216 10580 35225
rect 10444 35176 10540 35216
rect 10348 35167 10388 35176
rect 10252 35082 10292 35167
rect 10443 34964 10485 34973
rect 10443 34924 10444 34964
rect 10484 34924 10485 34964
rect 10443 34915 10485 34924
rect 10347 34880 10389 34889
rect 10347 34840 10348 34880
rect 10388 34840 10389 34880
rect 10347 34831 10389 34840
rect 10251 34460 10293 34469
rect 10251 34420 10252 34460
rect 10292 34420 10293 34460
rect 10251 34411 10293 34420
rect 10252 34376 10292 34411
rect 10252 34325 10292 34336
rect 10348 34376 10388 34831
rect 10348 34327 10388 34336
rect 10155 34124 10197 34133
rect 10155 34084 10156 34124
rect 10196 34084 10292 34124
rect 10155 34075 10197 34084
rect 10059 34040 10101 34049
rect 10059 34000 10060 34040
rect 10100 34000 10101 34040
rect 10059 33991 10101 34000
rect 9868 33916 10004 33956
rect 9388 30892 9524 30932
rect 9196 28960 9332 29000
rect 9388 30764 9428 30773
rect 8907 28580 8949 28589
rect 8907 28540 8908 28580
rect 8948 28540 8949 28580
rect 8907 28531 8949 28540
rect 8852 26776 9044 26816
rect 8812 26767 8852 26776
rect 8716 25556 8756 26104
rect 8716 25516 8852 25556
rect 8715 25388 8757 25397
rect 8715 25348 8716 25388
rect 8756 25348 8763 25388
rect 8715 25339 8763 25348
rect 8723 25187 8763 25339
rect 8716 25178 8763 25187
rect 8756 25138 8763 25178
rect 8716 25096 8763 25138
rect 8812 25136 8852 25516
rect 8807 25096 8852 25136
rect 8807 25052 8847 25096
rect 8716 25012 8847 25052
rect 8619 24380 8661 24389
rect 8619 24340 8620 24380
rect 8660 24340 8661 24380
rect 8619 24331 8661 24340
rect 8620 24221 8660 24331
rect 8619 24212 8661 24221
rect 8619 24172 8620 24212
rect 8660 24172 8661 24212
rect 8619 24163 8661 24172
rect 8716 23288 8756 25012
rect 8908 24632 8948 24641
rect 9004 24632 9044 26776
rect 9099 26480 9141 26489
rect 9099 26440 9100 26480
rect 9140 26440 9141 26480
rect 9099 26431 9141 26440
rect 8620 23248 8756 23288
rect 8812 24592 8908 24632
rect 8948 24592 9044 24632
rect 8523 23120 8565 23129
rect 8523 23080 8524 23120
rect 8564 23080 8565 23120
rect 8523 23071 8565 23080
rect 8523 22952 8565 22961
rect 8523 22912 8524 22952
rect 8564 22912 8565 22952
rect 8523 22903 8565 22912
rect 8331 21944 8373 21953
rect 8331 21904 8332 21944
rect 8372 21904 8373 21944
rect 8331 21895 8373 21904
rect 7892 21400 8276 21440
rect 7852 21391 7892 21400
rect 7851 21188 7893 21197
rect 7851 21148 7852 21188
rect 7892 21148 7893 21188
rect 7851 21139 7893 21148
rect 7852 20096 7892 21139
rect 8524 20945 8564 22903
rect 8331 20936 8373 20945
rect 8331 20896 8332 20936
rect 8372 20896 8373 20936
rect 8331 20887 8373 20896
rect 8523 20936 8565 20945
rect 8523 20896 8524 20936
rect 8564 20896 8565 20936
rect 8523 20887 8565 20896
rect 8332 20768 8372 20887
rect 8332 20719 8372 20728
rect 8620 20609 8660 23248
rect 8715 23120 8757 23129
rect 8715 23080 8716 23120
rect 8756 23080 8757 23120
rect 8715 23071 8757 23080
rect 8716 21197 8756 23071
rect 8812 21869 8852 24592
rect 8908 24583 8948 24592
rect 9004 23129 9044 23214
rect 8908 23120 8948 23129
rect 8908 22625 8948 23080
rect 9003 23120 9045 23129
rect 9003 23080 9004 23120
rect 9044 23080 9045 23120
rect 9100 23120 9140 26431
rect 9196 24053 9236 28960
rect 9388 28841 9428 30724
rect 9484 30269 9524 30892
rect 9483 30260 9525 30269
rect 9483 30220 9484 30260
rect 9524 30220 9525 30260
rect 9483 30211 9525 30220
rect 9580 29000 9620 33328
rect 9676 32192 9716 32203
rect 9676 32117 9716 32152
rect 9675 32108 9717 32117
rect 9675 32068 9676 32108
rect 9716 32068 9717 32108
rect 9675 32059 9717 32068
rect 9484 28960 9620 29000
rect 9387 28832 9429 28841
rect 9387 28792 9388 28832
rect 9428 28792 9429 28832
rect 9387 28783 9429 28792
rect 9292 26821 9332 26830
rect 9484 26816 9524 28960
rect 9292 26321 9332 26781
rect 9388 26776 9524 26816
rect 9676 27656 9716 27665
rect 9291 26312 9333 26321
rect 9291 26272 9292 26312
rect 9332 26272 9333 26312
rect 9291 26263 9333 26272
rect 9388 24716 9428 26776
rect 9292 24676 9428 24716
rect 9484 26648 9524 26657
rect 9195 24044 9237 24053
rect 9195 24004 9196 24044
rect 9236 24004 9237 24044
rect 9195 23995 9237 24004
rect 9292 23969 9332 24676
rect 9388 24618 9428 24627
rect 9388 24044 9428 24578
rect 9388 23995 9428 24004
rect 9291 23960 9333 23969
rect 9291 23920 9292 23960
rect 9332 23920 9333 23960
rect 9291 23911 9333 23920
rect 9195 23876 9237 23885
rect 9195 23836 9196 23876
rect 9236 23836 9237 23876
rect 9195 23827 9237 23836
rect 9196 23792 9236 23827
rect 9196 23741 9236 23752
rect 9484 23633 9524 26608
rect 9580 24716 9620 24725
rect 9580 23969 9620 24676
rect 9579 23960 9621 23969
rect 9579 23920 9580 23960
rect 9620 23920 9621 23960
rect 9579 23911 9621 23920
rect 9676 23885 9716 27616
rect 9772 24137 9812 33832
rect 9867 32360 9909 32369
rect 9867 32320 9868 32360
rect 9908 32320 9909 32360
rect 9867 32311 9909 32320
rect 9868 32226 9908 32311
rect 9867 28496 9909 28505
rect 9867 28456 9868 28496
rect 9908 28456 9909 28496
rect 9867 28447 9909 28456
rect 9868 27740 9908 28447
rect 9868 27691 9908 27700
rect 9964 26480 10004 33916
rect 10060 32864 10100 32873
rect 10060 32369 10100 32824
rect 10155 32864 10197 32873
rect 10155 32824 10156 32864
rect 10196 32824 10197 32864
rect 10155 32815 10197 32824
rect 10156 32730 10196 32815
rect 10059 32360 10101 32369
rect 10059 32320 10060 32360
rect 10100 32320 10101 32360
rect 10059 32311 10101 32320
rect 10156 32192 10196 32201
rect 10252 32192 10292 34084
rect 10347 33956 10389 33965
rect 10347 33916 10348 33956
rect 10388 33916 10389 33956
rect 10347 33907 10389 33916
rect 10060 32152 10156 32192
rect 10196 32152 10292 32192
rect 10060 27413 10100 32152
rect 10156 32143 10196 32152
rect 10348 32108 10388 33907
rect 10444 32948 10484 34915
rect 10540 33545 10580 35176
rect 10636 34469 10676 36688
rect 10732 35477 10772 36847
rect 10828 36728 10868 38443
rect 10924 37661 10964 39698
rect 11020 38912 11060 38921
rect 10923 37652 10965 37661
rect 10923 37612 10924 37652
rect 10964 37612 10965 37652
rect 10923 37603 10965 37612
rect 11020 36905 11060 38872
rect 11019 36896 11061 36905
rect 11019 36856 11020 36896
rect 11060 36856 11061 36896
rect 11019 36847 11061 36856
rect 10924 36728 10964 36737
rect 10828 36688 10924 36728
rect 10924 36679 10964 36688
rect 11019 36728 11061 36737
rect 11019 36688 11020 36728
rect 11060 36688 11061 36728
rect 11019 36679 11061 36688
rect 10923 36560 10965 36569
rect 10923 36520 10924 36560
rect 10964 36520 10965 36560
rect 10923 36511 10965 36520
rect 10731 35468 10773 35477
rect 10731 35428 10732 35468
rect 10772 35428 10773 35468
rect 10731 35419 10773 35428
rect 10732 34889 10772 35419
rect 10731 34880 10773 34889
rect 10731 34840 10732 34880
rect 10772 34840 10773 34880
rect 10731 34831 10773 34840
rect 10635 34460 10677 34469
rect 10635 34420 10636 34460
rect 10676 34420 10677 34460
rect 10635 34411 10677 34420
rect 10731 34376 10773 34385
rect 10731 34336 10732 34376
rect 10772 34336 10773 34376
rect 10731 34327 10773 34336
rect 10828 34376 10868 34385
rect 10732 34242 10772 34327
rect 10635 34208 10677 34217
rect 10635 34168 10636 34208
rect 10676 34168 10677 34208
rect 10635 34159 10677 34168
rect 10539 33536 10581 33545
rect 10539 33496 10540 33536
rect 10580 33496 10581 33536
rect 10539 33487 10581 33496
rect 10636 32957 10676 34159
rect 10828 33872 10868 34336
rect 10732 33832 10868 33872
rect 10732 33629 10772 33832
rect 10827 33704 10869 33713
rect 10827 33664 10828 33704
rect 10868 33664 10869 33704
rect 10827 33655 10869 33664
rect 10731 33620 10773 33629
rect 10731 33580 10732 33620
rect 10772 33580 10773 33620
rect 10731 33571 10773 33580
rect 10540 32948 10580 32957
rect 10444 32908 10540 32948
rect 10540 32899 10580 32908
rect 10635 32948 10677 32957
rect 10635 32908 10636 32948
rect 10676 32908 10677 32948
rect 10635 32899 10677 32908
rect 10636 32814 10676 32899
rect 10731 32864 10773 32873
rect 10731 32824 10732 32864
rect 10772 32824 10773 32864
rect 10731 32815 10773 32824
rect 10252 32068 10388 32108
rect 10155 31352 10197 31361
rect 10155 31312 10156 31352
rect 10196 31312 10197 31352
rect 10155 31303 10197 31312
rect 10156 31218 10196 31303
rect 10252 31100 10292 32068
rect 10636 31352 10676 31361
rect 10348 31268 10388 31277
rect 10636 31268 10676 31312
rect 10388 31228 10676 31268
rect 10732 31352 10772 32815
rect 10828 32696 10868 33655
rect 10924 33041 10964 36511
rect 10923 33032 10965 33041
rect 10923 32992 10924 33032
rect 10964 32992 10965 33032
rect 10923 32983 10965 32992
rect 10924 32873 10964 32983
rect 10923 32864 10965 32873
rect 10923 32824 10924 32864
rect 10964 32824 10965 32864
rect 10923 32815 10965 32824
rect 11020 32789 11060 36679
rect 11116 32864 11156 39796
rect 11211 38240 11253 38249
rect 11211 38200 11212 38240
rect 11252 38200 11253 38240
rect 11211 38191 11253 38200
rect 11212 38106 11252 38191
rect 11500 37820 11540 41476
rect 11788 41432 11828 41551
rect 11595 41348 11637 41357
rect 11595 41308 11596 41348
rect 11636 41308 11637 41348
rect 11595 41299 11637 41308
rect 11404 37780 11540 37820
rect 11211 37148 11253 37157
rect 11211 37108 11212 37148
rect 11252 37108 11253 37148
rect 11211 37099 11253 37108
rect 11212 34805 11252 37099
rect 11307 36476 11349 36485
rect 11307 36436 11308 36476
rect 11348 36436 11349 36476
rect 11307 36427 11349 36436
rect 11308 36342 11348 36427
rect 11307 36224 11349 36233
rect 11307 36184 11308 36224
rect 11348 36184 11349 36224
rect 11307 36175 11349 36184
rect 11308 35804 11348 36175
rect 11404 35981 11444 37780
rect 11499 36812 11541 36821
rect 11499 36772 11500 36812
rect 11540 36772 11541 36812
rect 11499 36763 11541 36772
rect 11500 36728 11540 36763
rect 11500 36653 11540 36688
rect 11499 36644 11541 36653
rect 11499 36604 11500 36644
rect 11540 36604 11541 36644
rect 11499 36595 11541 36604
rect 11499 36476 11541 36485
rect 11499 36436 11500 36476
rect 11540 36436 11541 36476
rect 11499 36427 11541 36436
rect 11403 35972 11445 35981
rect 11403 35932 11404 35972
rect 11444 35932 11445 35972
rect 11403 35923 11445 35932
rect 11308 35764 11444 35804
rect 11211 34796 11253 34805
rect 11211 34756 11212 34796
rect 11252 34756 11253 34796
rect 11211 34747 11253 34756
rect 11404 34553 11444 35764
rect 11500 35561 11540 36427
rect 11499 35552 11541 35561
rect 11499 35512 11500 35552
rect 11540 35512 11541 35552
rect 11499 35503 11541 35512
rect 11403 34544 11445 34553
rect 11403 34504 11404 34544
rect 11444 34504 11445 34544
rect 11403 34495 11445 34504
rect 11308 34376 11348 34385
rect 11212 34336 11308 34376
rect 11212 34217 11252 34336
rect 11308 34327 11348 34336
rect 11211 34208 11253 34217
rect 11211 34168 11212 34208
rect 11252 34168 11253 34208
rect 11211 34159 11253 34168
rect 11403 33872 11445 33881
rect 11403 33832 11404 33872
rect 11444 33832 11445 33872
rect 11403 33823 11445 33832
rect 11211 32948 11253 32957
rect 11211 32908 11212 32948
rect 11252 32908 11253 32948
rect 11211 32899 11253 32908
rect 11019 32780 11061 32789
rect 11019 32740 11020 32780
rect 11060 32740 11061 32780
rect 11019 32731 11061 32740
rect 10828 32656 10964 32696
rect 10348 31219 10388 31228
rect 10156 31060 10292 31100
rect 10156 28328 10196 31060
rect 10732 30848 10772 31312
rect 10444 30808 10772 30848
rect 10347 29840 10389 29849
rect 10347 29800 10348 29840
rect 10388 29800 10389 29840
rect 10347 29791 10389 29800
rect 10348 29706 10388 29791
rect 10252 29168 10292 29177
rect 10252 28505 10292 29128
rect 10348 29168 10388 29177
rect 10444 29168 10484 30808
rect 10636 30680 10676 30689
rect 10540 30092 10580 30101
rect 10636 30092 10676 30640
rect 10732 30680 10772 30808
rect 10732 30631 10772 30640
rect 10827 30680 10869 30689
rect 10827 30640 10828 30680
rect 10868 30640 10869 30680
rect 10827 30631 10869 30640
rect 10580 30052 10676 30092
rect 10540 30043 10580 30052
rect 10539 29924 10581 29933
rect 10539 29884 10540 29924
rect 10580 29884 10581 29924
rect 10539 29875 10581 29884
rect 10388 29128 10484 29168
rect 10348 29119 10388 29128
rect 10444 29000 10484 29128
rect 10348 28960 10484 29000
rect 10251 28496 10293 28505
rect 10251 28456 10252 28496
rect 10292 28456 10293 28496
rect 10251 28447 10293 28456
rect 10251 28328 10293 28337
rect 10156 28288 10252 28328
rect 10292 28288 10293 28328
rect 10251 28279 10293 28288
rect 10252 28194 10292 28279
rect 10156 27656 10196 27665
rect 10059 27404 10101 27413
rect 10059 27364 10060 27404
rect 10100 27364 10101 27404
rect 10059 27355 10101 27364
rect 10059 27236 10101 27245
rect 10059 27196 10060 27236
rect 10100 27196 10101 27236
rect 10059 27187 10101 27196
rect 10060 26816 10100 27187
rect 10060 26767 10100 26776
rect 9964 26440 10100 26480
rect 9963 26144 10005 26153
rect 9963 26104 9964 26144
rect 10004 26104 10005 26144
rect 9963 26095 10005 26104
rect 9964 26010 10004 26095
rect 9964 24632 10004 24641
rect 10060 24632 10100 26440
rect 10156 26312 10196 27616
rect 10156 26263 10196 26272
rect 10252 27656 10292 27665
rect 10348 27656 10388 28960
rect 10443 28328 10485 28337
rect 10443 28288 10444 28328
rect 10484 28288 10485 28328
rect 10443 28279 10485 28288
rect 10292 27616 10388 27656
rect 10004 24592 10100 24632
rect 10156 25304 10196 25313
rect 9964 24473 10004 24592
rect 9963 24464 10005 24473
rect 9963 24424 9964 24464
rect 10004 24424 10005 24464
rect 9963 24415 10005 24424
rect 9771 24128 9813 24137
rect 9771 24088 9772 24128
rect 9812 24088 9813 24128
rect 9771 24079 9813 24088
rect 10156 23969 10196 25264
rect 9963 23960 10005 23969
rect 9963 23920 9964 23960
rect 10004 23920 10005 23960
rect 9963 23911 10005 23920
rect 10155 23960 10197 23969
rect 10155 23920 10156 23960
rect 10196 23920 10197 23960
rect 10155 23911 10197 23920
rect 9675 23876 9717 23885
rect 9675 23836 9676 23876
rect 9716 23836 9812 23876
rect 9675 23827 9717 23836
rect 9772 23792 9812 23836
rect 9812 23752 9908 23792
rect 9772 23743 9812 23752
rect 9675 23708 9717 23717
rect 9675 23668 9676 23708
rect 9716 23668 9717 23708
rect 9675 23659 9717 23668
rect 9483 23624 9525 23633
rect 9483 23584 9484 23624
rect 9524 23584 9525 23624
rect 9483 23575 9525 23584
rect 9580 23624 9620 23633
rect 9580 23465 9620 23584
rect 9579 23456 9621 23465
rect 9579 23416 9580 23456
rect 9620 23416 9621 23456
rect 9579 23407 9621 23416
rect 9387 23372 9429 23381
rect 9387 23332 9388 23372
rect 9428 23332 9429 23372
rect 9387 23323 9429 23332
rect 9291 23288 9333 23297
rect 9291 23248 9292 23288
rect 9332 23248 9333 23288
rect 9291 23239 9333 23248
rect 9292 23154 9332 23239
rect 9196 23120 9236 23129
rect 9100 23080 9196 23120
rect 9003 23071 9045 23080
rect 9196 23036 9236 23080
rect 9388 23120 9428 23323
rect 9676 23288 9716 23659
rect 9388 23071 9428 23080
rect 9484 23248 9676 23288
rect 9484 23120 9524 23248
rect 9676 23239 9716 23248
rect 9484 23071 9524 23080
rect 9771 23120 9813 23129
rect 9771 23080 9772 23120
rect 9812 23080 9813 23120
rect 9771 23071 9813 23080
rect 9868 23120 9908 23752
rect 9196 22996 9332 23036
rect 9004 22952 9044 22961
rect 9044 22912 9243 22952
rect 9004 22903 9044 22912
rect 9203 22868 9243 22912
rect 9196 22828 9243 22868
rect 8907 22616 8949 22625
rect 8907 22576 8908 22616
rect 8948 22576 8949 22616
rect 8907 22567 8949 22576
rect 9196 22541 9236 22828
rect 9195 22532 9237 22541
rect 9195 22492 9196 22532
rect 9236 22492 9237 22532
rect 9195 22483 9237 22492
rect 9292 22364 9332 22996
rect 9387 22868 9429 22877
rect 9387 22828 9388 22868
rect 9428 22828 9429 22868
rect 9387 22819 9429 22828
rect 9196 22324 9332 22364
rect 8811 21860 8853 21869
rect 8811 21820 8812 21860
rect 8852 21820 8853 21860
rect 8811 21811 8853 21820
rect 9196 21440 9236 22324
rect 9388 22280 9428 22819
rect 9772 22700 9812 23071
rect 9868 22877 9908 23080
rect 9867 22868 9909 22877
rect 9867 22828 9868 22868
rect 9908 22828 9909 22868
rect 9867 22819 9909 22828
rect 9772 22660 9908 22700
rect 9579 22616 9621 22625
rect 9579 22576 9580 22616
rect 9620 22576 9621 22616
rect 9579 22567 9621 22576
rect 9580 22532 9620 22567
rect 9580 22481 9620 22492
rect 9771 22532 9813 22541
rect 9771 22492 9772 22532
rect 9812 22492 9813 22532
rect 9771 22483 9813 22492
rect 9292 21608 9332 21617
rect 9388 21608 9428 22240
rect 9483 22280 9525 22289
rect 9483 22240 9484 22280
rect 9524 22240 9525 22280
rect 9483 22231 9525 22240
rect 9772 22280 9812 22483
rect 9868 22289 9908 22660
rect 9772 22231 9812 22240
rect 9867 22280 9909 22289
rect 9867 22240 9868 22280
rect 9908 22240 9909 22280
rect 9867 22231 9909 22240
rect 9484 21776 9524 22231
rect 9964 22112 10004 23911
rect 10155 22616 10197 22625
rect 10155 22576 10156 22616
rect 10196 22576 10197 22616
rect 10155 22567 10197 22576
rect 9484 21727 9524 21736
rect 9868 22072 10004 22112
rect 10060 22280 10100 22289
rect 9675 21692 9717 21701
rect 9675 21652 9676 21692
rect 9716 21652 9717 21692
rect 9675 21643 9717 21652
rect 9676 21608 9716 21643
rect 9332 21568 9524 21608
rect 9292 21559 9332 21568
rect 9196 21400 9332 21440
rect 8715 21188 8757 21197
rect 8715 21148 8716 21188
rect 8756 21148 8757 21188
rect 8715 21139 8757 21148
rect 9195 21188 9237 21197
rect 9195 21148 9196 21188
rect 9236 21148 9237 21188
rect 9195 21139 9237 21148
rect 8524 20600 8564 20609
rect 8524 20273 8564 20560
rect 8619 20600 8661 20609
rect 8619 20560 8620 20600
rect 8660 20560 8661 20600
rect 8619 20551 8661 20560
rect 8620 20441 8660 20551
rect 8619 20432 8661 20441
rect 8619 20392 8620 20432
rect 8660 20392 8661 20432
rect 8619 20383 8661 20392
rect 7947 20264 7989 20273
rect 8523 20264 8565 20273
rect 7947 20224 7948 20264
rect 7988 20224 7989 20264
rect 7947 20215 7989 20224
rect 8236 20224 8468 20264
rect 7852 18257 7892 20056
rect 7948 18677 7988 20215
rect 8043 20096 8085 20105
rect 8043 20056 8044 20096
rect 8084 20056 8085 20096
rect 8043 20047 8085 20056
rect 8140 20096 8180 20105
rect 8236 20096 8276 20224
rect 8180 20056 8276 20096
rect 8140 20047 8180 20056
rect 8044 19676 8084 20047
rect 8139 19928 8181 19937
rect 8139 19888 8140 19928
rect 8180 19888 8181 19928
rect 8139 19879 8181 19888
rect 8140 19794 8180 19879
rect 8044 19636 8180 19676
rect 8044 19349 8084 19380
rect 8043 19340 8085 19349
rect 8043 19300 8044 19340
rect 8084 19300 8085 19340
rect 8043 19291 8085 19300
rect 8044 19256 8084 19291
rect 7947 18668 7989 18677
rect 7947 18628 7948 18668
rect 7988 18628 7989 18668
rect 7947 18619 7989 18628
rect 8044 18584 8084 19216
rect 8140 18752 8180 19636
rect 8236 19508 8276 20056
rect 8332 20096 8372 20107
rect 8332 20021 8372 20056
rect 8428 20096 8468 20224
rect 8523 20224 8524 20264
rect 8564 20224 8565 20264
rect 8523 20215 8565 20224
rect 8812 20264 8852 20273
rect 8852 20224 9044 20264
rect 8812 20215 8852 20224
rect 8716 20096 8756 20105
rect 8428 20047 8468 20056
rect 8572 20081 8612 20090
rect 8331 20012 8373 20021
rect 8331 19972 8332 20012
rect 8372 19972 8373 20012
rect 8331 19963 8373 19972
rect 8572 19937 8612 20041
rect 8709 20056 8716 20081
rect 8709 20041 8756 20056
rect 8873 20081 8913 20090
rect 8913 20041 8948 20081
rect 8709 20021 8749 20041
rect 8873 20032 8948 20041
rect 8667 20012 8749 20021
rect 8667 19972 8668 20012
rect 8708 19972 8749 20012
rect 8667 19963 8709 19972
rect 8571 19928 8613 19937
rect 8571 19888 8572 19928
rect 8612 19888 8613 19928
rect 8571 19879 8613 19888
rect 8811 19760 8853 19769
rect 8811 19720 8812 19760
rect 8852 19720 8853 19760
rect 8811 19711 8853 19720
rect 8236 19459 8276 19468
rect 8812 19256 8852 19711
rect 8908 19685 8948 20032
rect 8907 19676 8949 19685
rect 8907 19636 8908 19676
rect 8948 19636 8949 19676
rect 8907 19627 8949 19636
rect 8812 19207 8852 19216
rect 8331 19088 8373 19097
rect 8331 19048 8332 19088
rect 8372 19048 8373 19088
rect 8331 19039 8373 19048
rect 8236 18752 8276 18761
rect 8140 18712 8236 18752
rect 8236 18703 8276 18712
rect 8084 18544 8276 18584
rect 8044 18535 8084 18544
rect 7947 18416 7989 18425
rect 7947 18376 7948 18416
rect 7988 18376 7989 18416
rect 7947 18367 7989 18376
rect 7851 18248 7893 18257
rect 7851 18208 7852 18248
rect 7892 18208 7893 18248
rect 7851 18199 7893 18208
rect 7755 17912 7797 17921
rect 7755 17872 7756 17912
rect 7796 17872 7797 17912
rect 7755 17863 7797 17872
rect 7700 17704 7796 17744
rect 7660 17695 7700 17704
rect 7563 17576 7605 17585
rect 7563 17536 7564 17576
rect 7604 17536 7605 17576
rect 7563 17527 7605 17536
rect 7467 17408 7509 17417
rect 7467 17368 7468 17408
rect 7508 17368 7509 17408
rect 7467 17359 7509 17368
rect 6988 17032 7084 17072
rect 6891 16736 6933 16745
rect 6891 16696 6892 16736
rect 6932 16696 6933 16736
rect 6891 16687 6933 16696
rect 6988 16409 7028 17032
rect 7084 17023 7124 17032
rect 7180 17284 7412 17324
rect 7083 16736 7125 16745
rect 7083 16696 7084 16736
rect 7124 16696 7125 16736
rect 7083 16687 7125 16696
rect 6987 16400 7029 16409
rect 6987 16360 6988 16400
rect 7028 16360 7029 16400
rect 6987 16351 7029 16360
rect 6796 16232 6836 16241
rect 6988 16232 7028 16351
rect 6836 16192 7028 16232
rect 6796 16183 6836 16192
rect 6988 16064 7028 16073
rect 6700 16024 6836 16064
rect 6603 14972 6645 14981
rect 6603 14932 6604 14972
rect 6644 14932 6645 14972
rect 6603 14923 6645 14932
rect 6604 14048 6644 14923
rect 6700 14720 6740 14729
rect 6700 14057 6740 14680
rect 6796 14393 6836 16024
rect 6892 16024 6988 16064
rect 6892 15560 6932 16024
rect 6988 16015 7028 16024
rect 6892 15511 6932 15520
rect 6987 15560 7029 15569
rect 6987 15520 6988 15560
rect 7028 15520 7029 15560
rect 6987 15511 7029 15520
rect 6988 15233 7028 15511
rect 6987 15224 7029 15233
rect 6987 15184 6988 15224
rect 7028 15184 7029 15224
rect 6987 15175 7029 15184
rect 6795 14384 6837 14393
rect 6795 14344 6796 14384
rect 6836 14344 6837 14384
rect 6795 14335 6837 14344
rect 6795 14132 6837 14141
rect 6795 14092 6796 14132
rect 6836 14092 6837 14132
rect 6795 14083 6837 14092
rect 6604 13889 6644 14008
rect 6699 14048 6741 14057
rect 6699 14008 6700 14048
rect 6740 14008 6741 14048
rect 6699 13999 6741 14008
rect 6603 13880 6645 13889
rect 6603 13840 6604 13880
rect 6644 13840 6645 13880
rect 6603 13831 6645 13840
rect 6699 13544 6741 13553
rect 6699 13504 6700 13544
rect 6740 13504 6741 13544
rect 6699 13495 6741 13504
rect 6700 13222 6740 13495
rect 6507 13208 6549 13217
rect 6507 13168 6508 13208
rect 6548 13168 6549 13208
rect 6700 13173 6740 13182
rect 6507 13159 6549 13168
rect 6411 12872 6453 12881
rect 6411 12832 6412 12872
rect 6452 12832 6453 12872
rect 6411 12823 6453 12832
rect 6412 12536 6452 12545
rect 6452 12496 6548 12536
rect 6412 12487 6452 12496
rect 6124 12076 6260 12116
rect 6124 11537 6164 12076
rect 6219 11948 6261 11957
rect 6219 11908 6220 11948
rect 6260 11908 6261 11948
rect 6219 11899 6261 11908
rect 6411 11948 6453 11957
rect 6411 11908 6412 11948
rect 6452 11908 6453 11948
rect 6411 11899 6453 11908
rect 6220 11696 6260 11899
rect 6412 11814 6452 11899
rect 6123 11528 6165 11537
rect 6123 11488 6124 11528
rect 6164 11488 6165 11528
rect 6123 11479 6165 11488
rect 6220 11453 6260 11656
rect 6219 11444 6261 11453
rect 6219 11404 6220 11444
rect 6260 11404 6261 11444
rect 6219 11395 6261 11404
rect 6508 11201 6548 12496
rect 6604 12368 6644 12377
rect 6604 11705 6644 12328
rect 6796 11948 6836 14083
rect 6987 13880 7029 13889
rect 6987 13840 6988 13880
rect 7028 13840 7029 13880
rect 6987 13831 7029 13840
rect 6891 13124 6933 13133
rect 6891 13084 6892 13124
rect 6932 13084 6933 13124
rect 6891 13075 6933 13084
rect 6892 12990 6932 13075
rect 6988 12620 7028 13831
rect 7084 13292 7124 16687
rect 7180 14384 7220 17284
rect 7276 17156 7316 17165
rect 7316 17116 7604 17156
rect 7276 17107 7316 17116
rect 7564 17072 7604 17116
rect 7564 17023 7604 17032
rect 7659 17072 7701 17081
rect 7659 17032 7660 17072
rect 7700 17032 7701 17072
rect 7659 17023 7701 17032
rect 7660 16938 7700 17023
rect 7659 16736 7701 16745
rect 7659 16696 7660 16736
rect 7700 16696 7701 16736
rect 7659 16687 7701 16696
rect 7563 16568 7605 16577
rect 7563 16528 7564 16568
rect 7604 16528 7605 16568
rect 7563 16519 7605 16528
rect 7275 16400 7317 16409
rect 7275 16360 7276 16400
rect 7316 16360 7317 16400
rect 7275 16351 7317 16360
rect 7276 14729 7316 16351
rect 7372 15476 7412 15485
rect 7372 15317 7412 15436
rect 7467 15476 7509 15485
rect 7467 15436 7468 15476
rect 7508 15436 7509 15476
rect 7467 15427 7509 15436
rect 7468 15342 7508 15427
rect 7371 15308 7413 15317
rect 7371 15268 7372 15308
rect 7412 15268 7413 15308
rect 7371 15259 7413 15268
rect 7564 15224 7604 16519
rect 7468 15184 7604 15224
rect 7660 16232 7700 16687
rect 7275 14720 7317 14729
rect 7275 14680 7276 14720
rect 7316 14680 7317 14720
rect 7275 14671 7317 14680
rect 7180 14344 7316 14384
rect 7179 14216 7221 14225
rect 7179 14176 7180 14216
rect 7220 14176 7221 14216
rect 7179 14167 7221 14176
rect 7180 13460 7220 14167
rect 7180 13411 7220 13420
rect 7084 13252 7220 13292
rect 7084 13197 7124 13206
rect 7084 13133 7124 13157
rect 7083 13124 7125 13133
rect 7083 13084 7084 13124
rect 7124 13084 7125 13124
rect 7083 13075 7125 13084
rect 7084 13062 7124 13075
rect 7180 12965 7220 13252
rect 7179 12956 7221 12965
rect 7179 12916 7180 12956
rect 7220 12916 7221 12956
rect 7179 12907 7221 12916
rect 7083 12872 7125 12881
rect 7083 12832 7084 12872
rect 7124 12832 7125 12872
rect 7083 12823 7125 12832
rect 6988 12571 7028 12580
rect 6892 11948 6932 11957
rect 6796 11908 6892 11948
rect 6892 11899 6932 11908
rect 6603 11696 6645 11705
rect 6603 11656 6604 11696
rect 6644 11656 6645 11696
rect 6603 11647 6645 11656
rect 6891 11696 6933 11705
rect 6891 11656 6892 11696
rect 6932 11656 6933 11696
rect 6891 11647 6933 11656
rect 7084 11696 7124 12823
rect 7276 12704 7316 14344
rect 7371 13040 7413 13049
rect 7371 13000 7372 13040
rect 7412 13000 7413 13040
rect 7371 12991 7413 13000
rect 7372 12906 7412 12991
rect 7468 12881 7508 15184
rect 7563 15056 7605 15065
rect 7563 15016 7564 15056
rect 7604 15016 7605 15056
rect 7563 15007 7605 15016
rect 7564 13208 7604 15007
rect 7660 13712 7700 16192
rect 7756 14309 7796 17704
rect 7851 16820 7893 16829
rect 7851 16780 7852 16820
rect 7892 16780 7893 16820
rect 7851 16771 7893 16780
rect 7755 14300 7797 14309
rect 7755 14260 7756 14300
rect 7796 14260 7797 14300
rect 7755 14251 7797 14260
rect 7852 14048 7892 16771
rect 7948 15560 7988 18367
rect 8139 17912 8181 17921
rect 8139 17872 8140 17912
rect 8180 17872 8181 17912
rect 8139 17863 8181 17872
rect 8140 17744 8180 17863
rect 8140 17695 8180 17704
rect 8043 17576 8085 17585
rect 8043 17536 8044 17576
rect 8084 17536 8085 17576
rect 8043 17527 8085 17536
rect 7948 15401 7988 15520
rect 8044 16988 8084 17527
rect 8139 17408 8181 17417
rect 8139 17368 8140 17408
rect 8180 17368 8181 17408
rect 8139 17359 8181 17368
rect 7947 15392 7989 15401
rect 7947 15352 7948 15392
rect 7988 15352 7989 15392
rect 7947 15343 7989 15352
rect 8044 15149 8084 16948
rect 8140 16988 8180 17359
rect 8140 16829 8180 16948
rect 8139 16820 8181 16829
rect 8139 16780 8140 16820
rect 8180 16780 8181 16820
rect 8139 16771 8181 16780
rect 8236 15821 8276 18544
rect 8332 16241 8372 19039
rect 8619 18668 8661 18677
rect 8619 18628 8620 18668
rect 8660 18628 8661 18668
rect 8619 18619 8661 18628
rect 8427 18164 8469 18173
rect 8427 18124 8428 18164
rect 8468 18124 8469 18164
rect 8427 18115 8469 18124
rect 8428 17669 8468 18115
rect 8523 17912 8565 17921
rect 8523 17872 8524 17912
rect 8564 17872 8565 17912
rect 8523 17863 8565 17872
rect 8427 17660 8469 17669
rect 8427 17620 8428 17660
rect 8468 17620 8469 17660
rect 8427 17611 8469 17620
rect 8524 17072 8564 17863
rect 8620 17758 8660 18619
rect 8716 18593 8756 18678
rect 8715 18584 8757 18593
rect 8715 18544 8716 18584
rect 8756 18544 8757 18584
rect 8715 18535 8757 18544
rect 8620 17709 8660 17718
rect 9004 17669 9044 20224
rect 9099 20096 9141 20105
rect 9099 20056 9100 20096
rect 9140 20056 9141 20096
rect 9099 20047 9141 20056
rect 9196 20096 9236 21139
rect 9100 19962 9140 20047
rect 9196 19844 9236 20056
rect 9100 19804 9236 19844
rect 9100 19181 9140 19804
rect 9292 19601 9332 21400
rect 9388 20264 9428 20273
rect 9388 19937 9428 20224
rect 9387 19928 9429 19937
rect 9387 19888 9388 19928
rect 9428 19888 9429 19928
rect 9387 19879 9429 19888
rect 9291 19592 9333 19601
rect 9291 19552 9292 19592
rect 9332 19552 9333 19592
rect 9291 19543 9333 19552
rect 9099 19172 9141 19181
rect 9099 19132 9100 19172
rect 9140 19132 9141 19172
rect 9099 19123 9141 19132
rect 9003 17660 9045 17669
rect 9003 17620 9004 17660
rect 9044 17620 9045 17660
rect 9003 17611 9045 17620
rect 9100 17576 9140 19123
rect 9484 18929 9524 21568
rect 9676 21557 9716 21568
rect 9771 21608 9813 21617
rect 9771 21568 9772 21608
rect 9812 21568 9813 21608
rect 9771 21559 9813 21568
rect 9772 21197 9812 21559
rect 9771 21188 9813 21197
rect 9771 21148 9772 21188
rect 9812 21148 9813 21188
rect 9771 21139 9813 21148
rect 9580 20777 9620 20862
rect 9579 20768 9621 20777
rect 9579 20728 9580 20768
rect 9620 20728 9621 20768
rect 9579 20719 9621 20728
rect 9579 20600 9621 20609
rect 9579 20560 9580 20600
rect 9620 20560 9621 20600
rect 9579 20551 9621 20560
rect 9483 18920 9525 18929
rect 9483 18880 9484 18920
rect 9524 18880 9525 18920
rect 9483 18871 9525 18880
rect 9195 18164 9237 18173
rect 9195 18124 9196 18164
rect 9236 18124 9237 18164
rect 9195 18115 9237 18124
rect 9196 18005 9236 18115
rect 9195 17996 9237 18005
rect 9195 17956 9196 17996
rect 9236 17956 9237 17996
rect 9195 17947 9237 17956
rect 9196 17749 9236 17947
rect 9483 17912 9525 17921
rect 9483 17872 9484 17912
rect 9524 17872 9525 17912
rect 9483 17863 9525 17872
rect 9196 17700 9236 17709
rect 9387 17744 9429 17753
rect 9387 17704 9388 17744
rect 9428 17704 9429 17744
rect 9387 17695 9429 17704
rect 9484 17744 9524 17863
rect 9291 17660 9333 17669
rect 9291 17620 9292 17660
rect 9332 17620 9333 17660
rect 9291 17611 9333 17620
rect 8812 17534 8852 17543
rect 9100 17536 9236 17576
rect 8715 17408 8757 17417
rect 8812 17408 8852 17494
rect 8715 17368 8716 17408
rect 8756 17368 8852 17408
rect 8715 17359 8757 17368
rect 9003 17240 9045 17249
rect 9003 17200 9004 17240
rect 9044 17200 9045 17240
rect 9003 17191 9045 17200
rect 8620 17072 8660 17081
rect 8524 17032 8620 17072
rect 8620 17023 8660 17032
rect 8907 16400 8949 16409
rect 8907 16360 8908 16400
rect 8948 16360 8949 16400
rect 8907 16351 8949 16360
rect 8331 16232 8373 16241
rect 8331 16192 8332 16232
rect 8372 16192 8373 16232
rect 8331 16183 8373 16192
rect 8908 16232 8948 16351
rect 8908 16183 8948 16192
rect 8235 15812 8277 15821
rect 8235 15772 8236 15812
rect 8276 15772 8277 15812
rect 8235 15763 8277 15772
rect 8043 15140 8085 15149
rect 8043 15100 8044 15140
rect 8084 15100 8085 15140
rect 8043 15091 8085 15100
rect 7947 15056 7989 15065
rect 7947 15016 7948 15056
rect 7988 15016 7989 15056
rect 7947 15007 7989 15016
rect 7948 14729 7988 15007
rect 8139 14972 8181 14981
rect 8139 14932 8140 14972
rect 8180 14932 8181 14972
rect 8139 14923 8181 14932
rect 8140 14838 8180 14923
rect 7947 14720 7989 14729
rect 7947 14680 7948 14720
rect 7988 14680 7989 14720
rect 7947 14671 7989 14680
rect 7948 14141 7988 14671
rect 8043 14468 8085 14477
rect 8043 14428 8044 14468
rect 8084 14428 8085 14468
rect 8043 14419 8085 14428
rect 8044 14216 8084 14419
rect 8044 14167 8084 14176
rect 8235 14216 8277 14225
rect 8235 14176 8236 14216
rect 8276 14176 8277 14216
rect 8235 14167 8277 14176
rect 7947 14132 7989 14141
rect 7947 14092 7948 14132
rect 7988 14092 7989 14132
rect 7947 14083 7989 14092
rect 8236 14082 8276 14167
rect 7852 13973 7892 14008
rect 7851 13964 7893 13973
rect 7851 13924 7852 13964
rect 7892 13924 7893 13964
rect 7851 13915 7893 13924
rect 8044 13796 8084 13805
rect 7660 13672 7796 13712
rect 7659 13544 7701 13553
rect 7659 13504 7660 13544
rect 7700 13504 7701 13544
rect 7659 13495 7701 13504
rect 7467 12872 7509 12881
rect 7467 12832 7468 12872
rect 7508 12832 7509 12872
rect 7467 12823 7509 12832
rect 7084 11647 7124 11656
rect 7180 12664 7316 12704
rect 7371 12704 7413 12713
rect 7371 12664 7372 12704
rect 7412 12664 7413 12704
rect 6604 11562 6644 11647
rect 6892 11562 6932 11647
rect 6700 11528 6740 11537
rect 6603 11444 6645 11453
rect 6603 11404 6604 11444
rect 6644 11404 6645 11444
rect 6603 11395 6645 11404
rect 6604 11285 6644 11395
rect 6603 11276 6645 11285
rect 6603 11236 6604 11276
rect 6644 11236 6645 11276
rect 6603 11227 6645 11236
rect 5931 11192 5973 11201
rect 5931 11152 5932 11192
rect 5972 11152 5973 11192
rect 5931 11143 5973 11152
rect 6124 11192 6164 11201
rect 6507 11192 6549 11201
rect 6164 11152 6260 11192
rect 6124 11143 6164 11152
rect 5492 10816 5588 10856
rect 5452 10807 5492 10816
rect 5644 10772 5684 10781
rect 5548 10732 5644 10772
rect 5355 10604 5397 10613
rect 5355 10564 5356 10604
rect 5396 10564 5397 10604
rect 5355 10555 5397 10564
rect 5548 10436 5588 10732
rect 5644 10723 5684 10732
rect 5356 10396 5588 10436
rect 4780 10135 4820 10144
rect 4875 10184 4917 10193
rect 4875 10144 4876 10184
rect 4916 10144 4917 10184
rect 4875 10135 4917 10144
rect 5159 10184 5199 10193
rect 4876 10050 4916 10135
rect 5159 10025 5199 10144
rect 5259 10184 5301 10193
rect 5259 10144 5260 10184
rect 5300 10144 5301 10184
rect 5259 10135 5301 10144
rect 5356 10184 5396 10396
rect 5643 10352 5685 10361
rect 5643 10312 5644 10352
rect 5684 10312 5685 10352
rect 5643 10303 5685 10312
rect 5356 10135 5396 10144
rect 5451 10184 5493 10193
rect 5451 10144 5452 10184
rect 5492 10144 5493 10184
rect 5451 10135 5493 10144
rect 5548 10184 5588 10193
rect 5260 10050 5300 10135
rect 5158 10016 5200 10025
rect 5158 9976 5159 10016
rect 5199 9976 5200 10016
rect 5158 9967 5200 9976
rect 5356 10016 5396 10025
rect 4928 9848 5296 9857
rect 4684 9773 4724 9817
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4683 9764 4725 9773
rect 4683 9724 4684 9764
rect 4724 9724 4725 9764
rect 4683 9722 4725 9724
rect 4683 9715 4684 9722
rect 4724 9715 4725 9722
rect 4684 9673 4724 9682
rect 5356 9680 5396 9976
rect 5068 9640 5396 9680
rect 5452 9680 5492 10135
rect 5548 9848 5588 10144
rect 5644 10184 5684 10303
rect 5644 10135 5684 10144
rect 5740 9848 5780 10975
rect 5836 10949 5876 10984
rect 5932 11024 5972 11143
rect 5972 10984 6068 11024
rect 5932 10975 5972 10984
rect 5835 10940 5877 10949
rect 5835 10900 5836 10940
rect 5876 10900 5877 10940
rect 5835 10891 5877 10900
rect 5836 10889 5876 10891
rect 6028 10184 6068 10984
rect 6028 10109 6068 10144
rect 6027 10100 6069 10109
rect 6027 10060 6028 10100
rect 6068 10060 6069 10100
rect 6027 10051 6069 10060
rect 5931 10016 5973 10025
rect 6028 10020 6068 10051
rect 5931 9976 5932 10016
rect 5972 9976 5973 10016
rect 5931 9967 5973 9976
rect 6124 10016 6164 10025
rect 5548 9808 5780 9848
rect 5644 9680 5684 9689
rect 5452 9640 5644 9680
rect 4876 9512 4916 9521
rect 4876 9017 4916 9472
rect 4972 9512 5012 9521
rect 4875 9008 4917 9017
rect 4875 8968 4876 9008
rect 4916 8968 4917 9008
rect 4875 8959 4917 8968
rect 4972 8933 5012 9472
rect 5068 9512 5108 9640
rect 5644 9631 5684 9640
rect 5068 9463 5108 9472
rect 5163 9512 5205 9521
rect 5163 9472 5164 9512
rect 5204 9472 5205 9512
rect 5163 9463 5205 9472
rect 5548 9512 5588 9521
rect 5164 9378 5204 9463
rect 4971 8924 5013 8933
rect 4971 8884 4972 8924
rect 5012 8884 5013 8924
rect 4971 8875 5013 8884
rect 5548 8849 5588 9472
rect 4779 8840 4821 8849
rect 4779 8800 4780 8840
rect 4820 8800 4821 8840
rect 4779 8791 4821 8800
rect 5547 8840 5589 8849
rect 5547 8800 5548 8840
rect 5588 8800 5589 8840
rect 5547 8791 5589 8800
rect 4683 8756 4725 8765
rect 4683 8716 4684 8756
rect 4724 8716 4725 8756
rect 4683 8707 4725 8716
rect 4684 8672 4724 8707
rect 4684 8621 4724 8632
rect 4780 8597 4820 8791
rect 4875 8672 4917 8681
rect 4875 8632 4876 8672
rect 4916 8632 4917 8672
rect 4875 8623 4917 8632
rect 4779 8588 4821 8597
rect 4779 8548 4780 8588
rect 4820 8548 4821 8588
rect 4779 8539 4821 8548
rect 4683 8420 4725 8429
rect 4683 8380 4684 8420
rect 4724 8380 4725 8420
rect 4683 8371 4725 8380
rect 4684 8000 4724 8371
rect 4684 7951 4724 7960
rect 4780 8000 4820 8539
rect 4876 8538 4916 8623
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4684 7832 4724 7841
rect 4588 7792 4684 7832
rect 4684 7783 4724 7792
rect 4396 7624 4532 7664
rect 4396 7160 4436 7624
rect 4780 7589 4820 7960
rect 4971 8000 5013 8009
rect 4971 7960 4972 8000
rect 5012 7960 5013 8000
rect 4971 7951 5013 7960
rect 4972 7866 5012 7951
rect 4779 7580 4821 7589
rect 4779 7540 4780 7580
rect 4820 7540 4821 7580
rect 4779 7531 4821 7540
rect 4492 7421 4532 7506
rect 4683 7496 4725 7505
rect 4683 7456 4684 7496
rect 4724 7456 4725 7496
rect 4683 7447 4725 7456
rect 4491 7412 4533 7421
rect 4491 7372 4492 7412
rect 4532 7372 4533 7412
rect 4491 7363 4533 7372
rect 4492 7160 4532 7169
rect 4396 7120 4492 7160
rect 4492 7111 4532 7120
rect 4300 2500 4532 2540
rect 4107 1952 4149 1961
rect 4107 1912 4108 1952
rect 4148 1912 4149 1952
rect 4107 1903 4149 1912
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 3244 1156 3764 1196
rect 3531 860 3573 869
rect 3531 820 3532 860
rect 3572 820 3573 860
rect 3531 811 3573 820
rect 3339 104 3381 113
rect 3339 80 3340 104
rect 1784 0 1864 80
rect 1976 0 2056 80
rect 2168 0 2248 80
rect 2360 0 2440 80
rect 2552 0 2632 80
rect 2744 0 2824 80
rect 2936 0 3016 80
rect 3128 0 3208 80
rect 3320 64 3340 80
rect 3380 80 3381 104
rect 3532 80 3572 811
rect 3724 80 3764 1156
rect 3915 356 3957 365
rect 3915 316 3916 356
rect 3956 316 3957 356
rect 3915 307 3957 316
rect 3916 80 3956 307
rect 4108 80 4148 1903
rect 4299 524 4341 533
rect 4299 484 4300 524
rect 4340 484 4341 524
rect 4299 475 4341 484
rect 4300 80 4340 475
rect 4492 80 4532 2500
rect 4684 80 4724 7447
rect 5740 7421 5780 9808
rect 5835 9848 5877 9857
rect 5835 9808 5836 9848
rect 5876 9808 5877 9848
rect 5835 9799 5877 9808
rect 5836 9512 5876 9799
rect 5836 8429 5876 9472
rect 5932 9344 5972 9967
rect 6124 9764 6164 9976
rect 6028 9724 6164 9764
rect 6028 9512 6068 9724
rect 6220 9722 6260 11152
rect 6507 11152 6508 11192
rect 6548 11152 6549 11192
rect 6507 11143 6549 11152
rect 6315 11024 6357 11033
rect 6315 10984 6316 11024
rect 6356 10984 6357 11024
rect 6315 10975 6357 10984
rect 6412 11024 6452 11033
rect 6316 10890 6356 10975
rect 6412 10697 6452 10984
rect 6411 10688 6453 10697
rect 6411 10648 6412 10688
rect 6452 10648 6453 10688
rect 6411 10639 6453 10648
rect 6316 10184 6356 10193
rect 6508 10184 6548 11143
rect 6700 11024 6740 11488
rect 7180 11453 7220 12664
rect 7371 12655 7413 12664
rect 7276 12536 7316 12545
rect 7276 11957 7316 12496
rect 7372 12536 7412 12655
rect 7372 12487 7412 12496
rect 7467 12200 7509 12209
rect 7467 12160 7468 12200
rect 7508 12160 7509 12200
rect 7467 12151 7509 12160
rect 7275 11948 7317 11957
rect 7275 11908 7276 11948
rect 7316 11908 7317 11948
rect 7275 11899 7317 11908
rect 7179 11444 7221 11453
rect 7179 11404 7180 11444
rect 7220 11404 7221 11444
rect 7179 11395 7221 11404
rect 7083 11276 7125 11285
rect 7083 11236 7084 11276
rect 7124 11236 7125 11276
rect 7083 11227 7125 11236
rect 6603 10772 6645 10781
rect 6603 10732 6604 10772
rect 6644 10732 6645 10772
rect 6603 10723 6645 10732
rect 6604 10638 6644 10723
rect 6356 10144 6548 10184
rect 6316 10135 6356 10144
rect 6315 10016 6357 10025
rect 6315 9976 6316 10016
rect 6356 9976 6357 10016
rect 6315 9967 6357 9976
rect 6700 10016 6740 10984
rect 6892 10856 6932 10865
rect 6219 9682 6260 9722
rect 6219 9680 6259 9682
rect 6028 9463 6068 9472
rect 6124 9640 6259 9680
rect 6028 9344 6068 9353
rect 5932 9304 6028 9344
rect 6028 9295 6068 9304
rect 6124 9176 6164 9640
rect 6316 9512 6356 9967
rect 6700 9680 6740 9976
rect 6700 9631 6740 9640
rect 6796 10816 6892 10856
rect 6220 9498 6260 9507
rect 6316 9463 6356 9472
rect 6411 9512 6453 9521
rect 6411 9472 6412 9512
rect 6452 9472 6453 9512
rect 6411 9463 6453 9472
rect 6220 9353 6260 9458
rect 6219 9344 6261 9353
rect 6219 9304 6220 9344
rect 6260 9304 6261 9344
rect 6219 9295 6261 9304
rect 6028 9136 6164 9176
rect 5835 8420 5877 8429
rect 5835 8380 5836 8420
rect 5876 8380 5877 8420
rect 5835 8371 5877 8380
rect 5835 8252 5877 8261
rect 5835 8212 5836 8252
rect 5876 8212 5877 8252
rect 5835 8203 5877 8212
rect 5739 7412 5781 7421
rect 5739 7372 5740 7412
rect 5780 7372 5781 7412
rect 5739 7363 5781 7372
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 5739 2120 5781 2129
rect 5739 2080 5740 2120
rect 5780 2080 5781 2120
rect 5739 2071 5781 2080
rect 5740 1986 5780 2071
rect 5355 1028 5397 1037
rect 5355 988 5356 1028
rect 5396 988 5397 1028
rect 5355 979 5397 988
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 5356 524 5396 979
rect 5643 776 5685 785
rect 5643 736 5644 776
rect 5684 736 5685 776
rect 5643 727 5685 736
rect 5451 608 5493 617
rect 5451 568 5452 608
rect 5492 568 5493 608
rect 5451 559 5493 568
rect 5260 484 5396 524
rect 5067 272 5109 281
rect 5067 232 5068 272
rect 5108 232 5109 272
rect 5067 223 5109 232
rect 4875 188 4917 197
rect 4875 148 4876 188
rect 4916 148 4917 188
rect 4875 139 4917 148
rect 4876 80 4916 139
rect 5068 80 5108 223
rect 5260 80 5300 484
rect 5452 80 5492 559
rect 5644 80 5684 727
rect 5836 80 5876 8203
rect 6028 8177 6068 9136
rect 6316 8924 6356 8933
rect 6412 8924 6452 9463
rect 6356 8884 6452 8924
rect 6316 8875 6356 8884
rect 6123 8840 6165 8849
rect 6123 8800 6124 8840
rect 6164 8800 6165 8840
rect 6123 8791 6165 8800
rect 6124 8672 6164 8791
rect 6315 8756 6357 8765
rect 6315 8716 6316 8756
rect 6356 8716 6357 8756
rect 6315 8707 6357 8716
rect 6124 8623 6164 8632
rect 6316 8429 6356 8707
rect 6604 8504 6644 8513
rect 6796 8504 6836 10816
rect 6892 10807 6932 10816
rect 7084 10772 7124 11227
rect 7179 11024 7221 11033
rect 7179 10984 7180 11024
rect 7220 10984 7221 11024
rect 7179 10975 7221 10984
rect 7180 10890 7220 10975
rect 7084 10732 7220 10772
rect 6988 10361 7028 10446
rect 6987 10352 7029 10361
rect 6987 10312 6988 10352
rect 7028 10312 7029 10352
rect 6987 10303 7029 10312
rect 6988 10184 7028 10193
rect 6988 9773 7028 10144
rect 7084 10184 7124 10193
rect 7084 9857 7124 10144
rect 7083 9848 7125 9857
rect 7083 9808 7084 9848
rect 7124 9808 7125 9848
rect 7083 9799 7125 9808
rect 6987 9764 7029 9773
rect 6987 9724 6988 9764
rect 7028 9724 7029 9764
rect 6987 9715 7029 9724
rect 6987 9512 7029 9521
rect 6987 9472 6988 9512
rect 7028 9472 7029 9512
rect 6987 9463 7029 9472
rect 7084 9512 7124 9521
rect 6988 9378 7028 9463
rect 6891 9344 6933 9353
rect 6891 9304 6892 9344
rect 6932 9304 6933 9344
rect 6891 9295 6933 9304
rect 6892 8672 6932 9295
rect 6987 9176 7029 9185
rect 6987 9136 6988 9176
rect 7028 9136 7029 9176
rect 6987 9127 7029 9136
rect 6892 8623 6932 8632
rect 6644 8464 6836 8504
rect 6315 8420 6357 8429
rect 6315 8380 6316 8420
rect 6356 8380 6357 8420
rect 6315 8371 6357 8380
rect 6027 8168 6069 8177
rect 6027 8128 6028 8168
rect 6068 8128 6069 8168
rect 6027 8119 6069 8128
rect 6316 7832 6356 7841
rect 6316 7673 6356 7792
rect 6604 7832 6644 8464
rect 6604 7673 6644 7792
rect 6315 7664 6357 7673
rect 6315 7624 6316 7664
rect 6356 7624 6357 7664
rect 6315 7615 6357 7624
rect 6603 7664 6645 7673
rect 6603 7624 6604 7664
rect 6644 7624 6645 7664
rect 6603 7615 6645 7624
rect 6508 7160 6548 7169
rect 6604 7160 6644 7615
rect 6548 7120 6644 7160
rect 6508 7111 6548 7120
rect 6604 6656 6644 7120
rect 6604 5816 6644 6616
rect 6988 5825 7028 9127
rect 7084 8765 7124 9472
rect 7083 8756 7125 8765
rect 7083 8716 7084 8756
rect 7124 8716 7125 8756
rect 7083 8707 7125 8716
rect 7180 8345 7220 10732
rect 7275 10268 7317 10277
rect 7275 10228 7276 10268
rect 7316 10228 7317 10268
rect 7275 10219 7317 10228
rect 7276 10184 7316 10219
rect 7276 10133 7316 10144
rect 7468 9596 7508 12151
rect 7564 12125 7604 13168
rect 7660 13208 7700 13495
rect 7660 13159 7700 13168
rect 7756 12620 7796 13672
rect 8044 13553 8084 13756
rect 8236 13796 8276 13805
rect 8043 13544 8085 13553
rect 8043 13504 8044 13544
rect 8084 13504 8085 13544
rect 8043 13495 8085 13504
rect 7851 13208 7893 13217
rect 7851 13168 7852 13208
rect 7892 13168 7893 13208
rect 7851 13159 7893 13168
rect 7948 13208 7988 13217
rect 7852 13074 7892 13159
rect 7948 13049 7988 13168
rect 8140 13208 8180 13217
rect 8236 13208 8276 13756
rect 8180 13168 8276 13208
rect 8332 13208 8372 16183
rect 8620 15644 8660 15653
rect 8523 15560 8565 15569
rect 8428 15546 8468 15555
rect 8523 15520 8524 15560
rect 8564 15520 8565 15560
rect 8523 15511 8565 15520
rect 8428 14981 8468 15506
rect 8427 14972 8469 14981
rect 8427 14932 8428 14972
rect 8468 14932 8469 14972
rect 8427 14923 8469 14932
rect 8524 14720 8564 15511
rect 8524 14477 8564 14680
rect 8523 14468 8565 14477
rect 8523 14428 8524 14468
rect 8564 14428 8565 14468
rect 8523 14419 8565 14428
rect 8428 14048 8468 14057
rect 8428 13973 8468 14008
rect 8427 13964 8469 13973
rect 8427 13924 8428 13964
rect 8468 13924 8469 13964
rect 8427 13915 8469 13924
rect 8140 13159 8180 13168
rect 8332 13124 8372 13168
rect 8236 13084 8372 13124
rect 7947 13040 7989 13049
rect 7947 13000 7948 13040
rect 7988 13000 7989 13040
rect 7947 12991 7989 13000
rect 8140 13040 8180 13051
rect 8140 12965 8180 13000
rect 8139 12956 8181 12965
rect 8139 12916 8140 12956
rect 8180 12916 8181 12956
rect 8139 12907 8181 12916
rect 7851 12872 7893 12881
rect 7851 12832 7852 12872
rect 7892 12832 7893 12872
rect 7851 12823 7893 12832
rect 7660 12580 7796 12620
rect 7563 12116 7605 12125
rect 7563 12076 7564 12116
rect 7604 12076 7605 12116
rect 7563 12067 7605 12076
rect 7563 11696 7605 11705
rect 7563 11656 7564 11696
rect 7604 11656 7605 11696
rect 7563 11647 7605 11656
rect 7564 11562 7604 11647
rect 7660 11360 7700 12580
rect 7852 12536 7892 12823
rect 7852 12487 7892 12496
rect 8139 12536 8181 12545
rect 8139 12496 8140 12536
rect 8180 12496 8181 12536
rect 8139 12487 8181 12496
rect 7756 12452 7796 12461
rect 7756 11537 7796 12412
rect 7947 12116 7989 12125
rect 7947 12076 7948 12116
rect 7988 12076 7989 12116
rect 7947 12067 7989 12076
rect 7755 11528 7797 11537
rect 7755 11488 7756 11528
rect 7796 11488 7797 11528
rect 7755 11479 7797 11488
rect 7564 11320 7700 11360
rect 7564 10193 7604 11320
rect 7563 10184 7605 10193
rect 7563 10144 7564 10184
rect 7604 10144 7605 10184
rect 7563 10135 7605 10144
rect 7564 10050 7604 10135
rect 7468 9556 7604 9596
rect 7564 9512 7604 9556
rect 7468 9470 7508 9479
rect 7564 9463 7604 9472
rect 7468 9428 7508 9430
rect 7276 9388 7508 9428
rect 7276 8429 7316 9388
rect 7467 9260 7509 9269
rect 7467 9220 7468 9260
rect 7508 9220 7509 9260
rect 7467 9211 7509 9220
rect 7371 9092 7413 9101
rect 7371 9052 7372 9092
rect 7412 9052 7413 9092
rect 7371 9043 7413 9052
rect 7275 8420 7317 8429
rect 7275 8380 7276 8420
rect 7316 8380 7317 8420
rect 7275 8371 7317 8380
rect 7179 8336 7221 8345
rect 7179 8296 7180 8336
rect 7220 8296 7221 8336
rect 7179 8287 7221 8296
rect 7179 8168 7221 8177
rect 7179 8128 7180 8168
rect 7220 8128 7221 8168
rect 7179 8119 7221 8128
rect 7180 8000 7220 8119
rect 7180 7951 7220 7960
rect 6604 5144 6644 5776
rect 6987 5816 7029 5825
rect 6987 5776 6988 5816
rect 7028 5776 7029 5816
rect 6987 5767 7029 5776
rect 6604 4304 6644 5104
rect 6411 3800 6453 3809
rect 6411 3760 6412 3800
rect 6452 3760 6453 3800
rect 6411 3751 6453 3760
rect 6123 2204 6165 2213
rect 6123 2164 6124 2204
rect 6164 2164 6165 2204
rect 6123 2155 6165 2164
rect 6124 2120 6164 2155
rect 6124 2069 6164 2080
rect 5932 1868 5972 1877
rect 5932 1541 5972 1828
rect 6316 1868 6356 1877
rect 5931 1532 5973 1541
rect 5931 1492 5932 1532
rect 5972 1492 5973 1532
rect 5931 1483 5973 1492
rect 6316 1457 6356 1828
rect 6315 1448 6357 1457
rect 6315 1408 6316 1448
rect 6356 1408 6357 1448
rect 6315 1399 6357 1408
rect 6027 1280 6069 1289
rect 6027 1240 6028 1280
rect 6068 1240 6069 1280
rect 6027 1231 6069 1240
rect 6028 80 6068 1231
rect 6412 953 6452 3751
rect 6604 3632 6644 4264
rect 6604 3583 6644 3592
rect 6891 2876 6933 2885
rect 6891 2836 6892 2876
rect 6932 2836 6933 2876
rect 6891 2827 6933 2836
rect 6892 2742 6932 2827
rect 7084 2708 7124 2717
rect 6507 2120 6549 2129
rect 6507 2080 6508 2120
rect 6548 2080 6549 2120
rect 6507 2071 6549 2080
rect 6891 2120 6933 2129
rect 6891 2080 6892 2120
rect 6932 2080 6933 2120
rect 6891 2071 6933 2080
rect 6508 1986 6548 2071
rect 6892 1986 6932 2071
rect 7084 2045 7124 2668
rect 7372 2540 7412 9043
rect 7468 7589 7508 9211
rect 7756 7757 7796 11479
rect 7851 11444 7893 11453
rect 7851 11404 7852 11444
rect 7892 11404 7893 11444
rect 7851 11395 7893 11404
rect 7755 7748 7797 7757
rect 7755 7708 7756 7748
rect 7796 7708 7797 7748
rect 7755 7699 7797 7708
rect 7467 7580 7509 7589
rect 7467 7540 7468 7580
rect 7508 7540 7509 7580
rect 7467 7531 7509 7540
rect 7755 7496 7797 7505
rect 7755 7456 7756 7496
rect 7796 7456 7797 7496
rect 7755 7447 7797 7456
rect 7756 7160 7796 7447
rect 7756 7111 7796 7120
rect 7852 3809 7892 11395
rect 7948 11360 7988 12067
rect 8140 11360 8180 12487
rect 8236 11873 8276 13084
rect 8332 12629 8372 12660
rect 8331 12620 8373 12629
rect 8331 12580 8332 12620
rect 8372 12580 8373 12620
rect 8331 12571 8373 12580
rect 8332 12536 8372 12571
rect 8235 11864 8277 11873
rect 8235 11824 8236 11864
rect 8276 11824 8277 11864
rect 8235 11815 8277 11824
rect 8332 11789 8372 12496
rect 8331 11780 8373 11789
rect 8331 11740 8332 11780
rect 8372 11740 8373 11780
rect 8331 11731 8373 11740
rect 7948 11320 8084 11360
rect 8140 11320 8276 11360
rect 8044 11276 8084 11320
rect 8044 11236 8180 11276
rect 8140 10697 8180 11236
rect 8139 10688 8181 10697
rect 8139 10648 8140 10688
rect 8180 10648 8181 10688
rect 8139 10639 8181 10648
rect 8043 9512 8085 9521
rect 8043 9472 8044 9512
rect 8084 9472 8085 9512
rect 8043 9463 8085 9472
rect 8044 9378 8084 9463
rect 8140 9260 8180 10639
rect 8044 9220 8180 9260
rect 8044 7925 8084 9220
rect 8139 8840 8181 8849
rect 8139 8800 8140 8840
rect 8180 8800 8181 8840
rect 8139 8791 8181 8800
rect 8140 8672 8180 8791
rect 8236 8756 8276 11320
rect 8428 11024 8468 13915
rect 8620 11360 8660 15604
rect 8907 15644 8949 15653
rect 8907 15604 8908 15644
rect 8948 15604 8949 15644
rect 8907 15595 8949 15604
rect 8908 15560 8948 15595
rect 8908 15317 8948 15520
rect 8907 15308 8949 15317
rect 8907 15268 8908 15308
rect 8948 15268 8949 15308
rect 8907 15259 8949 15268
rect 8715 15140 8757 15149
rect 8715 15100 8716 15140
rect 8756 15100 8757 15140
rect 8715 15091 8757 15100
rect 8716 14477 8756 15091
rect 8811 14888 8853 14897
rect 8811 14848 8812 14888
rect 8852 14848 8857 14888
rect 8811 14839 8857 14848
rect 8817 14729 8857 14839
rect 8812 14720 8857 14729
rect 8852 14689 8857 14720
rect 8812 14671 8852 14680
rect 8908 14636 8948 14645
rect 8715 14468 8757 14477
rect 8715 14428 8716 14468
rect 8756 14428 8757 14468
rect 8715 14419 8757 14428
rect 8908 13553 8948 14596
rect 8907 13544 8949 13553
rect 8907 13504 8908 13544
rect 8948 13504 8949 13544
rect 8907 13495 8949 13504
rect 8716 13301 8756 13320
rect 8715 13292 8757 13301
rect 9004 13292 9044 17191
rect 9100 17058 9140 17067
rect 9100 16484 9140 17018
rect 9100 16435 9140 16444
rect 9196 16316 9236 17536
rect 9292 17526 9332 17611
rect 9100 16276 9236 16316
rect 9292 17156 9332 17165
rect 9100 16157 9140 16276
rect 9099 16148 9141 16157
rect 9099 16108 9100 16148
rect 9140 16108 9141 16148
rect 9099 16099 9141 16108
rect 8715 13252 8716 13292
rect 8756 13252 9044 13292
rect 8715 13243 8757 13252
rect 9100 12713 9140 16099
rect 9196 14888 9236 14897
rect 9196 14729 9236 14848
rect 9195 14720 9237 14729
rect 9195 14680 9196 14720
rect 9236 14680 9237 14720
rect 9195 14671 9237 14680
rect 9099 12704 9141 12713
rect 9099 12664 9100 12704
rect 9140 12664 9141 12704
rect 9099 12655 9141 12664
rect 9003 12620 9045 12629
rect 9003 12580 9004 12620
rect 9044 12580 9045 12620
rect 9003 12571 9045 12580
rect 8812 12522 8852 12531
rect 9004 12486 9044 12571
rect 8812 12032 8852 12482
rect 9196 12368 9236 12377
rect 8812 11992 9044 12032
rect 9004 11948 9044 11992
rect 9004 11899 9044 11908
rect 8811 11864 8853 11873
rect 8811 11824 8812 11864
rect 8852 11824 8853 11864
rect 8811 11815 8853 11824
rect 8812 11696 8852 11815
rect 8907 11780 8949 11789
rect 8907 11740 8908 11780
rect 8948 11740 8949 11780
rect 8907 11731 8949 11740
rect 8812 11647 8852 11656
rect 8428 10949 8468 10984
rect 8524 11320 8660 11360
rect 8427 10940 8469 10949
rect 8427 10900 8428 10940
rect 8468 10900 8469 10940
rect 8427 10891 8469 10900
rect 8428 10889 8468 10891
rect 8524 9596 8564 11320
rect 8619 11108 8661 11117
rect 8619 11068 8620 11108
rect 8660 11068 8661 11108
rect 8619 11059 8661 11068
rect 8620 10974 8660 11059
rect 8811 10940 8853 10949
rect 8811 10900 8812 10940
rect 8852 10900 8853 10940
rect 8811 10891 8853 10900
rect 8812 10184 8852 10891
rect 8812 10135 8852 10144
rect 8715 9764 8757 9773
rect 8715 9724 8716 9764
rect 8756 9724 8757 9764
rect 8715 9715 8757 9724
rect 8716 9680 8756 9715
rect 8716 9629 8756 9640
rect 8524 9556 8660 9596
rect 8524 9498 8564 9507
rect 8332 8924 8372 8933
rect 8524 8924 8564 9458
rect 8372 8884 8564 8924
rect 8332 8875 8372 8884
rect 8236 8716 8372 8756
rect 8140 8623 8180 8632
rect 8043 7916 8085 7925
rect 8043 7876 8044 7916
rect 8084 7876 8085 7916
rect 8043 7867 8085 7876
rect 8236 7160 8276 7169
rect 7948 7076 7988 7085
rect 8236 7076 8276 7120
rect 7988 7036 8276 7076
rect 8332 7160 8372 8716
rect 8620 8336 8660 9556
rect 8524 8296 8660 8336
rect 8716 8672 8756 8681
rect 8428 8000 8468 8009
rect 8428 7505 8468 7960
rect 8427 7496 8469 7505
rect 8427 7456 8428 7496
rect 8468 7456 8469 7496
rect 8427 7447 8469 7456
rect 7948 7027 7988 7036
rect 7851 3800 7893 3809
rect 7851 3760 7852 3800
rect 7892 3760 7893 3800
rect 7851 3751 7893 3760
rect 7180 2500 7412 2540
rect 8332 2540 8372 7120
rect 8427 6488 8469 6497
rect 8427 6448 8428 6488
rect 8468 6448 8469 6488
rect 8427 6439 8469 6448
rect 8428 6354 8468 6439
rect 8524 2540 8564 8296
rect 8620 8168 8660 8177
rect 8716 8168 8756 8632
rect 8812 8672 8852 8681
rect 8812 8345 8852 8632
rect 8908 8513 8948 11731
rect 9196 11621 9236 12328
rect 9003 11612 9045 11621
rect 9003 11572 9004 11612
rect 9044 11572 9045 11612
rect 9003 11563 9045 11572
rect 9195 11612 9237 11621
rect 9195 11572 9196 11612
rect 9236 11572 9237 11612
rect 9195 11563 9237 11572
rect 9004 10520 9044 11563
rect 9196 11024 9236 11563
rect 9292 11285 9332 17116
rect 9388 16484 9428 17695
rect 9484 17240 9524 17704
rect 9484 17191 9524 17200
rect 9483 17072 9525 17081
rect 9483 17032 9484 17072
rect 9524 17032 9525 17072
rect 9483 17023 9525 17032
rect 9484 16577 9524 17023
rect 9483 16568 9525 16577
rect 9483 16528 9484 16568
rect 9524 16528 9525 16568
rect 9483 16519 9525 16528
rect 9388 16435 9428 16444
rect 9388 14720 9428 14729
rect 9388 14225 9428 14680
rect 9484 14468 9524 16519
rect 9580 16493 9620 20551
rect 9675 20096 9717 20105
rect 9675 20056 9676 20096
rect 9716 20056 9717 20096
rect 9675 20047 9717 20056
rect 9676 19962 9716 20047
rect 9675 19676 9717 19685
rect 9675 19636 9676 19676
rect 9716 19636 9717 19676
rect 9675 19627 9717 19636
rect 9676 19013 9716 19627
rect 9675 19004 9717 19013
rect 9675 18964 9676 19004
rect 9716 18964 9717 19004
rect 9675 18955 9717 18964
rect 9868 18509 9908 22072
rect 9964 21776 10004 21785
rect 10060 21776 10100 22240
rect 10156 22280 10196 22567
rect 10252 22541 10292 27616
rect 10347 27488 10389 27497
rect 10347 27448 10348 27488
rect 10388 27448 10389 27488
rect 10347 27439 10389 27448
rect 10348 24053 10388 27439
rect 10347 24044 10389 24053
rect 10347 24004 10348 24044
rect 10388 24004 10389 24044
rect 10347 23995 10389 24004
rect 10347 23204 10389 23213
rect 10347 23164 10348 23204
rect 10388 23164 10389 23204
rect 10347 23155 10389 23164
rect 10251 22532 10293 22541
rect 10251 22492 10252 22532
rect 10292 22492 10293 22532
rect 10251 22483 10293 22492
rect 10257 22280 10297 22289
rect 10156 22231 10196 22240
rect 10252 22240 10257 22280
rect 10252 22231 10297 22240
rect 10004 21736 10100 21776
rect 10156 22112 10196 22121
rect 9964 21727 10004 21736
rect 10156 20180 10196 22072
rect 10060 20140 10196 20180
rect 10060 19508 10100 20140
rect 10252 19769 10292 22231
rect 10348 21533 10388 23155
rect 10347 21524 10389 21533
rect 10347 21484 10348 21524
rect 10388 21484 10389 21524
rect 10347 21475 10389 21484
rect 10347 21104 10389 21113
rect 10347 21064 10348 21104
rect 10388 21064 10389 21104
rect 10347 21055 10389 21064
rect 10251 19760 10293 19769
rect 10251 19720 10252 19760
rect 10292 19720 10293 19760
rect 10251 19711 10293 19720
rect 10348 19685 10388 21055
rect 10347 19676 10389 19685
rect 10347 19636 10348 19676
rect 10388 19636 10389 19676
rect 10347 19627 10389 19636
rect 10444 19601 10484 28279
rect 10540 20105 10580 29875
rect 10828 29336 10868 30631
rect 10924 29672 10964 32656
rect 11116 31529 11156 32824
rect 11115 31520 11157 31529
rect 11115 31480 11116 31520
rect 11156 31480 11157 31520
rect 11115 31471 11157 31480
rect 11212 31436 11252 32899
rect 11307 32780 11349 32789
rect 11307 32740 11308 32780
rect 11348 32740 11349 32780
rect 11307 32731 11349 32740
rect 11212 31387 11252 31396
rect 11116 31352 11156 31361
rect 11116 30689 11156 31312
rect 11211 31016 11253 31025
rect 11211 30976 11212 31016
rect 11252 30976 11253 31016
rect 11211 30967 11253 30976
rect 11115 30680 11157 30689
rect 11115 30640 11116 30680
rect 11156 30640 11157 30680
rect 11115 30631 11157 30640
rect 11212 30680 11252 30967
rect 11212 30631 11252 30640
rect 11116 30546 11156 30631
rect 11019 29924 11061 29933
rect 11019 29884 11020 29924
rect 11060 29884 11061 29924
rect 11019 29875 11061 29884
rect 11020 29840 11060 29875
rect 11020 29789 11060 29800
rect 10924 29632 11060 29672
rect 10923 29504 10965 29513
rect 10923 29464 10924 29504
rect 10964 29464 10965 29504
rect 10923 29455 10965 29464
rect 10732 29296 10868 29336
rect 10732 29168 10772 29296
rect 10636 29128 10732 29168
rect 10636 27572 10676 29128
rect 10732 29119 10772 29128
rect 10828 29168 10868 29177
rect 10924 29168 10964 29455
rect 10868 29128 10964 29168
rect 10828 29119 10868 29128
rect 11020 29000 11060 29632
rect 11308 29168 11348 32731
rect 11404 32201 11444 33823
rect 11596 33368 11636 41299
rect 11691 38744 11733 38753
rect 11691 38704 11692 38744
rect 11732 38704 11733 38744
rect 11691 38695 11733 38704
rect 11692 38235 11732 38695
rect 11692 38186 11732 38195
rect 11788 37820 11828 41392
rect 11884 40349 11924 46264
rect 11980 44288 12020 46432
rect 12075 46432 12076 46472
rect 12116 46432 12117 46472
rect 12075 46423 12117 46432
rect 11980 44239 12020 44248
rect 11980 42776 12020 42787
rect 11980 42701 12020 42736
rect 11979 42692 12021 42701
rect 12172 42692 12212 46600
rect 12652 46397 12692 47944
rect 12651 46388 12693 46397
rect 12651 46348 12652 46388
rect 12692 46348 12693 46388
rect 12651 46339 12693 46348
rect 12651 45968 12693 45977
rect 12651 45928 12652 45968
rect 12692 45928 12693 45968
rect 12651 45919 12693 45928
rect 12652 45834 12692 45919
rect 12459 45800 12501 45809
rect 12459 45760 12460 45800
rect 12500 45760 12501 45800
rect 12459 45751 12501 45760
rect 11979 42652 11980 42692
rect 12020 42652 12021 42692
rect 11979 42643 12021 42652
rect 12076 42652 12212 42692
rect 11980 42449 12020 42643
rect 11979 42440 12021 42449
rect 11979 42400 11980 42440
rect 12020 42400 12021 42440
rect 11979 42391 12021 42400
rect 11979 41600 12021 41609
rect 11979 41560 11980 41600
rect 12020 41560 12021 41600
rect 11979 41551 12021 41560
rect 11980 41264 12020 41551
rect 12076 41357 12116 42652
rect 12172 42524 12212 42533
rect 12172 41936 12212 42484
rect 12268 41936 12308 41945
rect 12172 41896 12268 41936
rect 12268 41887 12308 41896
rect 12364 41936 12404 41945
rect 12364 41777 12404 41896
rect 12363 41768 12405 41777
rect 12363 41728 12364 41768
rect 12404 41728 12405 41768
rect 12363 41719 12405 41728
rect 12460 41432 12500 45751
rect 12652 44960 12692 44969
rect 12555 44036 12597 44045
rect 12652 44036 12692 44920
rect 12555 43996 12556 44036
rect 12596 43996 12692 44036
rect 12555 43987 12597 43996
rect 12556 43541 12596 43987
rect 12555 43532 12597 43541
rect 12555 43492 12556 43532
rect 12596 43492 12597 43532
rect 12555 43483 12597 43492
rect 12556 43448 12596 43483
rect 12748 43448 12788 49120
rect 12844 47816 12884 49288
rect 13036 48992 13076 50203
rect 13131 49496 13173 49505
rect 13131 49456 13132 49496
rect 13172 49456 13173 49496
rect 13131 49447 13173 49456
rect 13029 48952 13076 48992
rect 13132 48992 13172 49447
rect 13029 48908 13069 48952
rect 13132 48943 13172 48952
rect 12947 48868 13069 48908
rect 12947 48833 12987 48868
rect 12940 48824 12987 48833
rect 12980 48784 12987 48824
rect 12940 48665 12980 48784
rect 12939 48656 12981 48665
rect 12939 48616 12940 48656
rect 12980 48616 12981 48656
rect 12939 48607 12981 48616
rect 13035 48152 13077 48161
rect 13035 48112 13036 48152
rect 13076 48112 13077 48152
rect 13035 48103 13077 48112
rect 13036 48068 13076 48103
rect 13036 48017 13076 48028
rect 13132 48068 13172 48077
rect 13228 48068 13268 50539
rect 13419 49916 13461 49925
rect 13419 49876 13420 49916
rect 13460 49876 13461 49916
rect 13419 49867 13461 49876
rect 13420 49496 13460 49867
rect 13420 49447 13460 49456
rect 13419 48740 13461 48749
rect 13419 48700 13420 48740
rect 13460 48700 13461 48740
rect 13419 48691 13461 48700
rect 13323 48152 13365 48161
rect 13323 48112 13324 48152
rect 13364 48112 13365 48152
rect 13323 48103 13365 48112
rect 13172 48028 13268 48068
rect 13132 48019 13172 48028
rect 12844 47776 13172 47816
rect 12844 46472 12884 46481
rect 12844 46061 12884 46432
rect 12940 46472 12980 46483
rect 12940 46397 12980 46432
rect 12939 46388 12981 46397
rect 12939 46348 12940 46388
rect 12980 46348 12981 46388
rect 12939 46339 12981 46348
rect 12843 46052 12885 46061
rect 12843 46012 12844 46052
rect 12884 46012 12885 46052
rect 12843 46003 12885 46012
rect 12844 45800 12884 45809
rect 12884 45760 12980 45800
rect 12844 45751 12884 45760
rect 12844 44792 12884 44801
rect 12844 43961 12884 44752
rect 12940 44633 12980 45760
rect 12939 44624 12981 44633
rect 12939 44584 12940 44624
rect 12980 44584 12981 44624
rect 12939 44575 12981 44584
rect 12843 43952 12885 43961
rect 12843 43912 12844 43952
rect 12884 43912 12885 43952
rect 12843 43903 12885 43912
rect 12556 43397 12596 43408
rect 12652 43408 12788 43448
rect 12364 41392 12500 41432
rect 12075 41348 12117 41357
rect 12075 41308 12076 41348
rect 12116 41308 12117 41348
rect 12075 41299 12117 41308
rect 11980 41215 12020 41224
rect 11980 40424 12020 40433
rect 12020 40384 12116 40424
rect 11980 40375 12020 40384
rect 11883 40340 11925 40349
rect 11883 40300 11884 40340
rect 11924 40300 11925 40340
rect 11883 40291 11925 40300
rect 12076 38912 12116 40384
rect 12172 40256 12212 40265
rect 12172 39761 12212 40216
rect 12171 39752 12213 39761
rect 12171 39712 12172 39752
rect 12212 39712 12213 39752
rect 12171 39703 12213 39712
rect 12268 38912 12308 38921
rect 12076 38872 12268 38912
rect 12076 38417 12116 38872
rect 12268 38863 12308 38872
rect 12364 38744 12404 41392
rect 12652 40592 12692 43408
rect 12844 43373 12884 43903
rect 13132 43700 13172 47776
rect 13228 46145 13268 48028
rect 13324 46472 13364 48103
rect 13420 46556 13460 48691
rect 13420 46507 13460 46516
rect 13227 46136 13269 46145
rect 13227 46096 13228 46136
rect 13268 46096 13269 46136
rect 13227 46087 13269 46096
rect 13228 44456 13268 46087
rect 13324 46061 13364 46432
rect 13419 46388 13461 46397
rect 13419 46348 13420 46388
rect 13460 46348 13461 46388
rect 13419 46339 13461 46348
rect 13323 46052 13365 46061
rect 13323 46012 13324 46052
rect 13364 46012 13365 46052
rect 13323 46003 13365 46012
rect 13420 45473 13460 46339
rect 13419 45464 13461 45473
rect 13419 45424 13420 45464
rect 13460 45424 13461 45464
rect 13419 45415 13461 45424
rect 13324 44960 13364 44969
rect 13324 44633 13364 44920
rect 13420 44960 13460 45415
rect 13420 44911 13460 44920
rect 13323 44624 13365 44633
rect 13323 44584 13324 44624
rect 13364 44584 13365 44624
rect 13323 44575 13365 44584
rect 13516 44540 13556 50884
rect 13612 47993 13652 51220
rect 13708 51017 13748 51102
rect 13707 51008 13749 51017
rect 13707 50968 13708 51008
rect 13748 50968 13749 51008
rect 13707 50959 13749 50968
rect 13900 50849 13940 56176
rect 13995 56048 14037 56057
rect 13995 56008 13996 56048
rect 14036 56008 14037 56048
rect 13995 55999 14037 56008
rect 13996 54041 14036 55999
rect 13995 54032 14037 54041
rect 13995 53992 13996 54032
rect 14036 53992 14037 54032
rect 13995 53983 14037 53992
rect 13996 53898 14036 53983
rect 14092 52772 14132 57268
rect 14187 57056 14229 57065
rect 14187 57016 14188 57056
rect 14228 57016 14229 57056
rect 14187 57007 14229 57016
rect 14284 57056 14324 57065
rect 14324 57016 14420 57056
rect 14284 57007 14324 57016
rect 14188 56922 14228 57007
rect 14380 56813 14420 57016
rect 14379 56804 14421 56813
rect 14379 56764 14380 56804
rect 14420 56764 14421 56804
rect 14379 56755 14421 56764
rect 14283 56384 14325 56393
rect 14283 56344 14284 56384
rect 14324 56344 14325 56384
rect 14283 56335 14325 56344
rect 14380 56384 14420 56755
rect 14380 56335 14420 56344
rect 14284 56250 14324 56335
rect 14476 56132 14516 60628
rect 14284 56092 14516 56132
rect 14187 54956 14229 54965
rect 14187 54916 14188 54956
rect 14228 54916 14229 54956
rect 14187 54907 14229 54916
rect 14188 54872 14228 54907
rect 14188 54821 14228 54832
rect 14187 54032 14229 54041
rect 14187 53992 14188 54032
rect 14228 53992 14229 54032
rect 14187 53983 14229 53992
rect 14188 53360 14228 53983
rect 14188 53311 14228 53320
rect 13996 52732 14132 52772
rect 13707 50840 13749 50849
rect 13707 50800 13708 50840
rect 13748 50800 13749 50840
rect 13707 50791 13749 50800
rect 13899 50840 13941 50849
rect 13899 50800 13900 50840
rect 13940 50800 13941 50840
rect 13899 50791 13941 50800
rect 13708 48824 13748 50791
rect 13899 49664 13941 49673
rect 13899 49624 13900 49664
rect 13940 49624 13941 49664
rect 13996 49664 14036 52732
rect 14284 52688 14324 56092
rect 14476 55544 14516 55553
rect 14476 55385 14516 55504
rect 14475 55376 14517 55385
rect 14475 55336 14476 55376
rect 14516 55336 14517 55376
rect 14475 55327 14517 55336
rect 14380 54620 14420 54629
rect 14420 54580 14516 54620
rect 14380 54571 14420 54580
rect 14379 54452 14421 54461
rect 14379 54412 14380 54452
rect 14420 54412 14421 54452
rect 14379 54403 14421 54412
rect 14092 52648 14324 52688
rect 14092 51185 14132 52648
rect 14187 52520 14229 52529
rect 14187 52480 14188 52520
rect 14228 52480 14229 52520
rect 14187 52471 14229 52480
rect 14284 52520 14324 52529
rect 14188 52386 14228 52471
rect 14284 52193 14324 52480
rect 14283 52184 14325 52193
rect 14283 52144 14284 52184
rect 14324 52144 14325 52184
rect 14283 52135 14325 52144
rect 14187 51680 14229 51689
rect 14187 51640 14188 51680
rect 14228 51640 14229 51680
rect 14187 51631 14229 51640
rect 14091 51176 14133 51185
rect 14091 51136 14092 51176
rect 14132 51136 14133 51176
rect 14091 51127 14133 51136
rect 14188 51092 14228 51631
rect 14188 51043 14228 51052
rect 14091 51008 14133 51017
rect 14091 50968 14092 51008
rect 14132 50968 14133 51008
rect 14091 50959 14133 50968
rect 14284 51008 14324 51017
rect 14092 49925 14132 50959
rect 14284 50756 14324 50968
rect 14188 50716 14324 50756
rect 14091 49916 14133 49925
rect 14091 49876 14092 49916
rect 14132 49876 14133 49916
rect 14091 49867 14133 49876
rect 13996 49624 14132 49664
rect 13899 49615 13941 49624
rect 13611 47984 13653 47993
rect 13611 47944 13612 47984
rect 13652 47944 13653 47984
rect 13611 47935 13653 47944
rect 13612 47850 13652 47935
rect 13708 44885 13748 48784
rect 13900 49580 13940 49615
rect 13900 48749 13940 49540
rect 13996 49496 14036 49507
rect 13996 49421 14036 49456
rect 13995 49412 14037 49421
rect 13995 49372 13996 49412
rect 14036 49372 14037 49412
rect 13995 49363 14037 49372
rect 13899 48740 13941 48749
rect 13899 48700 13900 48740
rect 13940 48700 13941 48740
rect 13899 48691 13941 48700
rect 14092 48161 14132 49624
rect 14188 49421 14228 50716
rect 14284 50336 14324 50345
rect 14187 49412 14229 49421
rect 14187 49372 14188 49412
rect 14228 49372 14229 49412
rect 14187 49363 14229 49372
rect 14187 48656 14229 48665
rect 14187 48616 14188 48656
rect 14228 48616 14229 48656
rect 14187 48607 14229 48616
rect 14091 48152 14133 48161
rect 14091 48112 14092 48152
rect 14132 48112 14133 48152
rect 14091 48103 14133 48112
rect 13899 47984 13941 47993
rect 13899 47944 13900 47984
rect 13940 47944 13941 47984
rect 13899 47935 13941 47944
rect 14092 47989 14132 47998
rect 13803 47312 13845 47321
rect 13803 47272 13804 47312
rect 13844 47272 13845 47312
rect 13803 47263 13845 47272
rect 13804 47178 13844 47263
rect 13900 46472 13940 47935
rect 13996 47480 14036 47489
rect 14092 47480 14132 47949
rect 14036 47440 14132 47480
rect 13996 47431 14036 47440
rect 14091 46892 14133 46901
rect 14091 46852 14092 46892
rect 14132 46852 14133 46892
rect 14091 46843 14133 46852
rect 13900 46423 13940 46432
rect 13899 45968 13941 45977
rect 13899 45928 13900 45968
rect 13940 45928 13941 45968
rect 13899 45919 13941 45928
rect 13803 45044 13845 45053
rect 13803 45004 13804 45044
rect 13844 45004 13845 45044
rect 13803 44995 13845 45004
rect 13900 45044 13940 45919
rect 14092 45809 14132 46843
rect 14091 45800 14133 45809
rect 14091 45760 14092 45800
rect 14132 45760 14133 45800
rect 14091 45751 14133 45760
rect 14092 45666 14132 45751
rect 13900 44995 13940 45004
rect 13804 44910 13844 44995
rect 14188 44960 14228 48607
rect 14284 48245 14324 50296
rect 14380 49757 14420 54403
rect 14476 54046 14516 54580
rect 14476 53997 14516 54006
rect 14475 53360 14517 53369
rect 14475 53320 14476 53360
rect 14516 53320 14517 53360
rect 14475 53311 14517 53320
rect 14476 50597 14516 53311
rect 14572 51017 14612 60712
rect 14668 60593 14708 63895
rect 14764 62273 14804 64240
rect 14956 64028 14996 66835
rect 15244 66128 15284 66137
rect 15148 66088 15244 66128
rect 15148 64616 15188 66088
rect 15244 66079 15284 66088
rect 15436 65960 15476 65969
rect 15340 65920 15436 65960
rect 15340 65456 15380 65920
rect 15436 65911 15476 65920
rect 15292 65446 15380 65456
rect 15332 65416 15380 65446
rect 15436 65540 15476 65549
rect 15292 65397 15332 65406
rect 15436 65381 15476 65500
rect 15532 65465 15572 68020
rect 15628 67052 15668 68692
rect 15724 68480 15764 68692
rect 15724 68431 15764 68440
rect 15724 67724 15764 67733
rect 15724 67649 15764 67684
rect 15723 67640 15765 67649
rect 15723 67600 15724 67640
rect 15764 67600 15765 67640
rect 15723 67591 15765 67600
rect 15724 67229 15764 67591
rect 15723 67220 15765 67229
rect 15723 67180 15724 67220
rect 15764 67180 15765 67220
rect 15723 67171 15765 67180
rect 15628 67012 15764 67052
rect 15628 66926 15668 66935
rect 15627 66886 15628 66893
rect 15668 66886 15669 66893
rect 15627 66884 15669 66886
rect 15627 66844 15628 66884
rect 15668 66844 15669 66884
rect 15627 66835 15669 66844
rect 15531 65456 15573 65465
rect 15531 65416 15532 65456
rect 15572 65416 15573 65456
rect 15531 65407 15573 65416
rect 15435 65372 15477 65381
rect 15435 65332 15436 65372
rect 15476 65332 15477 65372
rect 15435 65323 15477 65332
rect 15244 64616 15284 64625
rect 15148 64576 15244 64616
rect 15148 64289 15188 64576
rect 15244 64567 15284 64576
rect 15436 64448 15476 64457
rect 15147 64280 15189 64289
rect 15147 64240 15148 64280
rect 15188 64240 15189 64280
rect 15147 64231 15189 64240
rect 14956 63953 14999 64028
rect 14955 63944 14999 63953
rect 14955 63904 14956 63944
rect 14996 63904 14999 63944
rect 15436 63939 15476 64408
rect 15628 64280 15668 66835
rect 15724 64625 15764 67012
rect 15820 66893 15860 74143
rect 15916 73025 15956 79771
rect 16108 79409 16148 79780
rect 16107 79400 16149 79409
rect 16107 79360 16108 79400
rect 16148 79360 16149 79400
rect 16107 79351 16149 79360
rect 16108 79073 16148 79351
rect 16107 79064 16149 79073
rect 16107 79024 16108 79064
rect 16148 79024 16149 79064
rect 16107 79015 16149 79024
rect 16011 78224 16053 78233
rect 16011 78184 16012 78224
rect 16052 78184 16053 78224
rect 16011 78175 16053 78184
rect 16012 78090 16052 78175
rect 16011 77804 16053 77813
rect 16011 77764 16012 77804
rect 16052 77764 16053 77804
rect 16011 77755 16053 77764
rect 16012 75704 16052 77755
rect 16108 77552 16148 79015
rect 16204 77729 16244 85936
rect 16299 80324 16341 80333
rect 16299 80284 16300 80324
rect 16340 80284 16341 80324
rect 16299 80275 16341 80284
rect 16300 77813 16340 80275
rect 16396 79409 16436 85936
rect 16492 79820 16532 79829
rect 16492 79493 16532 79780
rect 16491 79484 16533 79493
rect 16491 79444 16492 79484
rect 16532 79444 16533 79484
rect 16491 79435 16533 79444
rect 16395 79400 16437 79409
rect 16395 79360 16396 79400
rect 16436 79360 16437 79400
rect 16395 79351 16437 79360
rect 16588 79232 16628 85936
rect 16780 81920 16820 85936
rect 16972 85625 17012 85936
rect 16971 85616 17013 85625
rect 16971 85576 16972 85616
rect 17012 85576 17013 85616
rect 16971 85567 17013 85576
rect 17164 84449 17204 85936
rect 17356 84533 17396 85936
rect 17355 84524 17397 84533
rect 17355 84484 17356 84524
rect 17396 84484 17397 84524
rect 17355 84475 17397 84484
rect 17548 84449 17588 85936
rect 17740 84617 17780 85936
rect 17932 85121 17972 85936
rect 18027 85448 18069 85457
rect 18027 85408 18028 85448
rect 18068 85408 18069 85448
rect 18027 85399 18069 85408
rect 17931 85112 17973 85121
rect 17931 85072 17932 85112
rect 17972 85072 17973 85112
rect 17931 85063 17973 85072
rect 17739 84608 17781 84617
rect 17739 84568 17740 84608
rect 17780 84568 17781 84608
rect 17739 84559 17781 84568
rect 17163 84440 17205 84449
rect 17163 84400 17164 84440
rect 17204 84400 17205 84440
rect 17163 84391 17205 84400
rect 17547 84440 17589 84449
rect 17547 84400 17548 84440
rect 17588 84400 17589 84440
rect 17547 84391 17589 84400
rect 18028 83768 18068 85399
rect 18124 84449 18164 85936
rect 18316 84533 18356 85936
rect 18315 84524 18357 84533
rect 18315 84484 18316 84524
rect 18356 84484 18357 84524
rect 18315 84475 18357 84484
rect 18508 84449 18548 85936
rect 18700 84533 18740 85936
rect 18892 84953 18932 85936
rect 19083 85912 19084 85936
rect 19124 85936 19144 85952
rect 19256 85952 19336 86016
rect 19256 85936 19276 85952
rect 19124 85912 19125 85936
rect 19083 85903 19125 85912
rect 19275 85912 19276 85936
rect 19316 85936 19336 85952
rect 19448 85936 19528 86016
rect 19316 85912 19317 85936
rect 19275 85903 19317 85912
rect 19275 85784 19317 85793
rect 19275 85744 19276 85784
rect 19316 85744 19317 85784
rect 19275 85735 19317 85744
rect 18891 84944 18933 84953
rect 18891 84904 18892 84944
rect 18932 84904 18933 84944
rect 18891 84895 18933 84904
rect 18808 84692 19176 84701
rect 18848 84652 18890 84692
rect 18930 84652 18972 84692
rect 19012 84652 19054 84692
rect 19094 84652 19136 84692
rect 18808 84643 19176 84652
rect 18699 84524 18741 84533
rect 19276 84524 19316 85735
rect 18699 84484 18700 84524
rect 18740 84484 18741 84524
rect 18699 84475 18741 84484
rect 19180 84484 19316 84524
rect 18123 84440 18165 84449
rect 18123 84400 18124 84440
rect 18164 84400 18165 84440
rect 18123 84391 18165 84400
rect 18507 84440 18549 84449
rect 18507 84400 18508 84440
rect 18548 84400 18549 84440
rect 18507 84391 18549 84400
rect 18124 83768 18164 83777
rect 18028 83728 18124 83768
rect 18124 83719 18164 83728
rect 19180 83768 19220 84484
rect 19468 84449 19508 85936
rect 19563 85448 19605 85457
rect 19563 85408 19564 85448
rect 19604 85408 19605 85448
rect 19563 85399 19605 85408
rect 19467 84440 19509 84449
rect 19467 84400 19468 84440
rect 19508 84400 19509 84440
rect 19467 84391 19509 84400
rect 19180 83719 19220 83728
rect 19275 83768 19317 83777
rect 19275 83728 19276 83768
rect 19316 83728 19317 83768
rect 19275 83719 19317 83728
rect 19564 83768 19604 85399
rect 19851 84776 19893 84785
rect 19851 84736 19852 84776
rect 19892 84736 19893 84776
rect 19851 84727 19893 84736
rect 19564 83719 19604 83728
rect 18316 83516 18356 83525
rect 17836 83476 18316 83516
rect 16780 81880 17012 81920
rect 16683 80408 16725 80417
rect 16683 80368 16684 80408
rect 16724 80368 16725 80408
rect 16683 80359 16725 80368
rect 16684 79988 16724 80359
rect 16684 79939 16724 79948
rect 16875 79400 16917 79409
rect 16875 79360 16876 79400
rect 16916 79360 16917 79400
rect 16875 79351 16917 79360
rect 16396 79192 16628 79232
rect 16299 77804 16341 77813
rect 16299 77764 16300 77804
rect 16340 77764 16341 77804
rect 16299 77755 16341 77764
rect 16203 77720 16245 77729
rect 16203 77680 16204 77720
rect 16244 77680 16245 77720
rect 16203 77671 16245 77680
rect 16300 77552 16340 77561
rect 16108 77512 16300 77552
rect 16300 77503 16340 77512
rect 16396 77477 16436 79192
rect 16587 79064 16629 79073
rect 16587 79024 16588 79064
rect 16628 79024 16629 79064
rect 16587 79015 16629 79024
rect 16588 78930 16628 79015
rect 16780 78812 16820 78821
rect 16588 78772 16780 78812
rect 16588 78308 16628 78772
rect 16780 78763 16820 78772
rect 16540 78268 16628 78308
rect 16540 78266 16580 78268
rect 16540 78217 16580 78226
rect 16684 78056 16724 78065
rect 16588 78016 16684 78056
rect 16395 77468 16437 77477
rect 16395 77428 16396 77468
rect 16436 77428 16437 77468
rect 16395 77419 16437 77428
rect 16588 77384 16628 78016
rect 16684 78007 16724 78016
rect 16876 77888 16916 79351
rect 16684 77848 16916 77888
rect 16684 77720 16724 77848
rect 16684 77671 16724 77680
rect 16972 77636 17012 81880
rect 17067 77720 17109 77729
rect 17067 77680 17068 77720
rect 17108 77680 17109 77720
rect 17067 77671 17109 77680
rect 17739 77720 17781 77729
rect 17739 77680 17740 77720
rect 17780 77680 17781 77720
rect 17739 77671 17781 77680
rect 16780 77596 17012 77636
rect 16588 77344 16724 77384
rect 16492 77300 16532 77309
rect 16532 77260 16628 77300
rect 16492 77251 16532 77260
rect 16203 76964 16245 76973
rect 16203 76924 16204 76964
rect 16244 76924 16245 76964
rect 16203 76915 16245 76924
rect 16107 76712 16149 76721
rect 16107 76672 16108 76712
rect 16148 76672 16149 76712
rect 16107 76663 16149 76672
rect 16108 75965 16148 76663
rect 16107 75956 16149 75965
rect 16107 75916 16108 75956
rect 16148 75916 16149 75956
rect 16107 75907 16149 75916
rect 16012 75664 16148 75704
rect 16011 75536 16053 75545
rect 16011 75496 16012 75536
rect 16052 75496 16053 75536
rect 16011 75487 16053 75496
rect 16012 75377 16052 75487
rect 16011 75368 16053 75377
rect 16011 75328 16012 75368
rect 16052 75328 16053 75368
rect 16011 75319 16053 75328
rect 15915 73016 15957 73025
rect 15915 72976 15916 73016
rect 15956 72976 15957 73016
rect 15915 72967 15957 72976
rect 15915 71504 15957 71513
rect 15915 71464 15916 71504
rect 15956 71464 15957 71504
rect 15915 71455 15957 71464
rect 15916 71370 15956 71455
rect 16012 69236 16052 75319
rect 16108 74453 16148 75664
rect 16204 75293 16244 76915
rect 16588 76726 16628 77260
rect 16684 76889 16724 77344
rect 16683 76880 16725 76889
rect 16683 76840 16684 76880
rect 16724 76840 16725 76880
rect 16683 76831 16725 76840
rect 16780 76712 16820 77596
rect 17068 77586 17108 77671
rect 17740 77552 17780 77671
rect 16588 76677 16628 76686
rect 16684 76672 16820 76712
rect 16876 77468 16916 77477
rect 16684 76628 16724 76672
rect 16396 76588 16724 76628
rect 16203 75284 16245 75293
rect 16203 75244 16204 75284
rect 16244 75244 16245 75284
rect 16203 75235 16245 75244
rect 16300 74528 16340 74537
rect 16107 74444 16149 74453
rect 16107 74404 16108 74444
rect 16148 74404 16149 74444
rect 16107 74395 16149 74404
rect 16108 74201 16148 74395
rect 16107 74192 16149 74201
rect 16107 74152 16108 74192
rect 16148 74152 16149 74192
rect 16107 74143 16149 74152
rect 16300 73865 16340 74488
rect 16299 73856 16341 73865
rect 16299 73816 16300 73856
rect 16340 73816 16341 73856
rect 16299 73807 16341 73816
rect 16300 73709 16340 73718
rect 16204 73669 16300 73702
rect 16204 73662 16340 73669
rect 16204 73613 16244 73662
rect 16300 73660 16340 73662
rect 16203 73604 16245 73613
rect 16203 73564 16204 73604
rect 16244 73564 16245 73604
rect 16203 73555 16245 73564
rect 16204 73016 16244 73555
rect 16299 73100 16341 73109
rect 16299 73060 16300 73100
rect 16340 73060 16341 73100
rect 16396 73100 16436 76588
rect 16779 76544 16821 76553
rect 16779 76504 16780 76544
rect 16820 76504 16821 76544
rect 16779 76495 16821 76504
rect 16780 76410 16820 76495
rect 16876 76208 16916 77428
rect 17259 77468 17301 77477
rect 17259 77428 17260 77468
rect 17300 77428 17301 77468
rect 17259 77419 17301 77428
rect 17164 76712 17204 76721
rect 17260 76712 17300 77419
rect 17740 76973 17780 77512
rect 17739 76964 17781 76973
rect 17739 76924 17740 76964
rect 17780 76924 17781 76964
rect 17739 76915 17781 76924
rect 17547 76880 17589 76889
rect 17547 76840 17548 76880
rect 17588 76840 17589 76880
rect 17547 76831 17589 76840
rect 17204 76672 17300 76712
rect 16972 76544 17012 76553
rect 16972 76217 17012 76504
rect 16588 76168 16916 76208
rect 16971 76208 17013 76217
rect 16971 76168 16972 76208
rect 17012 76168 17013 76208
rect 16588 75200 16628 76168
rect 16971 76159 17013 76168
rect 16876 76040 16916 76049
rect 17164 76040 17204 76672
rect 17451 76628 17493 76637
rect 17451 76588 17452 76628
rect 17492 76588 17493 76628
rect 17451 76579 17493 76588
rect 16916 76000 17204 76040
rect 16876 75293 16916 76000
rect 17068 75797 17108 75882
rect 17260 75872 17300 75881
rect 17067 75788 17109 75797
rect 17067 75748 17068 75788
rect 17108 75748 17109 75788
rect 17067 75739 17109 75748
rect 17260 75629 17300 75832
rect 17067 75620 17109 75629
rect 17067 75580 17068 75620
rect 17108 75580 17109 75620
rect 17067 75571 17109 75580
rect 17259 75620 17301 75629
rect 17259 75580 17260 75620
rect 17300 75580 17301 75620
rect 17259 75571 17301 75580
rect 16875 75284 16917 75293
rect 16875 75244 16876 75284
rect 16916 75244 16917 75284
rect 16875 75235 16917 75244
rect 16588 73697 16628 75160
rect 16971 75200 17013 75209
rect 16971 75160 16972 75200
rect 17012 75160 17013 75200
rect 16971 75151 17013 75160
rect 16972 75066 17012 75151
rect 16780 75032 16820 75041
rect 16780 74523 16820 74992
rect 16780 74474 16820 74483
rect 16972 74612 17012 74621
rect 16972 74453 17012 74572
rect 16971 74444 17013 74453
rect 16971 74404 16972 74444
rect 17012 74404 17013 74444
rect 16971 74395 17013 74404
rect 16587 73688 16629 73697
rect 16587 73648 16588 73688
rect 16628 73648 16629 73688
rect 16587 73639 16629 73648
rect 16492 73520 16532 73529
rect 16532 73480 16724 73520
rect 16492 73471 16532 73480
rect 16396 73060 16532 73100
rect 16299 73051 16341 73060
rect 16107 72008 16149 72017
rect 16107 71968 16108 72008
rect 16148 71968 16149 72008
rect 16107 71959 16149 71968
rect 16108 70664 16148 71959
rect 16204 70673 16244 72976
rect 16108 70589 16148 70624
rect 16203 70664 16245 70673
rect 16203 70624 16204 70664
rect 16244 70624 16245 70664
rect 16203 70615 16245 70624
rect 16107 70580 16149 70589
rect 16107 70540 16108 70580
rect 16148 70540 16149 70580
rect 16107 70531 16149 70540
rect 16108 70500 16148 70531
rect 16300 70076 16340 73051
rect 16396 72764 16436 72773
rect 16396 72353 16436 72724
rect 16395 72344 16437 72353
rect 16395 72304 16396 72344
rect 16436 72304 16437 72344
rect 16395 72295 16437 72304
rect 16204 70036 16340 70076
rect 16107 69908 16149 69917
rect 16107 69868 16108 69908
rect 16148 69868 16149 69908
rect 16107 69859 16149 69868
rect 16204 69908 16244 70036
rect 16108 69774 16148 69859
rect 16204 69833 16244 69868
rect 16203 69824 16245 69833
rect 16203 69784 16204 69824
rect 16244 69784 16245 69824
rect 16203 69775 16245 69784
rect 16108 69245 16148 69289
rect 16107 69236 16149 69245
rect 16012 69196 16108 69236
rect 16148 69196 16149 69236
rect 16107 69194 16149 69196
rect 16107 69187 16108 69194
rect 16148 69187 16149 69194
rect 16108 69145 16148 69154
rect 16203 68228 16245 68237
rect 16203 68188 16204 68228
rect 16244 68188 16245 68228
rect 16203 68179 16245 68188
rect 15915 67892 15957 67901
rect 15915 67852 15916 67892
rect 15956 67852 15957 67892
rect 15915 67843 15957 67852
rect 15916 67758 15956 67843
rect 16204 67640 16244 68179
rect 16204 67591 16244 67600
rect 16300 67620 16340 67651
rect 16300 67565 16340 67580
rect 16299 67556 16341 67565
rect 16299 67516 16300 67556
rect 16340 67516 16341 67556
rect 16299 67507 16341 67516
rect 15915 67304 15957 67313
rect 15915 67264 15916 67304
rect 15956 67264 15957 67304
rect 15915 67255 15957 67264
rect 16395 67304 16437 67313
rect 16395 67264 16396 67304
rect 16436 67264 16437 67304
rect 16395 67255 16437 67264
rect 15819 66884 15861 66893
rect 15819 66844 15820 66884
rect 15860 66844 15861 66884
rect 15819 66835 15861 66844
rect 15723 64616 15765 64625
rect 15723 64576 15724 64616
rect 15764 64576 15765 64616
rect 15723 64567 15765 64576
rect 15724 64482 15764 64567
rect 15628 64240 15764 64280
rect 14955 63895 14997 63904
rect 15436 63890 15476 63899
rect 15628 64028 15668 64037
rect 15628 63869 15668 63988
rect 14859 63860 14901 63869
rect 14859 63820 14860 63860
rect 14900 63820 14901 63860
rect 14859 63811 14901 63820
rect 15627 63860 15669 63869
rect 15627 63820 15628 63860
rect 15668 63820 15669 63860
rect 15627 63811 15669 63820
rect 14763 62264 14805 62273
rect 14763 62224 14764 62264
rect 14804 62224 14805 62264
rect 14763 62215 14805 62224
rect 14860 60761 14900 63811
rect 15052 63104 15092 63115
rect 15052 63029 15092 63064
rect 15147 63104 15189 63113
rect 15147 63064 15148 63104
rect 15188 63064 15189 63104
rect 15147 63055 15189 63064
rect 15531 63104 15573 63113
rect 15531 63064 15532 63104
rect 15572 63064 15573 63104
rect 15531 63055 15573 63064
rect 15051 63020 15093 63029
rect 15051 62980 15052 63020
rect 15092 62980 15093 63020
rect 15051 62971 15093 62980
rect 15051 62852 15093 62861
rect 15051 62812 15052 62852
rect 15092 62812 15093 62852
rect 15051 62803 15093 62812
rect 14956 62432 14996 62441
rect 14956 62273 14996 62392
rect 14955 62264 14997 62273
rect 14955 62224 14956 62264
rect 14996 62224 14997 62264
rect 14955 62215 14997 62224
rect 14955 60836 14997 60845
rect 14955 60796 14956 60836
rect 14996 60796 14997 60836
rect 14955 60787 14997 60796
rect 14859 60752 14901 60761
rect 14859 60712 14860 60752
rect 14900 60712 14901 60752
rect 14859 60703 14901 60712
rect 14764 60668 14804 60677
rect 14667 60584 14709 60593
rect 14667 60544 14668 60584
rect 14708 60544 14709 60584
rect 14667 60535 14709 60544
rect 14667 60416 14709 60425
rect 14667 60376 14668 60416
rect 14708 60376 14709 60416
rect 14667 60367 14709 60376
rect 14668 60005 14708 60367
rect 14764 60094 14804 60628
rect 14764 60045 14804 60054
rect 14667 59996 14709 60005
rect 14667 59956 14668 59996
rect 14708 59956 14709 59996
rect 14667 59947 14709 59956
rect 14956 59996 14996 60787
rect 15052 60425 15092 62803
rect 15148 61097 15188 63055
rect 15532 62970 15572 63055
rect 15244 62936 15284 62945
rect 15284 62896 15476 62936
rect 15244 62887 15284 62896
rect 15436 62427 15476 62896
rect 15436 62378 15476 62387
rect 15628 62516 15668 62525
rect 15628 62357 15668 62476
rect 15627 62348 15669 62357
rect 15627 62308 15628 62348
rect 15668 62308 15669 62348
rect 15627 62299 15669 62308
rect 15627 61760 15669 61769
rect 15627 61720 15628 61760
rect 15668 61720 15669 61760
rect 15627 61711 15669 61720
rect 15147 61088 15189 61097
rect 15147 61048 15148 61088
rect 15188 61048 15189 61088
rect 15147 61039 15189 61048
rect 15051 60416 15093 60425
rect 15051 60376 15052 60416
rect 15092 60376 15093 60416
rect 15051 60367 15093 60376
rect 15628 60173 15668 61711
rect 15627 60164 15669 60173
rect 15627 60124 15628 60164
rect 15668 60124 15669 60164
rect 15627 60115 15669 60124
rect 15051 60080 15093 60089
rect 15148 60080 15188 60089
rect 15051 60040 15052 60080
rect 15092 60040 15148 60080
rect 15051 60031 15093 60040
rect 15148 60031 15188 60040
rect 15244 60080 15284 60089
rect 15435 60080 15477 60089
rect 15284 60040 15291 60080
rect 15244 60031 15291 60040
rect 15435 60040 15436 60080
rect 15476 60040 15477 60080
rect 15435 60031 15477 60040
rect 14956 59947 14996 59956
rect 14956 58568 14996 58577
rect 14763 58232 14805 58241
rect 14763 58192 14764 58232
rect 14804 58192 14805 58232
rect 14763 58183 14805 58192
rect 14667 57896 14709 57905
rect 14667 57856 14668 57896
rect 14708 57856 14709 57896
rect 14667 57847 14709 57856
rect 14668 56981 14708 57847
rect 14764 57056 14804 58183
rect 14956 57149 14996 58528
rect 14955 57140 14997 57149
rect 14955 57100 14956 57140
rect 14996 57100 14997 57140
rect 14955 57091 14997 57100
rect 14804 57016 14900 57056
rect 14764 57007 14804 57016
rect 14667 56972 14709 56981
rect 14667 56932 14668 56972
rect 14708 56932 14709 56972
rect 14667 56923 14709 56932
rect 14668 56561 14708 56923
rect 14667 56552 14709 56561
rect 14667 56512 14668 56552
rect 14708 56512 14709 56552
rect 14667 56503 14709 56512
rect 14667 56384 14709 56393
rect 14667 56344 14668 56384
rect 14708 56344 14709 56384
rect 14667 56335 14709 56344
rect 14860 56384 14900 57016
rect 14860 56335 14900 56344
rect 14668 56141 14708 56335
rect 14667 56132 14709 56141
rect 14667 56092 14668 56132
rect 14708 56092 14709 56132
rect 14667 56083 14709 56092
rect 14668 55376 14708 55385
rect 14708 55336 14804 55376
rect 14668 55327 14708 55336
rect 14667 53948 14709 53957
rect 14667 53908 14668 53948
rect 14708 53908 14709 53948
rect 14667 53899 14709 53908
rect 14668 53814 14708 53899
rect 14764 53360 14804 55336
rect 14860 54872 14900 54881
rect 14860 54377 14900 54832
rect 14859 54368 14901 54377
rect 14859 54328 14860 54368
rect 14900 54328 14901 54368
rect 14859 54319 14901 54328
rect 14860 53444 14900 53453
rect 14900 53404 14996 53444
rect 14860 53395 14900 53404
rect 14716 53350 14804 53360
rect 14756 53320 14804 53350
rect 14716 53301 14756 53310
rect 14763 52772 14805 52781
rect 14763 52732 14764 52772
rect 14804 52732 14805 52772
rect 14763 52723 14805 52732
rect 14668 52520 14708 52529
rect 14668 51773 14708 52480
rect 14764 51848 14804 52723
rect 14667 51764 14709 51773
rect 14667 51724 14668 51764
rect 14708 51724 14709 51764
rect 14764 51764 14804 51808
rect 14859 51764 14901 51773
rect 14764 51724 14860 51764
rect 14900 51724 14901 51764
rect 14667 51715 14709 51724
rect 14859 51715 14901 51724
rect 14571 51008 14613 51017
rect 14571 50968 14572 51008
rect 14612 50968 14613 51008
rect 14571 50959 14613 50968
rect 14668 51008 14708 51017
rect 14571 50840 14613 50849
rect 14571 50800 14572 50840
rect 14612 50800 14613 50840
rect 14571 50791 14613 50800
rect 14475 50588 14517 50597
rect 14475 50548 14476 50588
rect 14516 50548 14517 50588
rect 14475 50539 14517 50548
rect 14379 49748 14421 49757
rect 14379 49708 14380 49748
rect 14420 49708 14421 49748
rect 14379 49699 14421 49708
rect 14380 49589 14420 49620
rect 14379 49580 14421 49589
rect 14379 49540 14380 49580
rect 14420 49540 14421 49580
rect 14379 49531 14421 49540
rect 14380 49496 14420 49531
rect 14283 48236 14325 48245
rect 14283 48196 14284 48236
rect 14324 48196 14325 48236
rect 14283 48187 14325 48196
rect 14283 47900 14325 47909
rect 14283 47860 14284 47900
rect 14324 47860 14325 47900
rect 14283 47851 14325 47860
rect 14284 47766 14324 47851
rect 14380 46817 14420 49456
rect 14475 49496 14517 49505
rect 14475 49456 14476 49496
rect 14516 49456 14517 49496
rect 14475 49447 14517 49456
rect 14476 49362 14516 49447
rect 14379 46808 14421 46817
rect 14379 46768 14380 46808
rect 14420 46768 14421 46808
rect 14379 46759 14421 46768
rect 14572 46640 14612 50791
rect 14668 49589 14708 50968
rect 14764 51008 14804 51017
rect 14764 50429 14804 50968
rect 14763 50420 14805 50429
rect 14763 50380 14764 50420
rect 14804 50380 14805 50420
rect 14763 50371 14805 50380
rect 14956 50093 14996 53404
rect 14955 50084 14997 50093
rect 14955 50044 14956 50084
rect 14996 50044 14997 50084
rect 14955 50035 14997 50044
rect 15052 49916 15092 60031
rect 15251 59912 15291 60031
rect 15436 59946 15476 60031
rect 15244 59872 15291 59912
rect 15340 59912 15380 59921
rect 15244 59576 15284 59872
rect 15340 59744 15380 59872
rect 15340 59704 15668 59744
rect 15436 59576 15476 59585
rect 15244 59536 15436 59576
rect 15436 59417 15476 59536
rect 15244 59408 15284 59417
rect 15244 58988 15284 59368
rect 15435 59408 15477 59417
rect 15435 59368 15436 59408
rect 15476 59368 15477 59408
rect 15435 59359 15477 59368
rect 15628 59408 15668 59704
rect 15724 59576 15764 64240
rect 15820 61592 15860 61601
rect 15820 61349 15860 61552
rect 15819 61340 15861 61349
rect 15819 61300 15820 61340
rect 15860 61300 15861 61340
rect 15819 61291 15861 61300
rect 15916 59669 15956 67255
rect 16299 65624 16341 65633
rect 16299 65584 16300 65624
rect 16340 65584 16341 65624
rect 16299 65575 16341 65584
rect 16300 65490 16340 65575
rect 16299 64616 16341 64625
rect 16299 64576 16300 64616
rect 16340 64576 16341 64616
rect 16299 64567 16341 64576
rect 16300 61937 16340 64567
rect 16299 61928 16341 61937
rect 16299 61888 16300 61928
rect 16340 61888 16341 61928
rect 16299 61879 16341 61888
rect 16203 61592 16245 61601
rect 16203 61552 16204 61592
rect 16244 61552 16245 61592
rect 16203 61543 16245 61552
rect 16204 61458 16244 61543
rect 16012 61424 16052 61433
rect 16012 60920 16052 61384
rect 16108 60920 16148 60929
rect 16012 60880 16108 60920
rect 16108 60871 16148 60880
rect 16204 60920 16244 60929
rect 16204 60593 16244 60880
rect 16203 60584 16245 60593
rect 16203 60544 16204 60584
rect 16244 60544 16245 60584
rect 16203 60535 16245 60544
rect 16012 60080 16052 60091
rect 16012 60005 16052 60040
rect 16107 60080 16149 60089
rect 16107 60040 16108 60080
rect 16148 60040 16149 60080
rect 16107 60031 16149 60040
rect 16011 59996 16053 60005
rect 16011 59956 16012 59996
rect 16052 59956 16053 59996
rect 16011 59947 16053 59956
rect 16108 59669 16148 60031
rect 15915 59660 15957 59669
rect 15915 59620 15916 59660
rect 15956 59620 15957 59660
rect 16108 59660 16154 59669
rect 16108 59620 16113 59660
rect 16153 59620 16154 59660
rect 15915 59611 15957 59620
rect 16112 59611 16154 59620
rect 15724 59536 15860 59576
rect 15628 59359 15668 59368
rect 15724 59393 15764 59402
rect 15724 59165 15764 59353
rect 15628 59156 15668 59165
rect 15244 58948 15476 58988
rect 15339 58820 15381 58829
rect 15339 58780 15340 58820
rect 15380 58780 15381 58820
rect 15339 58771 15381 58780
rect 15340 58686 15380 58771
rect 15436 58568 15476 58948
rect 15532 58568 15572 58577
rect 15436 58528 15532 58568
rect 15148 58400 15188 58409
rect 15148 57728 15188 58360
rect 15244 57905 15284 57990
rect 15243 57896 15285 57905
rect 15243 57856 15244 57896
rect 15284 57856 15285 57896
rect 15243 57847 15285 57856
rect 15148 57688 15284 57728
rect 15244 57070 15284 57688
rect 15436 57644 15476 57653
rect 15244 57021 15284 57030
rect 15340 57604 15436 57644
rect 15340 56379 15380 57604
rect 15436 57595 15476 57604
rect 15435 56888 15477 56897
rect 15435 56848 15436 56888
rect 15476 56848 15477 56888
rect 15435 56839 15477 56848
rect 15436 56754 15476 56839
rect 15532 56636 15572 58528
rect 15628 58241 15668 59116
rect 15723 59156 15765 59165
rect 15723 59116 15724 59156
rect 15764 59116 15765 59156
rect 15723 59107 15765 59116
rect 15627 58232 15669 58241
rect 15627 58192 15628 58232
rect 15668 58192 15669 58232
rect 15627 58183 15669 58192
rect 15627 58064 15669 58073
rect 15627 58024 15628 58064
rect 15668 58024 15669 58064
rect 15627 58015 15669 58024
rect 15628 57980 15668 58015
rect 15628 57929 15668 57940
rect 15724 57896 15764 57905
rect 15820 57896 15860 59536
rect 15915 59408 15957 59417
rect 15915 59368 15916 59408
rect 15956 59368 15957 59408
rect 15915 59359 15957 59368
rect 16012 59408 16052 59417
rect 15916 59274 15956 59359
rect 16012 58073 16052 59368
rect 16113 59408 16153 59611
rect 16113 59359 16153 59368
rect 16203 58988 16245 58997
rect 16203 58948 16204 58988
rect 16244 58948 16245 58988
rect 16203 58939 16245 58948
rect 16011 58064 16053 58073
rect 16011 58024 16012 58064
rect 16052 58024 16053 58064
rect 16011 58015 16053 58024
rect 15916 57896 15956 57905
rect 15820 57856 15916 57896
rect 15627 57476 15669 57485
rect 15627 57436 15628 57476
rect 15668 57436 15669 57476
rect 15627 57427 15669 57436
rect 15628 57065 15668 57427
rect 15627 57056 15669 57065
rect 15627 57016 15628 57056
rect 15668 57016 15669 57056
rect 15627 57007 15669 57016
rect 15340 56330 15380 56339
rect 15436 56596 15572 56636
rect 15436 56216 15476 56596
rect 15244 56176 15476 56216
rect 15532 56468 15572 56477
rect 15147 54200 15189 54209
rect 15244 54200 15284 56176
rect 15532 55460 15572 56428
rect 15436 55420 15572 55460
rect 15340 54209 15380 54294
rect 15147 54160 15148 54200
rect 15188 54160 15284 54200
rect 15339 54200 15381 54209
rect 15339 54160 15340 54200
rect 15380 54160 15381 54200
rect 15147 54151 15189 54160
rect 15339 54151 15381 54160
rect 15148 54032 15188 54041
rect 15340 54032 15380 54043
rect 15188 53992 15284 54023
rect 15148 53983 15284 53992
rect 15147 53864 15189 53873
rect 15147 53824 15148 53864
rect 15188 53824 15189 53864
rect 15147 53815 15189 53824
rect 15148 51857 15188 53815
rect 15244 53537 15284 53983
rect 15340 53957 15380 53992
rect 15339 53948 15381 53957
rect 15339 53908 15340 53948
rect 15380 53908 15381 53948
rect 15339 53899 15381 53908
rect 15436 53780 15476 55420
rect 15628 55208 15668 57007
rect 15724 55889 15764 57856
rect 15723 55880 15765 55889
rect 15723 55840 15724 55880
rect 15764 55840 15765 55880
rect 15723 55831 15765 55840
rect 15724 55553 15764 55638
rect 15819 55628 15861 55637
rect 15819 55588 15820 55628
rect 15860 55588 15861 55628
rect 15819 55579 15861 55588
rect 15723 55544 15765 55553
rect 15723 55504 15724 55544
rect 15764 55504 15765 55544
rect 15723 55495 15765 55504
rect 15820 55376 15860 55579
rect 15340 53740 15476 53780
rect 15532 55168 15668 55208
rect 15724 55336 15860 55376
rect 15532 54032 15572 55168
rect 15243 53528 15285 53537
rect 15243 53488 15244 53528
rect 15284 53488 15285 53528
rect 15243 53479 15285 53488
rect 15244 53394 15284 53479
rect 15147 51848 15189 51857
rect 15147 51808 15148 51848
rect 15188 51808 15189 51848
rect 15147 51799 15189 51808
rect 15147 50672 15189 50681
rect 15147 50632 15148 50672
rect 15188 50632 15189 50672
rect 15147 50623 15189 50632
rect 14860 49876 15092 49916
rect 14763 49748 14805 49757
rect 14763 49708 14764 49748
rect 14804 49708 14805 49748
rect 14763 49699 14805 49708
rect 14667 49580 14709 49589
rect 14667 49540 14668 49580
rect 14708 49540 14709 49580
rect 14667 49531 14709 49540
rect 14764 47984 14804 49699
rect 14764 46733 14804 47944
rect 14763 46724 14805 46733
rect 14763 46684 14764 46724
rect 14804 46684 14805 46724
rect 14763 46675 14805 46684
rect 14572 46600 14708 46640
rect 14380 46477 14420 46486
rect 14284 45968 14324 45977
rect 14380 45968 14420 46437
rect 14571 46388 14613 46397
rect 14571 46348 14572 46388
rect 14612 46348 14613 46388
rect 14571 46339 14613 46348
rect 14572 46254 14612 46339
rect 14668 46136 14708 46600
rect 14572 46096 14708 46136
rect 14324 45928 14420 45968
rect 14476 45968 14516 45977
rect 14284 45919 14324 45928
rect 14380 44960 14420 44969
rect 14188 44920 14380 44960
rect 14380 44911 14420 44920
rect 13707 44876 13749 44885
rect 13707 44836 13708 44876
rect 13748 44836 13749 44876
rect 13707 44827 13749 44836
rect 13899 44708 13941 44717
rect 13899 44668 13900 44708
rect 13940 44668 13941 44708
rect 13899 44659 13941 44668
rect 13803 44624 13845 44633
rect 13803 44584 13804 44624
rect 13844 44584 13845 44624
rect 13803 44575 13845 44584
rect 13515 44500 13556 44540
rect 13707 44540 13749 44549
rect 13707 44500 13708 44540
rect 13748 44500 13749 44540
rect 13228 44416 13364 44456
rect 13228 44288 13268 44297
rect 13228 44045 13268 44248
rect 13227 44036 13269 44045
rect 13227 43996 13228 44036
rect 13268 43996 13269 44036
rect 13227 43987 13269 43996
rect 12940 43660 13172 43700
rect 12843 43364 12885 43373
rect 12843 43324 12844 43364
rect 12884 43324 12885 43364
rect 12843 43315 12885 43324
rect 12747 43280 12789 43289
rect 12747 43240 12748 43280
rect 12788 43240 12789 43280
rect 12747 43231 12789 43240
rect 12748 43146 12788 43231
rect 12747 42776 12789 42785
rect 12747 42736 12748 42776
rect 12788 42736 12789 42776
rect 12747 42727 12789 42736
rect 12748 42642 12788 42727
rect 12843 42020 12885 42029
rect 12843 41980 12844 42020
rect 12884 41980 12885 42020
rect 12843 41971 12885 41980
rect 12747 41936 12789 41945
rect 12747 41896 12748 41936
rect 12788 41896 12789 41936
rect 12747 41887 12789 41896
rect 12748 41802 12788 41887
rect 12844 41886 12884 41971
rect 12652 40552 12788 40592
rect 12651 40424 12693 40433
rect 12651 40384 12652 40424
rect 12692 40384 12693 40424
rect 12651 40375 12693 40384
rect 12652 40290 12692 40375
rect 12651 40172 12693 40181
rect 12651 40132 12652 40172
rect 12692 40132 12693 40172
rect 12651 40123 12693 40132
rect 12459 39752 12501 39761
rect 12459 39712 12460 39752
rect 12500 39712 12501 39752
rect 12459 39703 12501 39712
rect 12556 39752 12596 39761
rect 12460 39618 12500 39703
rect 12556 39593 12596 39712
rect 12555 39584 12597 39593
rect 12555 39544 12556 39584
rect 12596 39544 12597 39584
rect 12555 39535 12597 39544
rect 12459 39080 12501 39089
rect 12459 39040 12460 39080
rect 12500 39040 12501 39080
rect 12459 39031 12501 39040
rect 12460 38946 12500 39031
rect 12652 38912 12692 40123
rect 12652 38828 12692 38872
rect 12172 38704 12404 38744
rect 12556 38788 12692 38828
rect 12075 38408 12117 38417
rect 12075 38368 12076 38408
rect 12116 38368 12117 38408
rect 12075 38359 12117 38368
rect 11884 38324 11924 38333
rect 11884 38081 11924 38284
rect 11883 38072 11925 38081
rect 11883 38032 11884 38072
rect 11924 38032 11925 38072
rect 11883 38023 11925 38032
rect 12076 37904 12116 38359
rect 11692 37780 11828 37820
rect 11884 37864 12116 37904
rect 11692 36317 11732 37780
rect 11884 37409 11924 37864
rect 12172 37820 12212 38704
rect 11980 37780 12212 37820
rect 12268 38240 12308 38249
rect 11883 37400 11925 37409
rect 11883 37360 11884 37400
rect 11924 37360 11925 37400
rect 11883 37351 11925 37360
rect 11787 37316 11829 37325
rect 11787 37276 11788 37316
rect 11828 37276 11829 37316
rect 11787 37267 11829 37276
rect 11691 36308 11733 36317
rect 11691 36268 11692 36308
rect 11732 36268 11733 36308
rect 11691 36259 11733 36268
rect 11691 35972 11733 35981
rect 11691 35932 11692 35972
rect 11732 35932 11733 35972
rect 11691 35923 11733 35932
rect 11692 35216 11732 35923
rect 11788 35888 11828 37267
rect 11884 37266 11924 37351
rect 11980 36233 12020 37780
rect 12076 37652 12116 37661
rect 12268 37652 12308 38200
rect 12116 37612 12308 37652
rect 12364 38240 12404 38249
rect 12076 37603 12116 37612
rect 12172 37400 12308 37409
rect 12172 37369 12268 37400
rect 12172 37325 12212 37369
rect 12268 37351 12308 37360
rect 12171 37316 12213 37325
rect 12171 37276 12172 37316
rect 12212 37276 12213 37316
rect 12171 37267 12213 37276
rect 12364 36569 12404 38200
rect 12363 36560 12405 36569
rect 12363 36520 12364 36560
rect 12404 36520 12405 36560
rect 12363 36511 12405 36520
rect 11979 36224 12021 36233
rect 11979 36184 11980 36224
rect 12020 36184 12021 36224
rect 11979 36175 12021 36184
rect 12171 36056 12213 36065
rect 12171 36016 12172 36056
rect 12212 36016 12213 36056
rect 12171 36007 12213 36016
rect 11788 35477 11828 35848
rect 11979 35888 12021 35897
rect 11979 35848 11980 35888
rect 12020 35848 12021 35888
rect 11979 35839 12021 35848
rect 12172 35888 12212 36007
rect 12556 35972 12596 38788
rect 12748 38744 12788 40552
rect 12940 40424 12980 43660
rect 13324 43616 13364 44416
rect 13515 44372 13555 44500
rect 13707 44491 13749 44500
rect 13612 44456 13652 44465
rect 13515 44332 13556 44372
rect 13419 44204 13461 44213
rect 13419 44164 13420 44204
rect 13460 44164 13461 44204
rect 13419 44155 13461 44164
rect 13420 44120 13460 44155
rect 13420 44069 13460 44080
rect 13132 43576 13364 43616
rect 13419 43616 13461 43625
rect 13419 43576 13420 43616
rect 13460 43576 13461 43616
rect 13132 43448 13172 43576
rect 13419 43567 13461 43576
rect 13323 43448 13365 43457
rect 13132 43399 13172 43408
rect 13228 43427 13268 43436
rect 13323 43408 13324 43448
rect 13364 43408 13365 43448
rect 13323 43399 13365 43408
rect 13420 43448 13460 43567
rect 13420 43399 13460 43408
rect 13228 43373 13268 43387
rect 13227 43364 13269 43373
rect 13227 43324 13228 43364
rect 13268 43324 13269 43364
rect 13227 43315 13269 43324
rect 13228 43292 13268 43315
rect 13324 43314 13364 43399
rect 13227 42776 13269 42785
rect 13227 42736 13228 42776
rect 13268 42736 13269 42776
rect 13227 42727 13269 42736
rect 13035 42020 13077 42029
rect 13035 41980 13036 42020
rect 13076 41980 13077 42020
rect 13035 41971 13077 41980
rect 12844 40384 12980 40424
rect 12844 40013 12884 40384
rect 12939 40256 12981 40265
rect 12939 40216 12940 40256
rect 12980 40216 12981 40256
rect 12939 40207 12981 40216
rect 12843 40004 12885 40013
rect 12843 39964 12844 40004
rect 12884 39964 12885 40004
rect 12843 39955 12885 39964
rect 12940 39677 12980 40207
rect 13036 39752 13076 41971
rect 13228 41693 13268 42727
rect 13516 42272 13556 44332
rect 13612 43448 13652 44416
rect 13708 44120 13748 44491
rect 13804 44288 13844 44575
rect 13804 44239 13844 44248
rect 13900 44288 13940 44659
rect 13995 44624 14037 44633
rect 13995 44584 13996 44624
rect 14036 44584 14037 44624
rect 13995 44575 14037 44584
rect 13900 44239 13940 44248
rect 13708 44080 13844 44120
rect 13708 43448 13748 43457
rect 13612 43408 13708 43448
rect 13708 43399 13748 43408
rect 13611 43280 13653 43289
rect 13804 43280 13844 44080
rect 13996 43961 14036 44575
rect 14091 44540 14133 44549
rect 14091 44500 14092 44540
rect 14132 44500 14133 44540
rect 14091 44491 14133 44500
rect 14092 44288 14132 44491
rect 14283 44456 14325 44465
rect 14283 44416 14284 44456
rect 14324 44416 14325 44456
rect 14283 44407 14325 44416
rect 14092 44239 14132 44248
rect 14188 44288 14228 44297
rect 14188 44120 14228 44248
rect 14284 44288 14324 44407
rect 14284 44213 14324 44248
rect 14379 44288 14421 44297
rect 14379 44248 14380 44288
rect 14420 44248 14421 44288
rect 14379 44239 14421 44248
rect 14283 44204 14325 44213
rect 14283 44164 14284 44204
rect 14324 44164 14325 44204
rect 14283 44155 14325 44164
rect 14284 44124 14324 44155
rect 14380 44154 14420 44239
rect 14092 44080 14228 44120
rect 13995 43952 14037 43961
rect 13995 43912 13996 43952
rect 14036 43912 14037 43952
rect 13995 43903 14037 43912
rect 13996 43448 14036 43903
rect 14092 43625 14132 44080
rect 14187 43952 14229 43961
rect 14187 43912 14188 43952
rect 14228 43912 14229 43952
rect 14187 43903 14229 43912
rect 14091 43616 14133 43625
rect 14091 43576 14092 43616
rect 14132 43576 14133 43616
rect 14091 43567 14133 43576
rect 14092 43448 14132 43457
rect 13996 43408 14092 43448
rect 14092 43399 14132 43408
rect 14188 43448 14228 43903
rect 14476 43457 14516 45928
rect 14188 43399 14228 43408
rect 14284 43448 14324 43457
rect 13611 43240 13612 43280
rect 13652 43240 13844 43280
rect 13900 43280 13940 43289
rect 14284 43280 14324 43408
rect 14475 43448 14517 43457
rect 14475 43408 14476 43448
rect 14516 43408 14517 43448
rect 14475 43399 14517 43408
rect 13940 43240 14324 43280
rect 14379 43280 14421 43289
rect 14379 43240 14380 43280
rect 14420 43240 14421 43280
rect 13611 43231 13653 43240
rect 13900 43231 13940 43240
rect 14379 43231 14421 43240
rect 13612 43146 13652 43231
rect 14380 43146 14420 43231
rect 13995 42776 14037 42785
rect 13995 42736 13996 42776
rect 14036 42736 14037 42776
rect 13995 42727 14037 42736
rect 14572 42776 14612 46096
rect 14763 46052 14805 46061
rect 14763 46012 14764 46052
rect 14804 46012 14805 46052
rect 14763 46003 14805 46012
rect 14668 45800 14708 45809
rect 14668 44633 14708 45760
rect 14764 45800 14804 46003
rect 14764 45751 14804 45760
rect 14860 45128 14900 49876
rect 15051 49580 15093 49589
rect 15051 49540 15052 49580
rect 15092 49540 15093 49580
rect 15051 49531 15093 49540
rect 15052 49496 15092 49531
rect 15052 49445 15092 49456
rect 15148 49076 15188 50623
rect 15243 49748 15285 49757
rect 15243 49708 15244 49748
rect 15284 49708 15285 49748
rect 15243 49699 15285 49708
rect 15244 49614 15284 49699
rect 15243 49496 15285 49505
rect 15243 49456 15244 49496
rect 15284 49456 15285 49496
rect 15243 49447 15285 49456
rect 15244 49362 15284 49447
rect 15340 49253 15380 53740
rect 15435 53612 15477 53621
rect 15435 53572 15436 53612
rect 15476 53572 15477 53612
rect 15435 53563 15477 53572
rect 15436 53360 15476 53563
rect 15436 53311 15476 53320
rect 15532 51689 15572 53992
rect 15628 54032 15668 54041
rect 15628 53873 15668 53992
rect 15724 54032 15764 55336
rect 15916 55217 15956 57856
rect 16107 55544 16149 55553
rect 16107 55504 16108 55544
rect 16148 55504 16149 55544
rect 16107 55495 16149 55504
rect 15915 55208 15957 55217
rect 15915 55168 15916 55208
rect 15956 55168 15957 55208
rect 15915 55159 15957 55168
rect 15915 55040 15957 55049
rect 15915 55000 15916 55040
rect 15956 55000 15957 55040
rect 15915 54991 15957 55000
rect 15724 53983 15764 53992
rect 15627 53864 15669 53873
rect 15627 53824 15628 53864
rect 15668 53824 15669 53864
rect 15627 53815 15669 53824
rect 15820 53864 15860 53873
rect 15627 53696 15669 53705
rect 15627 53656 15628 53696
rect 15668 53656 15669 53696
rect 15627 53647 15669 53656
rect 15531 51680 15573 51689
rect 15531 51640 15532 51680
rect 15572 51640 15573 51680
rect 15531 51631 15573 51640
rect 15531 51428 15573 51437
rect 15531 51388 15532 51428
rect 15572 51388 15573 51428
rect 15531 51379 15573 51388
rect 15532 51008 15572 51379
rect 15532 50959 15572 50968
rect 15628 50765 15668 53647
rect 15820 53369 15860 53824
rect 15819 53360 15861 53369
rect 15819 53320 15820 53360
rect 15860 53320 15861 53360
rect 15819 53311 15861 53320
rect 15723 53192 15765 53201
rect 15723 53152 15724 53192
rect 15764 53152 15765 53192
rect 15723 53143 15765 53152
rect 15627 50756 15669 50765
rect 15627 50716 15628 50756
rect 15668 50716 15669 50756
rect 15627 50707 15669 50716
rect 15531 50504 15573 50513
rect 15628 50504 15668 50707
rect 15724 50681 15764 53143
rect 15819 52940 15861 52949
rect 15819 52900 15820 52940
rect 15860 52900 15861 52940
rect 15819 52891 15861 52900
rect 15820 52016 15860 52891
rect 15916 52688 15956 54991
rect 16108 54872 16148 55495
rect 16011 53948 16053 53957
rect 16011 53908 16012 53948
rect 16052 53908 16053 53948
rect 16011 53899 16053 53908
rect 16012 53814 16052 53899
rect 16108 53621 16148 54832
rect 16204 54200 16244 58939
rect 16299 57980 16341 57989
rect 16299 57940 16300 57980
rect 16340 57940 16341 57980
rect 16299 57931 16341 57940
rect 16300 57065 16340 57931
rect 16299 57056 16341 57065
rect 16299 57016 16300 57056
rect 16340 57016 16341 57056
rect 16299 57007 16341 57016
rect 16300 56922 16340 57007
rect 16396 56645 16436 67255
rect 16492 62609 16532 73060
rect 16684 73016 16724 73480
rect 16684 72967 16724 72976
rect 16780 73016 16820 73025
rect 16780 72428 16820 72976
rect 16588 72388 16820 72428
rect 16588 70001 16628 72388
rect 16971 72344 17013 72353
rect 16780 72304 16972 72344
rect 17012 72304 17013 72344
rect 16780 72176 16820 72304
rect 16971 72295 17013 72304
rect 16780 72127 16820 72136
rect 16876 72156 17012 72176
rect 16916 72136 17012 72156
rect 16876 72107 16916 72116
rect 16683 71504 16725 71513
rect 16683 71464 16684 71504
rect 16724 71464 16725 71504
rect 16683 71455 16725 71464
rect 16587 69992 16629 70001
rect 16587 69952 16588 69992
rect 16628 69952 16629 69992
rect 16587 69943 16629 69952
rect 16684 69992 16724 71455
rect 16972 70580 17012 72136
rect 16684 68993 16724 69952
rect 16876 70540 17012 70580
rect 16876 69161 16916 70540
rect 16875 69152 16917 69161
rect 16875 69112 16876 69152
rect 16916 69112 16917 69152
rect 16875 69103 16917 69112
rect 16683 68984 16725 68993
rect 16683 68944 16684 68984
rect 16724 68944 16725 68984
rect 16683 68935 16725 68944
rect 16971 68984 17013 68993
rect 16971 68944 16972 68984
rect 17012 68944 17013 68984
rect 16971 68935 17013 68944
rect 16587 68480 16629 68489
rect 16587 68440 16588 68480
rect 16628 68440 16629 68480
rect 16587 68431 16629 68440
rect 16972 68480 17012 68935
rect 16588 67649 16628 68431
rect 16972 68321 17012 68440
rect 16971 68312 17013 68321
rect 16971 68272 16972 68312
rect 17012 68272 17013 68312
rect 16971 68263 17013 68272
rect 16779 68060 16821 68069
rect 16779 68020 16780 68060
rect 16820 68020 16821 68060
rect 16779 68011 16821 68020
rect 16587 67640 16629 67649
rect 16587 67600 16588 67640
rect 16628 67600 16629 67640
rect 16587 67591 16629 67600
rect 16684 67640 16724 67651
rect 16684 67565 16724 67600
rect 16780 67640 16820 68011
rect 16971 67724 17013 67733
rect 16971 67684 16972 67724
rect 17012 67684 17013 67724
rect 16971 67675 17013 67684
rect 16683 67556 16725 67565
rect 16683 67516 16684 67556
rect 16724 67516 16725 67556
rect 16683 67507 16725 67516
rect 16684 67061 16724 67507
rect 16780 67313 16820 67600
rect 16779 67304 16821 67313
rect 16779 67264 16780 67304
rect 16820 67264 16821 67304
rect 16779 67255 16821 67264
rect 16875 67220 16917 67229
rect 16875 67180 16876 67220
rect 16916 67180 16917 67220
rect 16875 67171 16917 67180
rect 16683 67052 16725 67061
rect 16683 67012 16684 67052
rect 16724 67012 16725 67052
rect 16683 67003 16725 67012
rect 16876 66977 16916 67171
rect 16875 66968 16917 66977
rect 16875 66928 16876 66968
rect 16916 66928 16917 66968
rect 16875 66919 16917 66928
rect 16876 66834 16916 66919
rect 16587 66716 16629 66725
rect 16587 66676 16588 66716
rect 16628 66676 16629 66716
rect 16587 66667 16629 66676
rect 16588 65456 16628 66667
rect 16683 66128 16725 66137
rect 16972 66128 17012 67675
rect 17068 66884 17108 75571
rect 17259 74360 17301 74369
rect 17259 74320 17260 74360
rect 17300 74320 17301 74360
rect 17259 74311 17301 74320
rect 17163 74108 17205 74117
rect 17163 74068 17164 74108
rect 17204 74068 17205 74108
rect 17163 74059 17205 74068
rect 17164 73688 17204 74059
rect 17164 73639 17204 73648
rect 17163 73100 17205 73109
rect 17163 73060 17164 73100
rect 17204 73060 17205 73100
rect 17163 73051 17205 73060
rect 17164 73016 17204 73051
rect 17164 72428 17204 72976
rect 17260 72932 17300 74311
rect 17260 72857 17300 72892
rect 17259 72848 17301 72857
rect 17259 72808 17260 72848
rect 17300 72808 17301 72848
rect 17259 72799 17301 72808
rect 17164 72388 17289 72428
rect 17249 72227 17289 72388
rect 17249 72218 17300 72227
rect 17249 72178 17260 72218
rect 17249 72155 17300 72178
rect 17356 72218 17396 72227
rect 17259 72008 17301 72017
rect 17259 71968 17260 72008
rect 17300 71968 17301 72008
rect 17259 71959 17301 71968
rect 17164 71504 17204 71513
rect 17164 71345 17204 71464
rect 17163 71336 17205 71345
rect 17163 71296 17164 71336
rect 17204 71296 17205 71336
rect 17163 71287 17205 71296
rect 17164 70841 17204 71287
rect 17163 70832 17205 70841
rect 17163 70792 17164 70832
rect 17204 70792 17205 70832
rect 17163 70783 17205 70792
rect 17163 70580 17205 70589
rect 17163 70540 17164 70580
rect 17204 70540 17205 70580
rect 17163 70531 17205 70540
rect 17164 69987 17204 70531
rect 17164 69938 17204 69947
rect 17260 69833 17300 71959
rect 17356 71597 17396 72178
rect 17355 71588 17397 71597
rect 17355 71548 17356 71588
rect 17396 71548 17397 71588
rect 17355 71539 17397 71548
rect 17452 71513 17492 76579
rect 17548 76049 17588 76831
rect 17643 76208 17685 76217
rect 17643 76168 17644 76208
rect 17684 76168 17685 76208
rect 17643 76159 17685 76168
rect 17547 76040 17589 76049
rect 17547 76000 17548 76040
rect 17588 76000 17589 76040
rect 17547 75991 17589 76000
rect 17644 76040 17684 76159
rect 17644 75991 17684 76000
rect 17740 76040 17780 76049
rect 17547 75788 17589 75797
rect 17547 75748 17548 75788
rect 17588 75748 17589 75788
rect 17547 75739 17589 75748
rect 17548 74528 17588 75739
rect 17740 75629 17780 76000
rect 17739 75620 17781 75629
rect 17739 75580 17740 75620
rect 17780 75580 17781 75620
rect 17739 75571 17781 75580
rect 17548 74479 17588 74488
rect 17644 74528 17684 74537
rect 17451 71504 17493 71513
rect 17451 71464 17452 71504
rect 17492 71464 17493 71504
rect 17451 71455 17493 71464
rect 17356 71252 17396 71261
rect 17396 71212 17492 71252
rect 17356 71203 17396 71212
rect 17355 70832 17397 70841
rect 17355 70792 17356 70832
rect 17396 70792 17397 70832
rect 17355 70783 17397 70792
rect 17356 70673 17396 70783
rect 17355 70664 17397 70673
rect 17355 70624 17356 70664
rect 17396 70624 17397 70664
rect 17452 70664 17492 71212
rect 17644 70841 17684 74488
rect 17740 73016 17780 73025
rect 17740 71849 17780 72976
rect 17836 72344 17876 83476
rect 18316 83467 18356 83476
rect 18988 83516 19028 83525
rect 18988 83357 19028 83476
rect 18987 83348 19029 83357
rect 18987 83308 18988 83348
rect 19028 83308 19029 83348
rect 18987 83299 19029 83308
rect 18808 83180 19176 83189
rect 18848 83140 18890 83180
rect 18930 83140 18972 83180
rect 19012 83140 19054 83180
rect 19094 83140 19136 83180
rect 18808 83131 19176 83140
rect 19180 83012 19220 83021
rect 19276 83012 19316 83719
rect 19372 83644 19508 83684
rect 19372 83516 19412 83644
rect 19468 83600 19508 83644
rect 19468 83560 19796 83600
rect 19372 83467 19412 83476
rect 19659 83432 19701 83441
rect 19659 83392 19660 83432
rect 19700 83392 19701 83432
rect 19659 83383 19701 83392
rect 19467 83348 19509 83357
rect 19467 83308 19468 83348
rect 19508 83308 19509 83348
rect 19467 83299 19509 83308
rect 19220 82972 19316 83012
rect 19180 82963 19220 82972
rect 18987 82844 19029 82853
rect 18987 82804 18988 82844
rect 19028 82804 19029 82844
rect 18987 82795 19029 82804
rect 19372 82844 19412 82853
rect 18988 82710 19028 82795
rect 19372 81761 19412 82804
rect 19371 81752 19413 81761
rect 19371 81712 19372 81752
rect 19412 81712 19413 81752
rect 19371 81703 19413 81712
rect 18808 81668 19176 81677
rect 18848 81628 18890 81668
rect 18930 81628 18972 81668
rect 19012 81628 19054 81668
rect 19094 81628 19136 81668
rect 18808 81619 19176 81628
rect 19083 81500 19125 81509
rect 19083 81460 19084 81500
rect 19124 81460 19125 81500
rect 19083 81451 19125 81460
rect 18988 81332 19028 81341
rect 18988 81173 19028 81292
rect 18987 81164 19029 81173
rect 18987 81124 18988 81164
rect 19028 81124 19029 81164
rect 18987 81115 19029 81124
rect 18891 81080 18933 81089
rect 18891 81040 18892 81080
rect 18932 81040 18933 81080
rect 18891 81031 18933 81040
rect 18700 80492 18740 80501
rect 18508 80452 18700 80492
rect 18411 78308 18453 78317
rect 18411 78268 18412 78308
rect 18452 78268 18453 78308
rect 18411 78259 18453 78268
rect 18412 76712 18452 78259
rect 18508 77561 18548 80452
rect 18700 80443 18740 80452
rect 18892 80408 18932 81031
rect 18892 80359 18932 80368
rect 19084 80333 19124 81451
rect 19179 81416 19221 81425
rect 19179 81376 19180 81416
rect 19220 81376 19221 81416
rect 19179 81367 19221 81376
rect 19180 81282 19220 81367
rect 19371 81332 19413 81341
rect 19371 81292 19372 81332
rect 19412 81292 19413 81332
rect 19371 81283 19413 81292
rect 19372 81198 19412 81283
rect 19468 80912 19508 83299
rect 19564 83012 19604 83021
rect 19660 83012 19700 83383
rect 19604 82972 19700 83012
rect 19564 82963 19604 82972
rect 19659 82340 19701 82349
rect 19659 82300 19660 82340
rect 19700 82300 19701 82340
rect 19659 82291 19701 82300
rect 19563 81752 19605 81761
rect 19563 81712 19564 81752
rect 19604 81712 19605 81752
rect 19563 81703 19605 81712
rect 19564 81500 19604 81703
rect 19564 81451 19604 81460
rect 19660 81425 19700 82291
rect 19659 81416 19701 81425
rect 19659 81376 19660 81416
rect 19700 81376 19701 81416
rect 19659 81367 19701 81376
rect 19180 80872 19508 80912
rect 19180 80585 19220 80872
rect 19275 80744 19317 80753
rect 19275 80704 19276 80744
rect 19316 80704 19317 80744
rect 19275 80695 19317 80704
rect 19179 80576 19221 80585
rect 19179 80536 19180 80576
rect 19220 80536 19221 80576
rect 19179 80527 19221 80536
rect 19083 80324 19125 80333
rect 19083 80284 19084 80324
rect 19124 80284 19125 80324
rect 19083 80275 19125 80284
rect 18808 80156 19176 80165
rect 18848 80116 18890 80156
rect 18930 80116 18972 80156
rect 19012 80116 19054 80156
rect 19094 80116 19136 80156
rect 18808 80107 19176 80116
rect 19180 79988 19220 79997
rect 19276 79988 19316 80695
rect 19756 80660 19796 83560
rect 19660 80620 19796 80660
rect 19467 80576 19509 80585
rect 19467 80536 19468 80576
rect 19508 80536 19509 80576
rect 19467 80527 19509 80536
rect 19372 80492 19412 80501
rect 19372 80249 19412 80452
rect 19371 80240 19413 80249
rect 19371 80200 19372 80240
rect 19412 80200 19413 80240
rect 19371 80191 19413 80200
rect 19220 79948 19316 79988
rect 19371 79988 19413 79997
rect 19371 79948 19372 79988
rect 19412 79948 19413 79988
rect 19180 79939 19220 79948
rect 19371 79939 19413 79948
rect 18987 79820 19029 79829
rect 18987 79780 18988 79820
rect 19028 79780 19029 79820
rect 18987 79771 19029 79780
rect 19372 79820 19412 79939
rect 19372 79771 19412 79780
rect 18988 79686 19028 79771
rect 19275 79736 19317 79745
rect 19275 79696 19276 79736
rect 19316 79696 19317 79736
rect 19275 79687 19317 79696
rect 19179 79400 19221 79409
rect 19179 79360 19180 79400
rect 19220 79360 19221 79400
rect 19179 79351 19221 79360
rect 19180 79232 19220 79351
rect 19180 79183 19220 79192
rect 19276 79157 19316 79687
rect 19275 79148 19317 79157
rect 19275 79108 19276 79148
rect 19316 79108 19317 79148
rect 19275 79099 19317 79108
rect 18699 79064 18741 79073
rect 18699 79024 18700 79064
rect 18740 79024 18741 79064
rect 18699 79015 18741 79024
rect 18700 78476 18740 79015
rect 18988 78980 19028 78989
rect 19372 78980 19412 78989
rect 18988 78821 19028 78940
rect 19276 78940 19372 78980
rect 18987 78812 19029 78821
rect 18987 78772 18988 78812
rect 19028 78772 19029 78812
rect 18987 78763 19029 78772
rect 18808 78644 19176 78653
rect 18848 78604 18890 78644
rect 18930 78604 18972 78644
rect 19012 78604 19054 78644
rect 19094 78604 19136 78644
rect 18808 78595 19176 78604
rect 18796 78476 18836 78485
rect 18700 78436 18796 78476
rect 18796 78427 18836 78436
rect 19179 78476 19221 78485
rect 19179 78436 19180 78476
rect 19220 78436 19221 78476
rect 19179 78427 19221 78436
rect 19180 78342 19220 78427
rect 18604 78308 18644 78317
rect 18507 77552 18549 77561
rect 18507 77512 18508 77552
rect 18548 77512 18549 77552
rect 18507 77503 18549 77512
rect 18604 76964 18644 78268
rect 18987 78308 19029 78317
rect 18987 78268 18988 78308
rect 19028 78268 19029 78308
rect 18987 78259 19029 78268
rect 18988 78174 19028 78259
rect 19276 77645 19316 78940
rect 19372 78931 19412 78940
rect 19372 78308 19412 78317
rect 19372 78149 19412 78268
rect 19371 78140 19413 78149
rect 19371 78100 19372 78140
rect 19412 78100 19413 78140
rect 19371 78091 19413 78100
rect 19275 77636 19317 77645
rect 19275 77596 19276 77636
rect 19316 77596 19317 77636
rect 19275 77587 19317 77596
rect 18988 77552 19028 77563
rect 18988 77477 19028 77512
rect 19354 77481 19394 77490
rect 18987 77468 19029 77477
rect 18987 77428 18988 77468
rect 19028 77428 19029 77468
rect 18987 77419 19029 77428
rect 19084 77441 19354 77468
rect 19084 77428 19394 77441
rect 19084 77309 19124 77428
rect 19468 77384 19508 80527
rect 19564 80324 19604 80333
rect 19564 80081 19604 80284
rect 19563 80072 19605 80081
rect 19563 80032 19564 80072
rect 19604 80032 19605 80072
rect 19563 80023 19605 80032
rect 19660 79745 19700 80620
rect 19755 80492 19797 80501
rect 19755 80452 19756 80492
rect 19796 80452 19797 80492
rect 19755 80443 19797 80452
rect 19756 80358 19796 80443
rect 19756 79820 19796 79829
rect 19659 79736 19701 79745
rect 19659 79696 19660 79736
rect 19700 79696 19701 79736
rect 19659 79687 19701 79696
rect 19756 79577 19796 79780
rect 19564 79568 19604 79577
rect 19755 79568 19797 79577
rect 19604 79528 19700 79568
rect 19564 79519 19604 79528
rect 19563 78812 19605 78821
rect 19563 78772 19564 78812
rect 19604 78772 19605 78812
rect 19563 78763 19605 78772
rect 19564 78678 19604 78763
rect 19660 78737 19700 79528
rect 19755 79528 19756 79568
rect 19796 79528 19797 79568
rect 19755 79519 19797 79528
rect 19852 79400 19892 84727
rect 20523 84440 20565 84449
rect 20523 84400 20524 84440
rect 20564 84400 20565 84440
rect 20523 84391 20565 84400
rect 20048 83936 20416 83945
rect 20088 83896 20130 83936
rect 20170 83896 20212 83936
rect 20252 83896 20294 83936
rect 20334 83896 20376 83936
rect 20048 83887 20416 83896
rect 20048 82424 20416 82433
rect 20088 82384 20130 82424
rect 20170 82384 20212 82424
rect 20252 82384 20294 82424
rect 20334 82384 20376 82424
rect 20048 82375 20416 82384
rect 19947 81416 19989 81425
rect 19947 81376 19948 81416
rect 19988 81376 19989 81416
rect 19947 81367 19989 81376
rect 19948 80408 19988 81367
rect 20048 80912 20416 80921
rect 20088 80872 20130 80912
rect 20170 80872 20212 80912
rect 20252 80872 20294 80912
rect 20334 80872 20376 80912
rect 20048 80863 20416 80872
rect 19948 80359 19988 80368
rect 19947 79736 19989 79745
rect 19947 79696 19948 79736
rect 19988 79696 19989 79736
rect 19947 79687 19989 79696
rect 19948 79568 19988 79687
rect 19948 79519 19988 79528
rect 20048 79400 20416 79409
rect 19852 79360 19988 79400
rect 19851 79232 19893 79241
rect 19851 79192 19852 79232
rect 19892 79192 19893 79232
rect 19851 79183 19893 79192
rect 19756 78980 19796 78989
rect 19659 78728 19701 78737
rect 19659 78688 19660 78728
rect 19700 78688 19701 78728
rect 19659 78679 19701 78688
rect 19756 78476 19796 78940
rect 19660 78436 19796 78476
rect 19563 78392 19605 78401
rect 19563 78352 19564 78392
rect 19604 78352 19605 78392
rect 19563 78343 19605 78352
rect 19564 78258 19604 78343
rect 19660 77729 19700 78436
rect 19756 78308 19796 78317
rect 19852 78308 19892 79183
rect 19948 78980 19988 79360
rect 20088 79360 20130 79400
rect 20170 79360 20212 79400
rect 20252 79360 20294 79400
rect 20334 79360 20376 79400
rect 20048 79351 20416 79360
rect 19948 78940 20084 78980
rect 19948 78812 19988 78821
rect 19948 78569 19988 78772
rect 19947 78560 19989 78569
rect 19947 78520 19948 78560
rect 19988 78520 19989 78560
rect 19947 78511 19989 78520
rect 19796 78268 19892 78308
rect 19756 78259 19796 78268
rect 20044 78224 20084 78940
rect 19852 78184 20084 78224
rect 19659 77720 19701 77729
rect 19659 77680 19660 77720
rect 19700 77680 19701 77720
rect 19659 77671 19701 77680
rect 19852 77477 19892 78184
rect 19948 78056 19988 78065
rect 19756 77468 19796 77477
rect 19372 77344 19508 77384
rect 19660 77428 19756 77468
rect 19083 77300 19125 77309
rect 19083 77260 19084 77300
rect 19124 77260 19125 77300
rect 19083 77251 19125 77260
rect 19180 77300 19220 77309
rect 19220 77260 19316 77300
rect 19180 77251 19220 77260
rect 18808 77132 19176 77141
rect 18848 77092 18890 77132
rect 18930 77092 18972 77132
rect 19012 77092 19054 77132
rect 19094 77092 19136 77132
rect 18808 77083 19176 77092
rect 17932 76672 18412 76712
rect 17932 73109 17972 76672
rect 18412 76663 18452 76672
rect 18508 76924 18644 76964
rect 18123 76544 18165 76553
rect 18123 76504 18124 76544
rect 18164 76504 18165 76544
rect 18123 76495 18165 76504
rect 18124 75956 18164 76495
rect 18219 76040 18261 76049
rect 18219 76000 18220 76040
rect 18260 76000 18356 76040
rect 18219 75991 18261 76000
rect 18027 74612 18069 74621
rect 18027 74572 18028 74612
rect 18068 74572 18069 74612
rect 18027 74563 18069 74572
rect 18028 74528 18068 74563
rect 18028 74477 18068 74488
rect 18124 74444 18164 75916
rect 18220 75906 18260 75991
rect 18220 75293 18260 75337
rect 18219 75284 18261 75293
rect 18219 75244 18220 75284
rect 18260 75244 18261 75284
rect 18219 75242 18261 75244
rect 18219 75235 18220 75242
rect 18260 75235 18261 75242
rect 18220 75193 18260 75202
rect 18316 75116 18356 76000
rect 18508 75461 18548 76924
rect 18603 76796 18645 76805
rect 18603 76756 18604 76796
rect 18644 76756 18645 76796
rect 18603 76747 18645 76756
rect 18988 76796 19028 76805
rect 18604 76662 18644 76747
rect 18795 76712 18837 76721
rect 18795 76672 18796 76712
rect 18836 76672 18837 76712
rect 18795 76663 18837 76672
rect 18699 76628 18741 76637
rect 18699 76588 18700 76628
rect 18740 76588 18741 76628
rect 18699 76579 18741 76588
rect 18700 76040 18740 76579
rect 18796 76544 18836 76663
rect 18796 76495 18836 76504
rect 18988 76469 19028 76756
rect 19180 76544 19220 76553
rect 18987 76460 19029 76469
rect 18987 76420 18988 76460
rect 19028 76420 19029 76460
rect 18987 76411 19029 76420
rect 19180 76217 19220 76504
rect 19179 76208 19221 76217
rect 19179 76168 19180 76208
rect 19220 76168 19221 76208
rect 19179 76159 19221 76168
rect 19276 76040 19316 77260
rect 19372 76469 19412 77344
rect 19564 77300 19604 77309
rect 19468 77260 19564 77300
rect 19371 76460 19413 76469
rect 19371 76420 19372 76460
rect 19412 76420 19413 76460
rect 19371 76411 19413 76420
rect 19468 76385 19508 77260
rect 19564 77251 19604 77260
rect 19564 76796 19604 76805
rect 19467 76376 19509 76385
rect 19467 76336 19468 76376
rect 19508 76336 19509 76376
rect 19467 76327 19509 76336
rect 19371 76124 19413 76133
rect 19564 76124 19604 76756
rect 19660 76133 19700 77428
rect 19756 77419 19796 77428
rect 19851 77468 19893 77477
rect 19851 77428 19852 77468
rect 19892 77428 19893 77468
rect 19948 77468 19988 78016
rect 20048 77888 20416 77897
rect 20088 77848 20130 77888
rect 20170 77848 20212 77888
rect 20252 77848 20294 77888
rect 20334 77848 20376 77888
rect 20048 77839 20416 77848
rect 19948 77428 20084 77468
rect 19851 77419 19893 77428
rect 19948 77300 19988 77309
rect 19852 77260 19948 77300
rect 19852 76805 19892 77260
rect 19948 77251 19988 77260
rect 20044 77057 20084 77428
rect 20043 77048 20085 77057
rect 20043 77008 20044 77048
rect 20084 77008 20085 77048
rect 20043 76999 20085 77008
rect 19851 76796 19893 76805
rect 19851 76756 19852 76796
rect 19892 76756 19893 76796
rect 19851 76747 19893 76756
rect 19948 76796 19988 76805
rect 19948 76553 19988 76756
rect 20140 76553 20180 76638
rect 19756 76544 19796 76553
rect 19947 76544 19989 76553
rect 19796 76504 19892 76544
rect 19756 76495 19796 76504
rect 19755 76292 19797 76301
rect 19755 76252 19756 76292
rect 19796 76252 19797 76292
rect 19755 76243 19797 76252
rect 19371 76084 19372 76124
rect 19412 76084 19413 76124
rect 19371 76075 19413 76084
rect 19468 76084 19604 76124
rect 19659 76124 19701 76133
rect 19659 76084 19660 76124
rect 19700 76084 19701 76124
rect 18700 75991 18740 76000
rect 19228 76030 19316 76040
rect 19268 76000 19316 76030
rect 19372 75990 19412 76075
rect 19228 75981 19268 75990
rect 18808 75620 19176 75629
rect 18848 75580 18890 75620
rect 18930 75580 18972 75620
rect 19012 75580 19054 75620
rect 19094 75580 19136 75620
rect 18808 75571 19176 75580
rect 18507 75452 18549 75461
rect 18507 75412 18508 75452
rect 18548 75412 18549 75452
rect 18507 75403 18549 75412
rect 18796 75293 18836 75324
rect 18795 75284 18837 75293
rect 18795 75244 18796 75284
rect 18836 75244 18837 75284
rect 18795 75235 18837 75244
rect 18796 75200 18836 75235
rect 18796 75116 18836 75160
rect 18124 73277 18164 74404
rect 18220 75076 18356 75116
rect 18700 75076 18836 75116
rect 18123 73268 18165 73277
rect 18123 73228 18124 73268
rect 18164 73228 18165 73268
rect 18123 73219 18165 73228
rect 17931 73100 17973 73109
rect 18220 73100 18260 75076
rect 18412 75032 18452 75041
rect 17931 73060 17932 73100
rect 17972 73060 17973 73100
rect 17931 73051 17973 73060
rect 18172 73060 18260 73100
rect 18316 74992 18412 75032
rect 18172 73016 18212 73060
rect 18316 73016 18356 74992
rect 18412 74983 18452 74992
rect 18603 75032 18645 75041
rect 18603 74992 18604 75032
rect 18644 74992 18645 75032
rect 18603 74983 18645 74992
rect 18604 74898 18644 74983
rect 18603 74780 18645 74789
rect 18603 74740 18604 74780
rect 18644 74740 18645 74780
rect 18603 74731 18645 74740
rect 18604 74528 18644 74731
rect 18412 73688 18452 73699
rect 18604 73697 18644 74488
rect 18412 73613 18452 73648
rect 18603 73688 18645 73697
rect 18603 73648 18604 73688
rect 18644 73648 18645 73688
rect 18603 73639 18645 73648
rect 18700 73613 18740 75076
rect 19083 75032 19125 75041
rect 19083 74992 19084 75032
rect 19124 74992 19125 75032
rect 19083 74983 19125 74992
rect 19084 74523 19124 74983
rect 19468 74780 19508 76084
rect 19659 76075 19701 76084
rect 19564 75956 19604 75965
rect 19756 75956 19796 76243
rect 19564 75881 19604 75916
rect 19553 75872 19604 75881
rect 19553 75832 19554 75872
rect 19594 75832 19604 75872
rect 19660 75916 19796 75956
rect 19553 75823 19595 75832
rect 19563 75704 19605 75713
rect 19563 75664 19564 75704
rect 19604 75664 19605 75704
rect 19563 75655 19605 75664
rect 19084 74474 19124 74483
rect 19180 74740 19508 74780
rect 19180 74276 19220 74740
rect 19276 74612 19316 74621
rect 19276 74444 19316 74572
rect 19450 74457 19490 74466
rect 19276 74417 19450 74444
rect 19276 74404 19490 74417
rect 19564 74360 19604 75655
rect 19660 74948 19700 75916
rect 19755 75788 19797 75797
rect 19755 75748 19756 75788
rect 19796 75748 19797 75788
rect 19755 75739 19797 75748
rect 19756 75654 19796 75739
rect 19852 75125 19892 76504
rect 19947 76504 19948 76544
rect 19988 76504 19989 76544
rect 19947 76495 19989 76504
rect 20139 76544 20181 76553
rect 20139 76504 20140 76544
rect 20180 76504 20181 76544
rect 20139 76495 20181 76504
rect 19947 76376 19989 76385
rect 19947 76336 19948 76376
rect 19988 76336 19989 76376
rect 19947 76327 19989 76336
rect 20048 76376 20416 76385
rect 20088 76336 20130 76376
rect 20170 76336 20212 76376
rect 20252 76336 20294 76376
rect 20334 76336 20376 76376
rect 20048 76327 20416 76336
rect 19948 76124 19988 76327
rect 19948 76084 20084 76124
rect 19947 75956 19989 75965
rect 19947 75916 19948 75956
rect 19988 75916 19989 75956
rect 19947 75907 19989 75916
rect 19948 75822 19988 75907
rect 20044 75713 20084 76084
rect 20140 75788 20180 75797
rect 20043 75704 20085 75713
rect 20043 75664 20044 75704
rect 20084 75664 20085 75704
rect 20043 75655 20085 75664
rect 20043 75536 20085 75545
rect 20043 75496 20044 75536
rect 20084 75496 20085 75536
rect 20043 75487 20085 75496
rect 20044 75200 20084 75487
rect 20044 75151 20084 75160
rect 19851 75116 19893 75125
rect 19851 75076 19852 75116
rect 19892 75076 19893 75116
rect 19851 75067 19893 75076
rect 20140 75041 20180 75748
rect 20139 75032 20181 75041
rect 20139 74992 20140 75032
rect 20180 74992 20181 75032
rect 20139 74983 20181 74992
rect 19660 74908 19988 74948
rect 19852 74453 19892 74538
rect 19851 74444 19893 74453
rect 19851 74404 19852 74444
rect 19892 74404 19893 74444
rect 19851 74395 19893 74404
rect 19372 74320 19604 74360
rect 19180 74236 19316 74276
rect 19276 74117 19316 74236
rect 18808 74108 19176 74117
rect 18848 74068 18890 74108
rect 18930 74068 18972 74108
rect 19012 74068 19054 74108
rect 19094 74068 19136 74108
rect 18808 74059 19176 74068
rect 19275 74108 19317 74117
rect 19275 74068 19276 74108
rect 19316 74068 19317 74108
rect 19275 74059 19317 74068
rect 18891 73940 18933 73949
rect 19372 73940 19412 74320
rect 19660 74276 19700 74285
rect 18891 73900 18892 73940
rect 18932 73900 18933 73940
rect 18891 73891 18933 73900
rect 19276 73900 19412 73940
rect 19468 74236 19660 74276
rect 18411 73604 18453 73613
rect 18411 73564 18412 73604
rect 18452 73564 18453 73604
rect 18411 73555 18453 73564
rect 18699 73604 18741 73613
rect 18699 73564 18700 73604
rect 18740 73564 18741 73604
rect 18699 73555 18741 73564
rect 18604 73520 18644 73529
rect 18412 73184 18452 73193
rect 18412 73025 18452 73144
rect 18604 73100 18644 73480
rect 18892 73100 18932 73891
rect 18988 73772 19028 73781
rect 18988 73109 19028 73732
rect 19179 73688 19221 73697
rect 19179 73648 19180 73688
rect 19220 73648 19221 73688
rect 19179 73639 19221 73648
rect 19180 73520 19220 73639
rect 19180 73471 19220 73480
rect 18508 73060 18644 73100
rect 18700 73060 18932 73100
rect 18987 73100 19029 73109
rect 18987 73060 18988 73100
rect 19028 73060 19029 73100
rect 18028 72976 18212 73016
rect 18268 73006 18356 73016
rect 17836 72304 17972 72344
rect 17836 72176 17876 72187
rect 17836 72101 17876 72136
rect 17835 72092 17877 72101
rect 17835 72052 17836 72092
rect 17876 72052 17877 72092
rect 17835 72043 17877 72052
rect 17739 71840 17781 71849
rect 17739 71800 17740 71840
rect 17780 71800 17781 71840
rect 17739 71791 17781 71800
rect 17740 71504 17780 71513
rect 17740 71009 17780 71464
rect 17739 71000 17781 71009
rect 17739 70960 17740 71000
rect 17780 70960 17781 71000
rect 17739 70951 17781 70960
rect 17643 70832 17685 70841
rect 17932 70832 17972 72304
rect 17643 70792 17644 70832
rect 17684 70792 17685 70832
rect 17643 70783 17685 70792
rect 17836 70792 17972 70832
rect 17452 70624 17684 70664
rect 17355 70615 17397 70624
rect 17356 70530 17396 70615
rect 17548 70496 17588 70505
rect 17355 70244 17397 70253
rect 17355 70204 17356 70244
rect 17396 70204 17397 70244
rect 17355 70195 17397 70204
rect 17356 70160 17396 70195
rect 17356 70109 17396 70120
rect 17259 69824 17301 69833
rect 17259 69784 17260 69824
rect 17300 69784 17301 69824
rect 17259 69775 17301 69784
rect 17548 69320 17588 70456
rect 17644 69992 17684 70624
rect 17739 70580 17781 70589
rect 17739 70540 17740 70580
rect 17780 70540 17781 70580
rect 17739 70531 17781 70540
rect 17740 70446 17780 70531
rect 17644 69943 17684 69952
rect 17739 69992 17781 70001
rect 17739 69952 17740 69992
rect 17780 69952 17781 69992
rect 17739 69943 17781 69952
rect 17740 69858 17780 69943
rect 17836 69329 17876 70792
rect 17931 70664 17973 70673
rect 17931 70624 17932 70664
rect 17972 70624 17973 70664
rect 17931 70615 17973 70624
rect 17932 70530 17972 70615
rect 17931 69992 17973 70001
rect 17931 69952 17932 69992
rect 17972 69952 17973 69992
rect 17931 69943 17973 69952
rect 17835 69320 17877 69329
rect 17548 69280 17684 69320
rect 17356 69152 17396 69161
rect 17356 68993 17396 69112
rect 17355 68984 17397 68993
rect 17355 68944 17356 68984
rect 17396 68944 17397 68984
rect 17355 68935 17397 68944
rect 17548 68984 17588 68993
rect 17548 68312 17588 68944
rect 17644 68480 17684 69280
rect 17835 69280 17836 69320
rect 17876 69280 17877 69320
rect 17835 69271 17877 69280
rect 17932 69320 17972 69943
rect 17932 69271 17972 69280
rect 17739 69236 17781 69245
rect 17739 69196 17740 69236
rect 17780 69196 17781 69236
rect 17739 69187 17781 69196
rect 17740 69102 17780 69187
rect 17739 68984 17781 68993
rect 17739 68944 17740 68984
rect 17780 68944 17781 68984
rect 17739 68935 17781 68944
rect 17740 68489 17780 68935
rect 17644 68431 17684 68440
rect 17739 68480 17781 68489
rect 17931 68480 17973 68489
rect 17739 68440 17740 68480
rect 17780 68440 17781 68480
rect 17739 68431 17781 68440
rect 17836 68440 17932 68480
rect 17972 68440 17973 68480
rect 17548 68272 17780 68312
rect 17164 68228 17204 68237
rect 17204 68188 17396 68228
rect 17164 68179 17204 68188
rect 17259 67976 17301 67985
rect 17259 67936 17260 67976
rect 17300 67936 17301 67976
rect 17259 67927 17301 67936
rect 17260 67733 17300 67927
rect 17259 67724 17301 67733
rect 17259 67684 17260 67724
rect 17300 67684 17301 67724
rect 17259 67675 17301 67684
rect 17260 67640 17300 67675
rect 17260 67589 17300 67600
rect 17259 67388 17301 67397
rect 17259 67348 17260 67388
rect 17300 67348 17301 67388
rect 17259 67339 17301 67348
rect 17260 66968 17300 67339
rect 17356 67136 17396 68188
rect 17643 68144 17685 68153
rect 17643 68104 17644 68144
rect 17684 68104 17685 68144
rect 17643 68095 17685 68104
rect 17547 67640 17589 67649
rect 17547 67600 17548 67640
rect 17588 67600 17589 67640
rect 17547 67591 17589 67600
rect 17356 67096 17492 67136
rect 17260 66919 17300 66928
rect 17068 66844 17204 66884
rect 17067 66716 17109 66725
rect 17067 66676 17068 66716
rect 17108 66676 17109 66716
rect 17067 66667 17109 66676
rect 17068 66582 17108 66667
rect 17164 66296 17204 66844
rect 17204 66256 17396 66296
rect 17164 66247 17204 66256
rect 17356 66137 17396 66256
rect 17355 66128 17397 66137
rect 16683 66088 16684 66128
rect 16724 66088 16725 66128
rect 16683 66079 16725 66088
rect 16780 66088 17204 66128
rect 16684 65633 16724 66079
rect 16683 65624 16725 65633
rect 16683 65584 16684 65624
rect 16724 65584 16725 65624
rect 16683 65575 16725 65584
rect 16588 65407 16628 65416
rect 16684 65456 16724 65575
rect 16684 64625 16724 65416
rect 16683 64616 16725 64625
rect 16683 64576 16684 64616
rect 16724 64576 16725 64616
rect 16683 64567 16725 64576
rect 16780 64280 16820 66088
rect 16875 65960 16917 65969
rect 16875 65920 16876 65960
rect 16916 65920 16917 65960
rect 16875 65911 16917 65920
rect 16684 64240 16820 64280
rect 16491 62600 16533 62609
rect 16491 62560 16492 62600
rect 16532 62560 16533 62600
rect 16491 62551 16533 62560
rect 16588 62348 16628 62357
rect 16588 61349 16628 62308
rect 16684 61760 16724 64240
rect 16780 63104 16820 63115
rect 16780 63029 16820 63064
rect 16779 63020 16821 63029
rect 16779 62980 16780 63020
rect 16820 62980 16821 63020
rect 16779 62971 16821 62980
rect 16779 62600 16821 62609
rect 16779 62560 16780 62600
rect 16820 62560 16821 62600
rect 16779 62551 16821 62560
rect 16780 62466 16820 62551
rect 16684 61720 16820 61760
rect 16587 61340 16629 61349
rect 16587 61300 16588 61340
rect 16628 61300 16629 61340
rect 16587 61291 16629 61300
rect 16588 60836 16628 60847
rect 16588 60761 16628 60796
rect 16684 60836 16724 60845
rect 16587 60752 16629 60761
rect 16587 60712 16588 60752
rect 16628 60712 16629 60752
rect 16587 60703 16629 60712
rect 16684 60593 16724 60796
rect 16683 60584 16725 60593
rect 16683 60544 16684 60584
rect 16724 60544 16725 60584
rect 16683 60535 16725 60544
rect 16587 60080 16629 60089
rect 16587 60040 16588 60080
rect 16628 60040 16629 60080
rect 16587 60031 16629 60040
rect 16395 56636 16437 56645
rect 16395 56596 16396 56636
rect 16436 56596 16437 56636
rect 16395 56587 16437 56596
rect 16491 56300 16533 56309
rect 16491 56260 16492 56300
rect 16532 56260 16533 56300
rect 16491 56251 16533 56260
rect 16492 56166 16532 56251
rect 16491 55796 16533 55805
rect 16491 55756 16492 55796
rect 16532 55756 16533 55796
rect 16491 55747 16533 55756
rect 16299 55040 16341 55049
rect 16299 55000 16300 55040
rect 16340 55000 16341 55040
rect 16299 54991 16341 55000
rect 16300 54906 16340 54991
rect 16204 54160 16340 54200
rect 16204 54037 16244 54046
rect 16204 53873 16244 53997
rect 16203 53864 16245 53873
rect 16203 53824 16204 53864
rect 16244 53824 16245 53864
rect 16203 53815 16245 53824
rect 16107 53612 16149 53621
rect 16107 53572 16108 53612
rect 16148 53572 16149 53612
rect 16107 53563 16149 53572
rect 16107 52856 16149 52865
rect 16107 52816 16108 52856
rect 16148 52816 16149 52856
rect 16107 52807 16149 52816
rect 16108 52772 16148 52807
rect 16108 52721 16148 52732
rect 15916 52648 16052 52688
rect 15916 52520 15956 52529
rect 15916 52109 15956 52480
rect 15915 52100 15957 52109
rect 15915 52060 15916 52100
rect 15956 52060 15957 52100
rect 15915 52051 15957 52060
rect 15820 51967 15860 51976
rect 15915 51932 15957 51941
rect 15915 51892 15916 51932
rect 15956 51892 15957 51932
rect 15915 51883 15957 51892
rect 15916 51848 15956 51883
rect 15916 51797 15956 51808
rect 15723 50672 15765 50681
rect 15723 50632 15724 50672
rect 15764 50632 15765 50672
rect 15723 50623 15765 50632
rect 15531 50464 15532 50504
rect 15572 50464 15668 50504
rect 15723 50504 15765 50513
rect 15723 50464 15724 50504
rect 15764 50464 15765 50504
rect 15531 50455 15573 50464
rect 15723 50455 15765 50464
rect 15435 50420 15477 50429
rect 15435 50380 15436 50420
rect 15476 50380 15477 50420
rect 15435 50371 15477 50380
rect 15436 49496 15476 50371
rect 15532 50336 15572 50345
rect 15532 50177 15572 50296
rect 15627 50336 15669 50345
rect 15627 50296 15628 50336
rect 15668 50296 15669 50336
rect 15627 50287 15669 50296
rect 15531 50168 15573 50177
rect 15531 50128 15532 50168
rect 15572 50128 15573 50168
rect 15531 50119 15573 50128
rect 15339 49244 15381 49253
rect 15339 49204 15340 49244
rect 15380 49204 15381 49244
rect 15339 49195 15381 49204
rect 15052 49036 15188 49076
rect 14956 48824 14996 48833
rect 14956 48749 14996 48784
rect 14955 48740 14997 48749
rect 14955 48700 14956 48740
rect 14996 48700 14997 48740
rect 15052 48740 15092 49036
rect 15148 48908 15188 48917
rect 15436 48908 15476 49456
rect 15532 49496 15572 49505
rect 15532 49169 15572 49456
rect 15628 49496 15668 50287
rect 15628 49447 15668 49456
rect 15724 49496 15764 50455
rect 16012 49664 16052 52648
rect 16300 52109 16340 54160
rect 16395 53696 16437 53705
rect 16395 53656 16396 53696
rect 16436 53656 16437 53696
rect 16395 53647 16437 53656
rect 16396 52184 16436 53647
rect 16492 52697 16532 55747
rect 16588 55460 16628 60031
rect 16684 59324 16724 59333
rect 16684 56981 16724 59284
rect 16780 58736 16820 61720
rect 16876 60005 16916 65911
rect 17067 65456 17109 65465
rect 17067 65416 17068 65456
rect 17108 65416 17109 65456
rect 17067 65407 17109 65416
rect 17164 65456 17204 66088
rect 17355 66088 17356 66128
rect 17396 66088 17397 66128
rect 17355 66079 17397 66088
rect 17452 66128 17492 67096
rect 17548 66296 17588 67591
rect 17644 67556 17684 68095
rect 17740 67654 17780 68272
rect 17740 67605 17780 67614
rect 17644 67516 17780 67556
rect 17548 66256 17684 66296
rect 17452 66079 17492 66088
rect 17547 66128 17589 66137
rect 17547 66088 17548 66128
rect 17588 66088 17589 66128
rect 17547 66079 17589 66088
rect 17548 65994 17588 66079
rect 17644 65876 17684 66256
rect 17164 65407 17204 65416
rect 17548 65836 17684 65876
rect 17068 65322 17108 65407
rect 16972 64616 17012 64656
rect 16972 64541 17012 64576
rect 17067 64616 17109 64625
rect 17067 64576 17068 64616
rect 17108 64576 17109 64616
rect 17067 64567 17109 64576
rect 16971 64532 17013 64541
rect 16971 64492 16972 64532
rect 17012 64492 17013 64532
rect 16971 64483 17013 64492
rect 16972 63197 17012 64483
rect 17068 63272 17108 64567
rect 17164 64448 17204 64457
rect 17204 64408 17492 64448
rect 17164 64399 17204 64408
rect 17452 63944 17492 64408
rect 17452 63895 17492 63904
rect 17548 63944 17588 65836
rect 17740 65792 17780 67516
rect 17739 65752 17780 65792
rect 17836 65792 17876 68440
rect 17931 68431 17973 68440
rect 17931 67976 17973 67985
rect 17931 67936 17932 67976
rect 17972 67936 17973 67976
rect 17931 67927 17973 67936
rect 17932 67556 17972 67927
rect 17932 67507 17972 67516
rect 18028 66212 18068 72976
rect 18308 72976 18356 73006
rect 18411 73016 18453 73025
rect 18411 72976 18412 73016
rect 18452 72976 18453 73016
rect 18411 72967 18453 72976
rect 18268 72957 18308 72966
rect 18412 72965 18452 72967
rect 18123 72848 18165 72857
rect 18123 72808 18124 72848
rect 18164 72808 18260 72848
rect 18123 72799 18165 72808
rect 18124 70085 18164 70087
rect 18123 70076 18165 70085
rect 18123 70036 18124 70076
rect 18164 70036 18165 70076
rect 18220 70076 18260 72808
rect 18364 72185 18404 72194
rect 18508 72176 18548 73060
rect 18604 72932 18644 72941
rect 18604 72605 18644 72892
rect 18603 72596 18645 72605
rect 18603 72556 18604 72596
rect 18644 72556 18645 72596
rect 18603 72547 18645 72556
rect 18404 72145 18548 72176
rect 18364 72136 18548 72145
rect 18411 72008 18453 72017
rect 18411 71968 18412 72008
rect 18452 71968 18453 72008
rect 18411 71959 18453 71968
rect 18508 72008 18548 72017
rect 18700 72008 18740 73060
rect 18987 73051 19029 73060
rect 18796 72857 18836 72942
rect 18987 72932 19029 72941
rect 18987 72892 18988 72932
rect 19028 72892 19029 72932
rect 18987 72883 19029 72892
rect 18795 72848 18837 72857
rect 18795 72808 18796 72848
rect 18836 72808 18837 72848
rect 18795 72799 18837 72808
rect 18988 72798 19028 72883
rect 19180 72857 19220 72942
rect 19179 72848 19221 72857
rect 19179 72808 19180 72848
rect 19220 72808 19221 72848
rect 19179 72799 19221 72808
rect 18808 72596 19176 72605
rect 18848 72556 18890 72596
rect 18930 72556 18972 72596
rect 19012 72556 19054 72596
rect 19094 72556 19136 72596
rect 18808 72547 19176 72556
rect 18795 72428 18837 72437
rect 18795 72388 18796 72428
rect 18836 72388 18837 72428
rect 18795 72379 18837 72388
rect 18987 72428 19029 72437
rect 18987 72388 18988 72428
rect 19028 72388 19029 72428
rect 18987 72379 19029 72388
rect 19180 72428 19220 72437
rect 19276 72428 19316 73900
rect 19372 73772 19412 73781
rect 19372 73193 19412 73732
rect 19371 73184 19413 73193
rect 19371 73144 19372 73184
rect 19412 73144 19413 73184
rect 19371 73135 19413 73144
rect 19220 72388 19316 72428
rect 19372 72932 19412 72941
rect 19372 72428 19412 72892
rect 19468 72689 19508 74236
rect 19660 74227 19700 74236
rect 19755 74276 19797 74285
rect 19755 74236 19756 74276
rect 19796 74236 19797 74276
rect 19755 74227 19797 74236
rect 19756 73940 19796 74227
rect 19948 74108 19988 74908
rect 20048 74864 20416 74873
rect 20088 74824 20130 74864
rect 20170 74824 20212 74864
rect 20252 74824 20294 74864
rect 20334 74824 20376 74864
rect 20048 74815 20416 74824
rect 20044 74285 20084 74370
rect 20043 74276 20085 74285
rect 20043 74236 20044 74276
rect 20084 74236 20085 74276
rect 20043 74227 20085 74236
rect 19948 74068 20084 74108
rect 19660 73900 19796 73940
rect 19947 73940 19989 73949
rect 19947 73900 19948 73940
rect 19988 73900 19989 73940
rect 19564 73520 19604 73529
rect 19564 73025 19604 73480
rect 19563 73016 19605 73025
rect 19563 72976 19564 73016
rect 19604 72976 19605 73016
rect 19563 72967 19605 72976
rect 19564 72764 19604 72773
rect 19467 72680 19509 72689
rect 19467 72640 19468 72680
rect 19508 72640 19509 72680
rect 19467 72631 19509 72640
rect 19372 72388 19508 72428
rect 19180 72379 19220 72388
rect 18548 71968 18740 72008
rect 18508 71959 18548 71968
rect 18220 70036 18356 70076
rect 18123 70027 18165 70036
rect 18124 69992 18164 70027
rect 18124 69943 18164 69952
rect 18220 69908 18260 69919
rect 18220 69833 18260 69868
rect 18219 69824 18261 69833
rect 18219 69784 18220 69824
rect 18260 69784 18261 69824
rect 18219 69775 18261 69784
rect 18123 69740 18165 69749
rect 18123 69700 18124 69740
rect 18164 69700 18165 69740
rect 18123 69691 18165 69700
rect 18124 69152 18164 69691
rect 18124 68657 18164 69112
rect 18123 68648 18165 68657
rect 18123 68608 18124 68648
rect 18164 68608 18165 68648
rect 18123 68599 18165 68608
rect 18220 68480 18260 68489
rect 18316 68480 18356 70036
rect 18412 68489 18452 71959
rect 18507 71840 18549 71849
rect 18507 71800 18508 71840
rect 18548 71800 18549 71840
rect 18507 71791 18549 71800
rect 18260 68440 18356 68480
rect 18220 68431 18260 68440
rect 18124 68396 18164 68405
rect 18124 68069 18164 68356
rect 18123 68060 18165 68069
rect 18123 68020 18124 68060
rect 18164 68020 18165 68060
rect 18123 68011 18165 68020
rect 17931 66128 17973 66137
rect 17931 66088 17932 66128
rect 17972 66088 17973 66128
rect 17931 66079 17973 66088
rect 17932 65994 17972 66079
rect 17836 65752 17972 65792
rect 17739 65708 17779 65752
rect 17739 65668 17876 65708
rect 17643 65624 17685 65633
rect 17643 65584 17644 65624
rect 17684 65584 17685 65624
rect 17643 65575 17685 65584
rect 17164 63272 17204 63281
rect 17068 63232 17164 63272
rect 17164 63223 17204 63232
rect 17259 63272 17301 63281
rect 17548 63272 17588 63904
rect 17644 65456 17684 65575
rect 17739 65540 17781 65549
rect 17739 65500 17740 65540
rect 17780 65500 17781 65540
rect 17739 65491 17781 65500
rect 17644 63281 17684 65416
rect 17740 64709 17780 65491
rect 17739 64700 17781 64709
rect 17739 64660 17740 64700
rect 17780 64660 17781 64700
rect 17739 64651 17781 64660
rect 17740 64616 17780 64651
rect 17740 64565 17780 64576
rect 17836 64280 17876 65668
rect 17932 65633 17972 65752
rect 17931 65624 17973 65633
rect 17931 65584 17932 65624
rect 17972 65584 17973 65624
rect 17931 65575 17973 65584
rect 18028 65288 18068 66172
rect 18124 67640 18164 67649
rect 18124 65717 18164 67600
rect 18316 67388 18356 68440
rect 18411 68480 18453 68489
rect 18411 68440 18412 68480
rect 18452 68440 18453 68480
rect 18411 68431 18453 68440
rect 18508 67733 18548 71791
rect 18796 71252 18836 72379
rect 18988 72260 19028 72379
rect 18988 72211 19028 72220
rect 19371 72260 19413 72269
rect 19371 72220 19372 72260
rect 19412 72220 19413 72260
rect 19371 72211 19413 72220
rect 19372 72126 19412 72211
rect 18891 71756 18933 71765
rect 18891 71716 18892 71756
rect 18932 71716 18933 71756
rect 18891 71707 18933 71716
rect 18892 71261 18932 71707
rect 19468 71681 19508 72388
rect 19564 72176 19604 72724
rect 19660 72353 19700 73900
rect 19947 73891 19989 73900
rect 19948 73806 19988 73891
rect 19755 73772 19797 73781
rect 19755 73732 19756 73772
rect 19796 73732 19797 73772
rect 19755 73723 19797 73732
rect 19756 73638 19796 73723
rect 20044 73520 20084 74068
rect 19948 73480 20084 73520
rect 19948 73100 19988 73480
rect 20048 73352 20416 73361
rect 20088 73312 20130 73352
rect 20170 73312 20212 73352
rect 20252 73312 20294 73352
rect 20334 73312 20376 73352
rect 20048 73303 20416 73312
rect 19852 73060 19988 73100
rect 19756 72932 19796 72941
rect 19756 72773 19796 72892
rect 19755 72764 19797 72773
rect 19755 72724 19756 72764
rect 19796 72724 19797 72764
rect 19755 72715 19797 72724
rect 19659 72344 19701 72353
rect 19659 72304 19660 72344
rect 19700 72304 19701 72344
rect 19659 72295 19701 72304
rect 19755 72260 19797 72269
rect 19755 72220 19756 72260
rect 19796 72220 19797 72260
rect 19755 72211 19797 72220
rect 19564 72136 19700 72176
rect 19563 72008 19605 72017
rect 19563 71968 19564 72008
rect 19604 71968 19605 72008
rect 19563 71959 19605 71968
rect 19564 71874 19604 71959
rect 19467 71672 19509 71681
rect 19467 71632 19468 71672
rect 19508 71632 19509 71672
rect 19467 71623 19509 71632
rect 18988 71504 19028 71513
rect 18988 71345 19028 71464
rect 19372 71420 19412 71429
rect 19412 71380 19508 71420
rect 19372 71371 19412 71380
rect 18987 71336 19029 71345
rect 18987 71296 18988 71336
rect 19028 71296 19029 71336
rect 18987 71287 19029 71296
rect 18700 71212 18836 71252
rect 18891 71252 18933 71261
rect 18891 71212 18892 71252
rect 18932 71212 18933 71252
rect 18700 69992 18740 71212
rect 18891 71203 18933 71212
rect 19180 71252 19220 71261
rect 19371 71252 19413 71261
rect 19220 71212 19316 71252
rect 19180 71203 19220 71212
rect 18808 71084 19176 71093
rect 18848 71044 18890 71084
rect 18930 71044 18972 71084
rect 19012 71044 19054 71084
rect 19094 71044 19136 71084
rect 18808 71035 19176 71044
rect 19179 70916 19221 70925
rect 19179 70876 19180 70916
rect 19220 70876 19221 70916
rect 19179 70867 19221 70876
rect 19180 70664 19220 70867
rect 19180 70615 19220 70624
rect 19276 69992 19316 71212
rect 19371 71212 19372 71252
rect 19412 71212 19413 71252
rect 19371 71203 19413 71212
rect 19372 70748 19412 71203
rect 19372 70699 19412 70708
rect 19468 70580 19508 71380
rect 19660 71345 19700 72136
rect 19756 72126 19796 72211
rect 19659 71336 19701 71345
rect 19659 71296 19660 71336
rect 19700 71296 19701 71336
rect 19659 71287 19701 71296
rect 19564 71252 19604 71261
rect 19564 70664 19604 71212
rect 19755 70748 19797 70757
rect 19755 70708 19756 70748
rect 19796 70708 19797 70748
rect 19755 70699 19797 70708
rect 19564 70624 19700 70664
rect 19372 70540 19508 70580
rect 19372 70253 19412 70540
rect 19564 70496 19604 70505
rect 19468 70456 19564 70496
rect 19371 70244 19413 70253
rect 19371 70204 19372 70244
rect 19412 70204 19413 70244
rect 19371 70195 19413 70204
rect 18700 69077 18740 69952
rect 19228 69982 19316 69992
rect 19268 69952 19316 69982
rect 19372 70076 19412 70085
rect 19228 69933 19268 69942
rect 18808 69572 19176 69581
rect 18848 69532 18890 69572
rect 18930 69532 18972 69572
rect 19012 69532 19054 69572
rect 19094 69532 19136 69572
rect 18808 69523 19176 69532
rect 19372 69329 19412 70036
rect 19468 69413 19508 70456
rect 19564 70447 19604 70456
rect 19660 70085 19700 70624
rect 19756 70614 19796 70699
rect 19659 70076 19701 70085
rect 19659 70036 19660 70076
rect 19700 70036 19701 70076
rect 19659 70027 19701 70036
rect 19564 69908 19604 69917
rect 19604 69868 19700 69908
rect 19564 69859 19604 69868
rect 19467 69404 19509 69413
rect 19467 69364 19468 69404
rect 19508 69364 19509 69404
rect 19467 69355 19509 69364
rect 19371 69320 19413 69329
rect 19371 69280 19372 69320
rect 19412 69280 19413 69320
rect 19371 69271 19413 69280
rect 18891 69152 18933 69161
rect 18891 69112 18892 69152
rect 18932 69112 18933 69152
rect 18891 69103 18933 69112
rect 19372 69152 19412 69161
rect 18699 69068 18741 69077
rect 18699 69028 18700 69068
rect 18740 69028 18741 69068
rect 18699 69019 18741 69028
rect 18700 68489 18740 68574
rect 18892 68573 18932 69103
rect 19372 69068 19412 69112
rect 19084 69028 19412 69068
rect 18891 68564 18933 68573
rect 18891 68524 18892 68564
rect 18932 68524 18933 68564
rect 18891 68515 18933 68524
rect 18699 68480 18741 68489
rect 18699 68440 18700 68480
rect 18740 68440 18741 68480
rect 18699 68431 18741 68440
rect 19084 68321 19124 69028
rect 19564 68984 19604 68993
rect 19276 68944 19564 68984
rect 19276 68480 19316 68944
rect 19564 68935 19604 68944
rect 19372 68648 19412 68657
rect 19660 68648 19700 69868
rect 19756 69740 19796 69749
rect 19756 69497 19796 69700
rect 19755 69488 19797 69497
rect 19755 69448 19756 69488
rect 19796 69448 19797 69488
rect 19755 69439 19797 69448
rect 19755 69320 19797 69329
rect 19755 69280 19756 69320
rect 19796 69280 19797 69320
rect 19755 69271 19797 69280
rect 19756 69236 19796 69271
rect 19756 69185 19796 69196
rect 19412 68608 19700 68648
rect 19372 68599 19412 68608
rect 19228 68470 19316 68480
rect 19268 68440 19316 68470
rect 19228 68421 19268 68430
rect 19563 68396 19605 68405
rect 19563 68356 19564 68396
rect 19604 68356 19605 68396
rect 19563 68347 19605 68356
rect 19083 68312 19125 68321
rect 19083 68272 19084 68312
rect 19124 68272 19125 68312
rect 19083 68263 19125 68272
rect 19371 68312 19413 68321
rect 19371 68272 19372 68312
rect 19412 68272 19413 68312
rect 19371 68263 19413 68272
rect 18808 68060 19176 68069
rect 18848 68020 18890 68060
rect 18930 68020 18972 68060
rect 19012 68020 19054 68060
rect 19094 68020 19136 68060
rect 18808 68011 19176 68020
rect 18507 67724 18549 67733
rect 18507 67684 18508 67724
rect 18548 67684 18644 67724
rect 18507 67675 18549 67684
rect 18316 67348 18452 67388
rect 18123 65708 18165 65717
rect 18123 65668 18124 65708
rect 18164 65668 18165 65708
rect 18123 65659 18165 65668
rect 18124 65465 18164 65546
rect 18315 65540 18357 65549
rect 18315 65500 18316 65540
rect 18356 65500 18357 65540
rect 18315 65491 18357 65500
rect 18123 65456 18165 65465
rect 18123 65411 18124 65456
rect 18164 65411 18165 65456
rect 18123 65407 18165 65411
rect 18124 65402 18164 65407
rect 18316 65406 18356 65491
rect 18028 65248 18356 65288
rect 18123 64364 18165 64373
rect 18123 64324 18124 64364
rect 18164 64324 18165 64364
rect 18123 64315 18165 64324
rect 17740 64240 17876 64280
rect 17259 63232 17260 63272
rect 17300 63232 17301 63272
rect 17259 63223 17301 63232
rect 17452 63232 17588 63272
rect 17643 63272 17685 63281
rect 17643 63232 17644 63272
rect 17684 63232 17685 63272
rect 16971 63188 17013 63197
rect 16971 63148 16972 63188
rect 17012 63148 17013 63188
rect 16971 63139 17013 63148
rect 17163 63104 17205 63113
rect 17068 63064 17164 63104
rect 17204 63064 17205 63104
rect 16972 63020 17012 63029
rect 17068 63020 17108 63064
rect 17163 63055 17205 63064
rect 17012 62980 17108 63020
rect 16972 62971 17012 62980
rect 17163 62936 17205 62945
rect 17163 62896 17164 62936
rect 17204 62896 17205 62936
rect 17163 62887 17205 62896
rect 17164 61760 17204 62887
rect 17068 61720 17204 61760
rect 16875 59996 16917 60005
rect 16875 59956 16876 59996
rect 16916 59956 16917 59996
rect 16875 59947 16917 59956
rect 16971 59660 17013 59669
rect 16971 59620 16972 59660
rect 17012 59620 17013 59660
rect 16971 59611 17013 59620
rect 16875 59576 16917 59585
rect 16875 59536 16876 59576
rect 16916 59536 16917 59576
rect 16875 59527 16917 59536
rect 16876 59442 16916 59527
rect 16972 58829 17012 59611
rect 17068 59240 17108 61720
rect 17164 60920 17204 60929
rect 17164 60677 17204 60880
rect 17163 60668 17205 60677
rect 17163 60628 17164 60668
rect 17204 60628 17205 60668
rect 17163 60619 17205 60628
rect 17260 60593 17300 63223
rect 17452 63020 17492 63232
rect 17643 63223 17685 63232
rect 17547 63104 17589 63113
rect 17547 63064 17548 63104
rect 17588 63064 17589 63104
rect 17547 63055 17589 63064
rect 17644 63104 17684 63113
rect 17356 62980 17492 63020
rect 17259 60584 17301 60593
rect 17259 60544 17260 60584
rect 17300 60544 17301 60584
rect 17259 60535 17301 60544
rect 17356 60509 17396 62980
rect 17548 62970 17588 63055
rect 17644 62945 17684 63064
rect 17643 62936 17685 62945
rect 17643 62896 17644 62936
rect 17684 62896 17685 62936
rect 17643 62887 17685 62896
rect 17740 62441 17780 64240
rect 18027 64196 18069 64205
rect 18027 64156 18028 64196
rect 18068 64156 18069 64196
rect 18027 64147 18069 64156
rect 17932 63860 17972 63871
rect 17932 63785 17972 63820
rect 18028 63860 18068 64147
rect 17931 63776 17973 63785
rect 17931 63736 17932 63776
rect 17972 63736 17973 63776
rect 17931 63727 17973 63736
rect 18028 63365 18068 63820
rect 18027 63356 18069 63365
rect 18027 63316 18028 63356
rect 18068 63316 18069 63356
rect 18027 63307 18069 63316
rect 18027 63104 18069 63113
rect 17932 63064 18028 63104
rect 18068 63064 18069 63104
rect 17739 62432 17781 62441
rect 17739 62392 17740 62432
rect 17780 62392 17781 62432
rect 17739 62383 17781 62392
rect 17452 61592 17492 61601
rect 17452 61349 17492 61552
rect 17644 61424 17684 61433
rect 17451 61340 17493 61349
rect 17451 61300 17452 61340
rect 17492 61300 17493 61340
rect 17451 61291 17493 61300
rect 17644 60915 17684 61384
rect 17644 60866 17684 60875
rect 17355 60500 17397 60509
rect 17355 60460 17356 60500
rect 17396 60460 17397 60500
rect 17355 60451 17397 60460
rect 17163 60332 17205 60341
rect 17163 60292 17164 60332
rect 17204 60292 17205 60332
rect 17163 60283 17205 60292
rect 17451 60332 17493 60341
rect 17451 60292 17452 60332
rect 17492 60292 17493 60332
rect 17451 60283 17493 60292
rect 17068 59081 17108 59200
rect 17067 59072 17109 59081
rect 17067 59032 17068 59072
rect 17108 59032 17109 59072
rect 17067 59023 17109 59032
rect 16971 58820 17013 58829
rect 16971 58780 16972 58820
rect 17012 58780 17013 58820
rect 16971 58771 17013 58780
rect 16780 58696 16916 58736
rect 16779 58568 16821 58577
rect 16779 58528 16780 58568
rect 16820 58528 16821 58568
rect 16779 58519 16821 58528
rect 16780 58434 16820 58519
rect 16779 57896 16821 57905
rect 16779 57856 16780 57896
rect 16820 57856 16821 57896
rect 16779 57847 16821 57856
rect 16683 56972 16725 56981
rect 16683 56932 16684 56972
rect 16724 56932 16725 56972
rect 16683 56923 16725 56932
rect 16683 56552 16725 56561
rect 16683 56512 16684 56552
rect 16724 56512 16725 56552
rect 16683 56503 16725 56512
rect 16684 56418 16724 56503
rect 16780 56393 16820 57847
rect 16876 56813 16916 58696
rect 16972 58568 17012 58771
rect 16972 58519 17012 58528
rect 17068 58568 17108 58577
rect 17164 58568 17204 60283
rect 17452 60198 17492 60283
rect 17259 60080 17301 60089
rect 17259 60040 17260 60080
rect 17300 60040 17301 60080
rect 17259 60031 17301 60040
rect 17260 59946 17300 60031
rect 17643 59996 17685 60005
rect 17643 59956 17644 59996
rect 17684 59956 17685 59996
rect 17643 59947 17685 59956
rect 17452 59408 17492 59417
rect 17356 59368 17452 59408
rect 17259 59156 17301 59165
rect 17259 59116 17260 59156
rect 17300 59116 17301 59156
rect 17259 59107 17301 59116
rect 17108 58528 17204 58568
rect 17068 58519 17108 58528
rect 17260 58400 17300 59107
rect 17260 58351 17300 58360
rect 17163 58064 17205 58073
rect 17163 58024 17164 58064
rect 17204 58024 17205 58064
rect 17163 58015 17205 58024
rect 17164 57896 17204 58015
rect 17356 57980 17396 59368
rect 17452 59359 17492 59368
rect 17548 59408 17588 59417
rect 17548 59081 17588 59368
rect 17547 59072 17589 59081
rect 17547 59032 17548 59072
rect 17588 59032 17589 59072
rect 17547 59023 17589 59032
rect 17644 58577 17684 59947
rect 17740 59240 17780 62383
rect 17835 61088 17877 61097
rect 17835 61048 17836 61088
rect 17876 61048 17877 61088
rect 17835 61039 17877 61048
rect 17836 60954 17876 61039
rect 17932 59408 17972 63064
rect 18027 63055 18069 63064
rect 18124 63104 18164 64315
rect 18028 62970 18068 63055
rect 18028 62441 18068 62526
rect 18027 62432 18069 62441
rect 18027 62392 18028 62432
rect 18068 62392 18069 62432
rect 18027 62383 18069 62392
rect 18124 62264 18164 63064
rect 17932 59359 17972 59368
rect 18028 62224 18164 62264
rect 18028 59408 18068 62224
rect 18124 60920 18164 60929
rect 18124 60341 18164 60880
rect 18220 60920 18260 60929
rect 18220 60509 18260 60880
rect 18219 60500 18261 60509
rect 18219 60460 18220 60500
rect 18260 60460 18261 60500
rect 18219 60451 18261 60460
rect 18123 60332 18165 60341
rect 18123 60292 18124 60332
rect 18164 60292 18165 60332
rect 18123 60283 18165 60292
rect 18124 60080 18164 60089
rect 18124 59753 18164 60040
rect 18219 59912 18261 59921
rect 18219 59872 18220 59912
rect 18260 59872 18261 59912
rect 18219 59863 18261 59872
rect 18123 59744 18165 59753
rect 18123 59704 18124 59744
rect 18164 59704 18165 59744
rect 18123 59695 18165 59704
rect 18028 59359 18068 59368
rect 17740 59200 18068 59240
rect 17643 58568 17685 58577
rect 17643 58528 17644 58568
rect 17684 58528 17685 58568
rect 17643 58519 17685 58528
rect 17644 58434 17684 58519
rect 17547 58148 17589 58157
rect 17547 58108 17548 58148
rect 17588 58108 17589 58148
rect 17547 58099 17589 58108
rect 17356 57931 17396 57940
rect 17548 57905 17588 58099
rect 18028 57989 18068 59200
rect 18027 57980 18069 57989
rect 18027 57940 18028 57980
rect 18068 57940 18069 57980
rect 18027 57931 18069 57940
rect 17068 57856 17164 57896
rect 16875 56804 16917 56813
rect 16875 56764 16876 56804
rect 16916 56764 16917 56804
rect 16875 56755 16917 56764
rect 16779 56384 16821 56393
rect 16779 56344 16780 56384
rect 16820 56344 16821 56384
rect 16779 56335 16821 56344
rect 16876 56384 16916 56755
rect 16876 56309 16916 56344
rect 16971 56384 17013 56393
rect 16971 56344 16972 56384
rect 17012 56344 17013 56384
rect 16971 56335 17013 56344
rect 16875 56300 16917 56309
rect 16875 56260 16876 56300
rect 16916 56260 16917 56300
rect 16875 56251 16917 56260
rect 16876 56220 16916 56251
rect 16972 56250 17012 56335
rect 16971 55544 17013 55553
rect 17068 55544 17108 57856
rect 17164 57847 17204 57856
rect 17547 57896 17589 57905
rect 17547 57856 17548 57896
rect 17588 57856 17589 57896
rect 17547 57847 17589 57856
rect 17644 57896 17684 57905
rect 17548 57762 17588 57847
rect 17644 57821 17684 57856
rect 17740 57896 17780 57905
rect 17643 57812 17685 57821
rect 17643 57772 17644 57812
rect 17684 57772 17685 57812
rect 17643 57763 17685 57772
rect 17163 57728 17205 57737
rect 17163 57688 17164 57728
rect 17204 57688 17205 57728
rect 17163 57679 17205 57688
rect 17164 56552 17204 57679
rect 17548 57056 17588 57067
rect 17548 56981 17588 57016
rect 17547 56972 17589 56981
rect 17547 56932 17548 56972
rect 17588 56932 17589 56972
rect 17547 56923 17589 56932
rect 17644 56720 17684 57763
rect 17740 57737 17780 57856
rect 17835 57896 17877 57905
rect 17835 57856 17836 57896
rect 17876 57856 17877 57896
rect 17835 57847 17877 57856
rect 18124 57896 18164 57907
rect 17836 57762 17876 57847
rect 18124 57821 18164 57856
rect 18123 57812 18165 57821
rect 18123 57772 18124 57812
rect 18164 57772 18165 57812
rect 18123 57763 18165 57772
rect 17739 57728 17781 57737
rect 17739 57688 17740 57728
rect 17780 57688 17781 57728
rect 17739 57679 17781 57688
rect 17739 57560 17781 57569
rect 17739 57520 17740 57560
rect 17780 57520 17781 57560
rect 17739 57511 17781 57520
rect 17740 57308 17780 57511
rect 17740 57259 17780 57268
rect 18123 57308 18165 57317
rect 18123 57268 18124 57308
rect 18164 57268 18165 57308
rect 18123 57259 18165 57268
rect 17931 57224 17973 57233
rect 17931 57184 17932 57224
rect 17972 57184 17973 57224
rect 17931 57175 17973 57184
rect 17932 57056 17972 57175
rect 18027 57140 18069 57149
rect 18027 57100 18028 57140
rect 18068 57100 18069 57140
rect 18027 57091 18069 57100
rect 17932 57007 17972 57016
rect 18028 57006 18068 57091
rect 18124 57056 18164 57259
rect 18220 57056 18260 59863
rect 18316 58073 18356 65248
rect 18412 58745 18452 67348
rect 18507 66968 18549 66977
rect 18507 66928 18508 66968
rect 18548 66928 18549 66968
rect 18507 66919 18549 66928
rect 18508 66834 18548 66919
rect 18508 66128 18548 66137
rect 18604 66128 18644 67684
rect 19372 67640 19412 68263
rect 19564 68262 19604 68347
rect 19756 68228 19796 68237
rect 19660 68188 19756 68228
rect 19660 67649 19700 68188
rect 19756 68179 19796 68188
rect 19756 67724 19796 67733
rect 19372 67591 19412 67600
rect 19659 67640 19701 67649
rect 19659 67600 19660 67640
rect 19700 67600 19701 67640
rect 19659 67591 19701 67600
rect 19564 67472 19604 67481
rect 19276 67432 19564 67472
rect 18548 66088 18644 66128
rect 18508 66079 18548 66088
rect 18604 64205 18644 66088
rect 18700 66716 18740 66725
rect 18700 65465 18740 66676
rect 18808 66548 19176 66557
rect 18848 66508 18890 66548
rect 18930 66508 18972 66548
rect 19012 66508 19054 66548
rect 19094 66508 19136 66548
rect 18808 66499 19176 66508
rect 19036 66137 19076 66146
rect 19276 66128 19316 67432
rect 19564 67423 19604 67432
rect 19756 67145 19796 67684
rect 19755 67136 19797 67145
rect 19755 67096 19756 67136
rect 19796 67096 19797 67136
rect 19755 67087 19797 67096
rect 19852 67136 19892 73060
rect 19948 72764 19988 72773
rect 19948 72269 19988 72724
rect 19947 72260 19989 72269
rect 19947 72220 19948 72260
rect 19988 72220 19989 72260
rect 19947 72211 19989 72220
rect 19948 72008 19988 72017
rect 19948 71588 19988 71968
rect 20048 71840 20416 71849
rect 20088 71800 20130 71840
rect 20170 71800 20212 71840
rect 20252 71800 20294 71840
rect 20334 71800 20376 71840
rect 20048 71791 20416 71800
rect 19948 71548 20084 71588
rect 19947 71420 19989 71429
rect 19947 71380 19948 71420
rect 19988 71380 19989 71420
rect 19947 71371 19989 71380
rect 19948 71286 19988 71371
rect 19947 70832 19989 70841
rect 19947 70792 19948 70832
rect 19988 70792 19989 70832
rect 19947 70783 19989 70792
rect 19948 70698 19988 70783
rect 20044 70673 20084 71548
rect 20140 71252 20180 71261
rect 20043 70664 20085 70673
rect 20043 70624 20044 70664
rect 20084 70624 20085 70664
rect 20043 70615 20085 70624
rect 20140 70589 20180 71212
rect 20139 70580 20181 70589
rect 20139 70540 20140 70580
rect 20180 70540 20181 70580
rect 20139 70531 20181 70540
rect 20048 70328 20416 70337
rect 20088 70288 20130 70328
rect 20170 70288 20212 70328
rect 20252 70288 20294 70328
rect 20334 70288 20376 70328
rect 20048 70279 20416 70288
rect 20043 70076 20085 70085
rect 20043 70036 20044 70076
rect 20084 70036 20085 70076
rect 20043 70027 20085 70036
rect 19948 69908 19988 69917
rect 19948 69161 19988 69868
rect 20044 69665 20084 70027
rect 20139 69740 20181 69749
rect 20139 69700 20140 69740
rect 20180 69700 20181 69740
rect 20139 69691 20181 69700
rect 20043 69656 20085 69665
rect 20043 69616 20044 69656
rect 20084 69616 20085 69656
rect 20043 69607 20085 69616
rect 20140 69606 20180 69691
rect 20043 69488 20085 69497
rect 20043 69448 20044 69488
rect 20084 69448 20085 69488
rect 20043 69439 20085 69448
rect 19947 69152 19989 69161
rect 19947 69112 19948 69152
rect 19988 69112 19989 69152
rect 19947 69103 19989 69112
rect 20044 68993 20084 69439
rect 19948 68984 19988 68993
rect 19948 68564 19988 68944
rect 20043 68984 20085 68993
rect 20043 68944 20044 68984
rect 20084 68944 20085 68984
rect 20043 68935 20085 68944
rect 20048 68816 20416 68825
rect 20088 68776 20130 68816
rect 20170 68776 20212 68816
rect 20252 68776 20294 68816
rect 20334 68776 20376 68816
rect 20048 68767 20416 68776
rect 19948 68524 20084 68564
rect 19948 68396 19988 68405
rect 19948 67985 19988 68356
rect 20044 68321 20084 68524
rect 20043 68312 20085 68321
rect 20043 68272 20044 68312
rect 20084 68272 20085 68312
rect 20043 68263 20085 68272
rect 20140 68228 20180 68237
rect 19947 67976 19989 67985
rect 19947 67936 19948 67976
rect 19988 67936 19989 67976
rect 19947 67927 19989 67936
rect 20140 67481 20180 68188
rect 19852 67087 19892 67096
rect 19948 67472 19988 67481
rect 19948 66977 19988 67432
rect 20139 67472 20181 67481
rect 20139 67432 20140 67472
rect 20180 67432 20181 67472
rect 20139 67423 20181 67432
rect 20048 67304 20416 67313
rect 20088 67264 20130 67304
rect 20170 67264 20212 67304
rect 20252 67264 20294 67304
rect 20334 67264 20376 67304
rect 20048 67255 20416 67264
rect 20236 67136 20276 67145
rect 20524 67136 20564 84391
rect 20619 84104 20661 84113
rect 20619 84064 20620 84104
rect 20660 84064 20661 84104
rect 20619 84055 20661 84064
rect 20620 80585 20660 84055
rect 21387 82760 21429 82769
rect 21387 82720 21388 82760
rect 21428 82720 21429 82760
rect 21387 82711 21429 82720
rect 21388 82265 21428 82711
rect 21387 82256 21429 82265
rect 21387 82216 21388 82256
rect 21428 82216 21429 82256
rect 21387 82207 21429 82216
rect 20619 80576 20661 80585
rect 20619 80536 20620 80576
rect 20660 80536 20661 80576
rect 20619 80527 20661 80536
rect 20619 76544 20661 76553
rect 20619 76504 20620 76544
rect 20660 76504 20661 76544
rect 20619 76495 20661 76504
rect 20620 75377 20660 76495
rect 20715 75788 20757 75797
rect 20715 75748 20716 75788
rect 20756 75748 20757 75788
rect 20715 75739 20757 75748
rect 20619 75368 20661 75377
rect 20619 75328 20620 75368
rect 20660 75328 20661 75368
rect 20619 75319 20661 75328
rect 20716 74369 20756 75739
rect 20715 74360 20757 74369
rect 20715 74320 20716 74360
rect 20756 74320 20757 74360
rect 20715 74311 20757 74320
rect 20619 72092 20661 72101
rect 20619 72052 20620 72092
rect 20660 72052 20661 72092
rect 20619 72043 20661 72052
rect 20620 71009 20660 72043
rect 20619 71000 20661 71009
rect 20619 70960 20620 71000
rect 20660 70960 20661 71000
rect 20619 70951 20661 70960
rect 21387 70832 21429 70841
rect 21387 70792 21388 70832
rect 21428 70792 21429 70832
rect 21387 70783 21429 70792
rect 20619 69740 20661 69749
rect 20619 69700 20620 69740
rect 20660 69700 20661 69740
rect 20619 69691 20661 69700
rect 20620 67985 20660 69691
rect 21388 68993 21428 70783
rect 21387 68984 21429 68993
rect 21387 68944 21388 68984
rect 21428 68944 21429 68984
rect 21387 68935 21429 68944
rect 20619 67976 20661 67985
rect 20619 67936 20620 67976
rect 20660 67936 20661 67976
rect 20619 67927 20661 67936
rect 20276 67096 20564 67136
rect 20236 67087 20276 67096
rect 19947 66968 19989 66977
rect 19947 66928 19948 66968
rect 19988 66928 19989 66968
rect 19947 66919 19989 66928
rect 19660 66884 19700 66893
rect 19467 66632 19509 66641
rect 19467 66592 19468 66632
rect 19508 66592 19509 66632
rect 19467 66583 19509 66592
rect 19076 66097 19316 66128
rect 19036 66088 19316 66097
rect 19372 66212 19412 66221
rect 19179 65960 19221 65969
rect 19179 65920 19180 65960
rect 19220 65920 19221 65960
rect 19179 65911 19221 65920
rect 19180 65826 19220 65911
rect 19372 65549 19412 66172
rect 19371 65540 19413 65549
rect 19371 65500 19372 65540
rect 19412 65500 19413 65540
rect 19371 65491 19413 65500
rect 18699 65456 18741 65465
rect 18699 65416 18700 65456
rect 18740 65416 18741 65456
rect 19468 65456 19508 66583
rect 19660 66305 19700 66844
rect 20044 66884 20084 66893
rect 19659 66296 19701 66305
rect 19659 66256 19660 66296
rect 19700 66256 19701 66296
rect 19659 66247 19701 66256
rect 19947 66296 19989 66305
rect 19947 66256 19948 66296
rect 19988 66256 19989 66296
rect 19947 66247 19989 66256
rect 19755 66212 19797 66221
rect 19755 66172 19756 66212
rect 19796 66172 19797 66212
rect 19755 66163 19797 66172
rect 19756 66078 19796 66163
rect 19948 66162 19988 66247
rect 19563 65960 19605 65969
rect 20044 65960 20084 66844
rect 19563 65920 19564 65960
rect 19604 65920 19605 65960
rect 19563 65911 19605 65920
rect 19852 65920 20084 65960
rect 19564 65826 19604 65911
rect 19468 65416 19604 65456
rect 18699 65407 18741 65416
rect 18988 65372 19028 65383
rect 18988 65297 19028 65332
rect 19372 65372 19412 65381
rect 19412 65332 19508 65372
rect 19372 65323 19412 65332
rect 18987 65288 19029 65297
rect 18987 65248 18988 65288
rect 19028 65248 19029 65288
rect 18987 65239 19029 65248
rect 19180 65204 19220 65213
rect 19220 65164 19316 65204
rect 19180 65155 19220 65164
rect 18808 65036 19176 65045
rect 18848 64996 18890 65036
rect 18930 64996 18972 65036
rect 19012 64996 19054 65036
rect 19094 64996 19136 65036
rect 18808 64987 19176 64996
rect 19276 64961 19316 65164
rect 19275 64952 19317 64961
rect 19275 64912 19276 64952
rect 19316 64912 19317 64952
rect 19275 64903 19317 64912
rect 19372 64700 19412 64709
rect 18988 64616 19028 64627
rect 18988 64541 19028 64576
rect 18987 64532 19029 64541
rect 18987 64492 18988 64532
rect 19028 64492 19029 64532
rect 18987 64483 19029 64492
rect 19180 64448 19220 64457
rect 19180 64280 19220 64408
rect 19372 64280 19412 64660
rect 19084 64240 19220 64280
rect 19276 64240 19412 64280
rect 18603 64196 18645 64205
rect 18603 64156 18604 64196
rect 18644 64156 18645 64196
rect 18603 64147 18645 64156
rect 18507 63944 18549 63953
rect 19084 63944 19124 64240
rect 19180 64112 19220 64121
rect 19276 64112 19316 64240
rect 19468 64121 19508 65332
rect 19564 65288 19604 65416
rect 19755 65372 19797 65381
rect 19755 65332 19756 65372
rect 19796 65332 19797 65372
rect 19755 65323 19797 65332
rect 19564 65239 19604 65248
rect 19756 65238 19796 65323
rect 19852 64877 19892 65920
rect 20048 65792 20416 65801
rect 20088 65752 20130 65792
rect 20170 65752 20212 65792
rect 20252 65752 20294 65792
rect 20334 65752 20376 65792
rect 20048 65743 20416 65752
rect 19947 65624 19989 65633
rect 19947 65584 19948 65624
rect 19988 65584 19989 65624
rect 19947 65575 19989 65584
rect 19948 65288 19988 65575
rect 19948 65239 19988 65248
rect 20043 65288 20085 65297
rect 20043 65248 20044 65288
rect 20084 65248 20085 65288
rect 20043 65239 20085 65248
rect 19851 64868 19893 64877
rect 19851 64828 19852 64868
rect 19892 64828 19893 64868
rect 19851 64819 19893 64828
rect 19948 64868 19988 64877
rect 20044 64868 20084 65239
rect 19988 64828 20084 64868
rect 19948 64819 19988 64828
rect 19756 64700 19796 64709
rect 19563 64616 19605 64625
rect 19563 64576 19564 64616
rect 19604 64576 19605 64616
rect 19563 64567 19605 64576
rect 19564 64448 19604 64567
rect 19659 64532 19701 64541
rect 19659 64492 19660 64532
rect 19700 64492 19701 64532
rect 19659 64483 19701 64492
rect 19564 64399 19604 64408
rect 19220 64072 19316 64112
rect 19467 64112 19509 64121
rect 19467 64072 19468 64112
rect 19508 64072 19509 64112
rect 19180 64063 19220 64072
rect 19467 64063 19509 64072
rect 19371 64028 19413 64037
rect 19371 63988 19372 64028
rect 19412 63988 19413 64028
rect 19371 63979 19413 63988
rect 18507 63904 18508 63944
rect 18548 63904 18740 63944
rect 18507 63895 18549 63904
rect 18508 63810 18548 63895
rect 18604 63104 18644 63113
rect 18507 63020 18549 63029
rect 18604 63020 18644 63064
rect 18507 62980 18508 63020
rect 18548 62980 18644 63020
rect 18507 62971 18549 62980
rect 18508 62273 18548 62971
rect 18700 62936 18740 63904
rect 19036 63934 19124 63944
rect 19076 63904 19124 63934
rect 19036 63885 19076 63894
rect 19372 63860 19412 63979
rect 19563 63944 19605 63953
rect 19563 63904 19564 63944
rect 19604 63904 19605 63944
rect 19563 63895 19605 63904
rect 19372 63811 19412 63820
rect 19564 63776 19604 63895
rect 19564 63727 19604 63736
rect 18808 63524 19176 63533
rect 18848 63484 18890 63524
rect 18930 63484 18972 63524
rect 19012 63484 19054 63524
rect 19094 63484 19136 63524
rect 18808 63475 19176 63484
rect 19660 63440 19700 64483
rect 19756 64457 19796 64660
rect 19755 64448 19797 64457
rect 19755 64408 19756 64448
rect 19796 64408 19797 64448
rect 19755 64399 19797 64408
rect 19947 64280 19989 64289
rect 19947 64240 19948 64280
rect 19988 64240 19989 64280
rect 19947 64231 19989 64240
rect 20048 64280 20416 64289
rect 20088 64240 20130 64280
rect 20170 64240 20212 64280
rect 20252 64240 20294 64280
rect 20334 64240 20376 64280
rect 20048 64231 20416 64240
rect 19948 64112 19988 64231
rect 19948 64063 19988 64072
rect 19755 63860 19797 63869
rect 19755 63820 19756 63860
rect 19796 63820 19797 63860
rect 19755 63811 19797 63820
rect 19756 63726 19796 63811
rect 19947 63608 19989 63617
rect 19947 63568 19948 63608
rect 19988 63568 19989 63608
rect 19947 63559 19989 63568
rect 19564 63400 19700 63440
rect 19468 63188 19508 63197
rect 19132 63113 19172 63122
rect 19172 63073 19220 63104
rect 19132 63064 19220 63073
rect 18604 62896 18740 62936
rect 18507 62264 18549 62273
rect 18507 62224 18508 62264
rect 18548 62224 18549 62264
rect 18507 62215 18549 62224
rect 18508 59408 18548 62215
rect 18604 61853 18644 62896
rect 19180 62684 19220 63064
rect 19276 63020 19316 63029
rect 19468 63020 19508 63148
rect 19316 62980 19508 63020
rect 19276 62971 19316 62980
rect 19180 62644 19508 62684
rect 19468 62600 19508 62644
rect 19468 62551 19508 62560
rect 19276 62432 19316 62441
rect 19564 62432 19604 63400
rect 19659 63272 19701 63281
rect 19659 63232 19660 63272
rect 19700 63232 19701 63272
rect 19659 63223 19701 63232
rect 19660 63138 19700 63223
rect 19659 62684 19701 62693
rect 19659 62644 19660 62684
rect 19700 62644 19701 62684
rect 19659 62635 19701 62644
rect 19316 62392 19604 62432
rect 18699 62264 18741 62273
rect 18699 62224 18700 62264
rect 18740 62224 18741 62264
rect 18699 62215 18741 62224
rect 18603 61844 18645 61853
rect 18603 61804 18604 61844
rect 18644 61804 18645 61844
rect 18603 61795 18645 61804
rect 18700 61760 18740 62215
rect 18808 62012 19176 62021
rect 18848 61972 18890 62012
rect 18930 61972 18972 62012
rect 19012 61972 19054 62012
rect 19094 61972 19136 62012
rect 18808 61963 19176 61972
rect 18796 61760 18836 61769
rect 18700 61720 18796 61760
rect 18796 61711 18836 61720
rect 19083 61760 19125 61769
rect 19083 61720 19084 61760
rect 19124 61720 19125 61760
rect 19083 61711 19125 61720
rect 18603 61676 18645 61685
rect 18603 61636 18604 61676
rect 18644 61636 18645 61676
rect 18603 61627 18645 61636
rect 18988 61676 19028 61685
rect 18604 61542 18644 61627
rect 18988 61097 19028 61636
rect 18987 61088 19029 61097
rect 18987 61048 18988 61088
rect 19028 61048 19029 61088
rect 18987 61039 19029 61048
rect 19084 60920 19124 61711
rect 19179 61592 19221 61601
rect 19179 61552 19180 61592
rect 19220 61552 19221 61592
rect 19179 61543 19221 61552
rect 19180 61424 19220 61543
rect 19180 61375 19220 61384
rect 19180 60920 19220 60929
rect 19084 60880 19180 60920
rect 18604 60836 18644 60847
rect 18604 60761 18644 60796
rect 18700 60836 18740 60845
rect 18603 60752 18645 60761
rect 18603 60712 18604 60752
rect 18644 60712 18645 60752
rect 18603 60703 18645 60712
rect 18603 60584 18645 60593
rect 18700 60584 18740 60796
rect 19180 60677 19220 60880
rect 19179 60668 19221 60677
rect 19179 60628 19180 60668
rect 19220 60628 19221 60668
rect 19179 60619 19221 60628
rect 18603 60544 18604 60584
rect 18644 60544 18740 60584
rect 18603 60535 18645 60544
rect 18508 59333 18548 59368
rect 18507 59324 18549 59333
rect 18507 59284 18508 59324
rect 18548 59284 18549 59324
rect 18507 59275 18549 59284
rect 18411 58736 18453 58745
rect 18411 58696 18412 58736
rect 18452 58696 18453 58736
rect 18411 58687 18453 58696
rect 18315 58064 18357 58073
rect 18315 58024 18316 58064
rect 18356 58024 18452 58064
rect 18315 58015 18357 58024
rect 18412 57896 18452 58024
rect 18508 57938 18548 57947
rect 18412 57847 18452 57856
rect 18503 57898 18508 57923
rect 18604 57923 18644 60535
rect 18808 60500 19176 60509
rect 18848 60460 18890 60500
rect 18930 60460 18972 60500
rect 19012 60460 19054 60500
rect 19094 60460 19136 60500
rect 18808 60451 19176 60460
rect 19276 60080 19316 62392
rect 19660 62348 19700 62635
rect 19851 62600 19893 62609
rect 19851 62560 19852 62600
rect 19892 62560 19893 62600
rect 19851 62551 19893 62560
rect 19852 62466 19892 62551
rect 19660 62299 19700 62308
rect 19948 62096 19988 63559
rect 20523 62936 20565 62945
rect 20523 62896 20524 62936
rect 20564 62896 20565 62936
rect 20523 62887 20565 62896
rect 20048 62768 20416 62777
rect 20088 62728 20130 62768
rect 20170 62728 20212 62768
rect 20252 62728 20294 62768
rect 20334 62728 20376 62768
rect 20048 62719 20416 62728
rect 20236 62600 20276 62609
rect 20524 62600 20564 62887
rect 20276 62560 20564 62600
rect 20236 62551 20276 62560
rect 20043 62348 20085 62357
rect 20043 62308 20044 62348
rect 20084 62308 20085 62348
rect 20043 62299 20085 62308
rect 20044 62214 20084 62299
rect 19852 62056 19988 62096
rect 19372 61676 19412 61685
rect 19372 61181 19412 61636
rect 19756 61676 19796 61685
rect 19563 61424 19605 61433
rect 19563 61384 19564 61424
rect 19604 61384 19605 61424
rect 19563 61375 19605 61384
rect 19564 61290 19604 61375
rect 19371 61172 19413 61181
rect 19371 61132 19372 61172
rect 19412 61132 19413 61172
rect 19371 61123 19413 61132
rect 19756 61088 19796 61636
rect 19852 61256 19892 62056
rect 19947 61928 19989 61937
rect 19947 61888 19948 61928
rect 19988 61888 19989 61928
rect 19947 61879 19989 61888
rect 19948 61760 19988 61879
rect 19948 61711 19988 61720
rect 20048 61256 20416 61265
rect 19852 61216 19988 61256
rect 19852 61088 19892 61097
rect 19756 61048 19852 61088
rect 19852 61039 19892 61048
rect 19467 60920 19509 60929
rect 19467 60880 19468 60920
rect 19508 60880 19509 60920
rect 19467 60871 19509 60880
rect 19660 60906 19700 60915
rect 19371 60080 19413 60089
rect 19276 60040 19372 60080
rect 19412 60040 19413 60080
rect 19371 60031 19413 60040
rect 19372 59946 19412 60031
rect 19180 59585 19220 59670
rect 19179 59576 19221 59585
rect 19179 59536 19180 59576
rect 19220 59536 19221 59576
rect 19179 59527 19221 59536
rect 19036 59398 19076 59407
rect 19076 59358 19316 59394
rect 19036 59354 19316 59358
rect 19036 59349 19076 59354
rect 18808 58988 19176 58997
rect 18848 58948 18890 58988
rect 18930 58948 18972 58988
rect 19012 58948 19054 58988
rect 19094 58948 19136 58988
rect 18808 58939 19176 58948
rect 19084 58820 19124 58829
rect 19276 58820 19316 59354
rect 19371 59324 19413 59333
rect 19371 59284 19372 59324
rect 19412 59284 19413 59324
rect 19371 59275 19413 59284
rect 19372 59190 19412 59275
rect 19124 58780 19316 58820
rect 19468 58820 19508 60871
rect 19564 60332 19604 60341
rect 19660 60332 19700 60866
rect 19604 60292 19700 60332
rect 19564 60283 19604 60292
rect 19756 60164 19796 60173
rect 19756 59837 19796 60124
rect 19948 60080 19988 61216
rect 20088 61216 20130 61256
rect 20170 61216 20212 61256
rect 20252 61216 20294 61256
rect 20334 61216 20376 61256
rect 20048 61207 20416 61216
rect 20043 60836 20085 60845
rect 20043 60796 20044 60836
rect 20084 60796 20085 60836
rect 20043 60787 20085 60796
rect 20044 60702 20084 60787
rect 20236 60668 20276 60677
rect 20236 60257 20276 60628
rect 21003 60584 21045 60593
rect 21003 60544 21004 60584
rect 21044 60544 21045 60584
rect 21003 60535 21045 60544
rect 20235 60248 20277 60257
rect 20235 60208 20236 60248
rect 20276 60208 20277 60248
rect 20235 60199 20277 60208
rect 19852 60040 19988 60080
rect 19755 59828 19797 59837
rect 19755 59788 19756 59828
rect 19796 59788 19797 59828
rect 19755 59779 19797 59788
rect 19852 59576 19892 60040
rect 19947 59912 19989 59921
rect 19947 59872 19948 59912
rect 19988 59872 19989 59912
rect 19947 59863 19989 59872
rect 19948 59778 19988 59863
rect 20048 59744 20416 59753
rect 20088 59704 20130 59744
rect 20170 59704 20212 59744
rect 20252 59704 20294 59744
rect 20334 59704 20376 59744
rect 20048 59695 20416 59704
rect 19564 59536 19892 59576
rect 19947 59576 19989 59585
rect 19947 59536 19948 59576
rect 19988 59536 19989 59576
rect 19564 59240 19604 59536
rect 19947 59527 19989 59536
rect 19948 59442 19988 59527
rect 19851 59408 19893 59417
rect 19851 59368 19852 59408
rect 19892 59368 19893 59408
rect 19851 59359 19893 59368
rect 19755 59324 19797 59333
rect 19755 59284 19756 59324
rect 19796 59284 19797 59324
rect 19755 59275 19797 59284
rect 19564 59191 19604 59200
rect 19756 59190 19796 59275
rect 19564 58820 19604 58829
rect 19468 58780 19564 58820
rect 19084 58771 19124 58780
rect 19564 58771 19604 58780
rect 18795 58736 18837 58745
rect 18795 58696 18796 58736
rect 18836 58696 18837 58736
rect 18795 58687 18837 58696
rect 18548 57898 18644 57923
rect 18503 57883 18644 57898
rect 18503 57728 18543 57883
rect 18796 57812 18836 58687
rect 19372 58652 19412 58661
rect 19755 58652 19797 58661
rect 19412 58612 19604 58652
rect 19372 58603 19412 58612
rect 18892 58568 18932 58577
rect 18892 57989 18932 58528
rect 19180 58024 19412 58064
rect 18891 57980 18933 57989
rect 18891 57940 18892 57980
rect 18932 57940 18933 57980
rect 18891 57931 18933 57940
rect 18988 57896 19028 57907
rect 18988 57821 19028 57856
rect 19083 57896 19125 57905
rect 19083 57856 19084 57896
rect 19124 57856 19125 57896
rect 19083 57847 19125 57856
rect 19180 57896 19220 58024
rect 19372 57980 19412 58024
rect 19372 57940 19508 57980
rect 19180 57847 19220 57856
rect 19276 57896 19316 57905
rect 18412 57688 18543 57728
rect 18604 57772 18836 57812
rect 18987 57812 19029 57821
rect 18987 57772 18988 57812
rect 19028 57772 19029 57812
rect 18316 57056 18356 57065
rect 18220 57016 18316 57056
rect 18124 57007 18164 57016
rect 18316 57007 18356 57016
rect 17740 56897 17780 56982
rect 17739 56888 17781 56897
rect 17739 56848 17740 56888
rect 17780 56848 17781 56888
rect 17739 56839 17781 56848
rect 17931 56888 17973 56897
rect 18412 56888 18452 57688
rect 17931 56848 17932 56888
rect 17972 56848 17973 56888
rect 17931 56839 17973 56848
rect 18220 56848 18452 56888
rect 17644 56680 17780 56720
rect 17644 56552 17684 56561
rect 17164 56503 17204 56512
rect 17548 56512 17644 56552
rect 17356 56384 17396 56395
rect 17356 56309 17396 56344
rect 17452 56384 17492 56393
rect 17355 56300 17397 56309
rect 17355 56260 17356 56300
rect 17396 56260 17397 56300
rect 17355 56251 17397 56260
rect 17452 55805 17492 56344
rect 17163 55796 17205 55805
rect 17163 55756 17164 55796
rect 17204 55756 17205 55796
rect 17163 55747 17205 55756
rect 17451 55796 17493 55805
rect 17451 55756 17452 55796
rect 17492 55756 17493 55796
rect 17451 55747 17493 55756
rect 17164 55662 17204 55747
rect 16971 55504 16972 55544
rect 17012 55504 17108 55544
rect 16971 55495 17013 55504
rect 16588 55420 16820 55460
rect 16684 54872 16724 54881
rect 16588 54832 16684 54872
rect 16588 54209 16628 54832
rect 16684 54823 16724 54832
rect 16683 54620 16725 54629
rect 16683 54580 16684 54620
rect 16724 54580 16725 54620
rect 16683 54571 16725 54580
rect 16684 54486 16724 54571
rect 16587 54200 16629 54209
rect 16587 54160 16588 54200
rect 16628 54160 16629 54200
rect 16587 54151 16629 54160
rect 16683 54116 16725 54125
rect 16683 54076 16684 54116
rect 16724 54076 16725 54116
rect 16683 54067 16725 54076
rect 16684 54032 16724 54067
rect 16684 53981 16724 53992
rect 16780 53705 16820 55420
rect 16972 55410 17012 55495
rect 17452 55460 17492 55747
rect 17548 55637 17588 56512
rect 17644 56503 17684 56512
rect 17740 56393 17780 56680
rect 17739 56384 17781 56393
rect 17739 56344 17740 56384
rect 17780 56344 17781 56384
rect 17739 56335 17781 56344
rect 17932 56384 17972 56839
rect 18027 56720 18069 56729
rect 18027 56680 18028 56720
rect 18068 56680 18069 56720
rect 18027 56671 18069 56680
rect 17932 56335 17972 56344
rect 18028 56384 18068 56671
rect 18028 56335 18068 56344
rect 18220 56057 18260 56848
rect 18508 56384 18548 56393
rect 18604 56384 18644 57772
rect 18987 57763 19029 57772
rect 19084 57762 19124 57847
rect 18699 57644 18741 57653
rect 18699 57604 18700 57644
rect 18740 57604 18836 57644
rect 18699 57595 18741 57604
rect 18796 57602 18836 57604
rect 18796 57553 18836 57562
rect 18808 57476 19176 57485
rect 18848 57436 18890 57476
rect 18930 57436 18972 57476
rect 19012 57436 19054 57476
rect 19094 57436 19136 57476
rect 18808 57427 19176 57436
rect 19276 57065 19316 57856
rect 19468 57896 19508 57940
rect 19371 57140 19413 57149
rect 19371 57100 19372 57140
rect 19412 57100 19413 57140
rect 19371 57091 19413 57100
rect 19275 57056 19317 57065
rect 19275 57016 19276 57056
rect 19316 57016 19317 57056
rect 19275 57007 19317 57016
rect 19275 56888 19317 56897
rect 19275 56848 19276 56888
rect 19316 56848 19317 56888
rect 19275 56839 19317 56848
rect 18987 56552 19029 56561
rect 18987 56512 18988 56552
rect 19028 56512 19029 56552
rect 18987 56503 19029 56512
rect 18548 56344 18644 56384
rect 18988 56384 19028 56503
rect 18412 56300 18452 56309
rect 18316 56260 18412 56300
rect 18219 56048 18261 56057
rect 18219 56008 18220 56048
rect 18260 56008 18261 56048
rect 18219 55999 18261 56008
rect 17547 55628 17589 55637
rect 17547 55588 17548 55628
rect 17588 55588 17589 55628
rect 17547 55579 17589 55588
rect 17644 55553 17684 55638
rect 17643 55544 17685 55553
rect 17643 55504 17644 55544
rect 17684 55504 17685 55544
rect 17643 55495 17685 55504
rect 17740 55544 17780 55553
rect 17452 55420 17588 55460
rect 17548 55376 17588 55420
rect 17740 55376 17780 55504
rect 17548 55336 17780 55376
rect 17932 55376 17972 55385
rect 17451 54956 17493 54965
rect 17451 54916 17452 54956
rect 17492 54916 17493 54956
rect 17451 54907 17493 54916
rect 16876 54872 16916 54881
rect 16779 53696 16821 53705
rect 16779 53656 16780 53696
rect 16820 53656 16821 53696
rect 16779 53647 16821 53656
rect 16876 53528 16916 54832
rect 16972 54872 17012 54881
rect 17356 54872 17396 54881
rect 17012 54832 17356 54872
rect 16972 54823 17012 54832
rect 17356 54823 17396 54832
rect 17452 54872 17492 54907
rect 17452 54821 17492 54832
rect 17548 54872 17588 54883
rect 17548 54797 17588 54832
rect 17644 54872 17684 55336
rect 17835 55040 17877 55049
rect 17547 54788 17589 54797
rect 17547 54748 17548 54788
rect 17588 54748 17589 54788
rect 17547 54739 17589 54748
rect 17163 54620 17205 54629
rect 17644 54620 17684 54832
rect 17163 54580 17164 54620
rect 17204 54580 17300 54620
rect 17163 54571 17205 54580
rect 17260 54209 17300 54580
rect 17452 54580 17684 54620
rect 17740 55000 17836 55040
rect 17876 55000 17877 55040
rect 17259 54200 17301 54209
rect 17259 54160 17260 54200
rect 17300 54160 17301 54200
rect 17259 54151 17301 54160
rect 17260 54116 17300 54151
rect 17260 54066 17300 54076
rect 17164 54032 17204 54043
rect 17164 53957 17204 53992
rect 17163 53948 17205 53957
rect 17163 53908 17164 53948
rect 17204 53908 17205 53948
rect 17163 53899 17205 53908
rect 17452 53873 17492 54580
rect 17547 54200 17589 54209
rect 17547 54160 17548 54200
rect 17588 54160 17589 54200
rect 17547 54151 17589 54160
rect 17451 53864 17493 53873
rect 17451 53824 17452 53864
rect 17492 53824 17493 53864
rect 17451 53815 17493 53824
rect 17259 53696 17301 53705
rect 17259 53656 17260 53696
rect 17300 53656 17301 53696
rect 17259 53647 17301 53656
rect 16588 53488 16916 53528
rect 16971 53528 17013 53537
rect 16971 53488 16972 53528
rect 17012 53488 17013 53528
rect 16588 53033 16628 53488
rect 16971 53479 17013 53488
rect 17163 53528 17205 53537
rect 17163 53488 17164 53528
rect 17204 53488 17205 53528
rect 17163 53479 17205 53488
rect 16876 53360 16916 53369
rect 16684 53318 16724 53327
rect 16684 53117 16724 53278
rect 16780 53320 16876 53360
rect 16683 53108 16725 53117
rect 16683 53068 16684 53108
rect 16724 53068 16725 53108
rect 16683 53059 16725 53068
rect 16587 53024 16629 53033
rect 16587 52984 16588 53024
rect 16628 52984 16629 53024
rect 16587 52975 16629 52984
rect 16683 52940 16725 52949
rect 16683 52900 16684 52940
rect 16724 52900 16725 52940
rect 16683 52891 16725 52900
rect 16491 52688 16533 52697
rect 16491 52648 16492 52688
rect 16532 52648 16533 52688
rect 16491 52639 16533 52648
rect 16588 52604 16628 52615
rect 16492 52520 16532 52531
rect 16588 52529 16628 52564
rect 16492 52445 16532 52480
rect 16587 52520 16629 52529
rect 16587 52480 16588 52520
rect 16628 52480 16629 52520
rect 16587 52471 16629 52480
rect 16684 52520 16724 52891
rect 16684 52471 16724 52480
rect 16491 52436 16533 52445
rect 16491 52396 16492 52436
rect 16532 52396 16533 52436
rect 16491 52387 16533 52396
rect 16396 52144 16628 52184
rect 16299 52100 16341 52109
rect 16299 52060 16300 52100
rect 16340 52060 16341 52100
rect 16299 52051 16341 52060
rect 16395 52016 16437 52025
rect 16395 51976 16396 52016
rect 16436 51976 16437 52016
rect 16395 51967 16437 51976
rect 16204 51848 16244 51857
rect 16204 51689 16244 51808
rect 16300 51848 16340 51859
rect 16300 51773 16340 51808
rect 16299 51764 16341 51773
rect 16299 51724 16300 51764
rect 16340 51724 16341 51764
rect 16299 51715 16341 51724
rect 16396 51689 16436 51967
rect 16203 51680 16245 51689
rect 16203 51640 16204 51680
rect 16244 51640 16245 51680
rect 16203 51631 16245 51640
rect 16395 51680 16437 51689
rect 16395 51640 16396 51680
rect 16436 51640 16437 51680
rect 16395 51631 16437 51640
rect 16299 51596 16341 51605
rect 16299 51556 16300 51596
rect 16340 51556 16341 51596
rect 16299 51547 16341 51556
rect 16203 50336 16245 50345
rect 16203 50296 16204 50336
rect 16244 50296 16245 50336
rect 16203 50287 16245 50296
rect 16012 49624 16148 49664
rect 15724 49447 15764 49456
rect 16012 49496 16052 49505
rect 16012 49253 16052 49456
rect 15627 49244 15669 49253
rect 15627 49204 15628 49244
rect 15668 49204 15669 49244
rect 15627 49195 15669 49204
rect 16011 49244 16053 49253
rect 16011 49204 16012 49244
rect 16052 49204 16053 49244
rect 16011 49195 16053 49204
rect 15531 49160 15573 49169
rect 15531 49120 15532 49160
rect 15572 49120 15573 49160
rect 15531 49111 15573 49120
rect 15188 48868 15476 48908
rect 15148 48859 15188 48868
rect 15436 48824 15476 48868
rect 15436 48775 15476 48784
rect 15532 48824 15572 48833
rect 15052 48700 15188 48740
rect 14955 48691 14997 48700
rect 14956 47993 14996 48691
rect 15051 48488 15093 48497
rect 15051 48448 15052 48488
rect 15092 48448 15093 48488
rect 15051 48439 15093 48448
rect 14955 47984 14997 47993
rect 14955 47944 14956 47984
rect 14996 47944 14997 47984
rect 14955 47935 14997 47944
rect 14956 47312 14996 47321
rect 14956 47069 14996 47272
rect 14955 47060 14997 47069
rect 14955 47020 14956 47060
rect 14996 47020 14997 47060
rect 14955 47011 14997 47020
rect 15052 46892 15092 48439
rect 14764 45088 14900 45128
rect 14956 46852 15092 46892
rect 14667 44624 14709 44633
rect 14667 44584 14668 44624
rect 14708 44584 14709 44624
rect 14667 44575 14709 44584
rect 14667 44372 14709 44381
rect 14667 44332 14668 44372
rect 14708 44332 14709 44372
rect 14667 44323 14709 44332
rect 14668 44288 14708 44323
rect 14668 44237 14708 44248
rect 14667 43868 14709 43877
rect 14667 43828 14668 43868
rect 14708 43828 14709 43868
rect 14667 43819 14709 43828
rect 14668 43448 14708 43819
rect 14668 43399 14708 43408
rect 14668 42776 14708 42785
rect 14572 42736 14668 42776
rect 13996 42642 14036 42727
rect 14188 42524 14228 42533
rect 14228 42484 14420 42524
rect 14188 42475 14228 42484
rect 13516 42232 13652 42272
rect 13324 41936 13364 41945
rect 13227 41684 13269 41693
rect 13227 41644 13228 41684
rect 13268 41644 13269 41684
rect 13227 41635 13269 41644
rect 13228 41264 13268 41635
rect 13324 41525 13364 41896
rect 13323 41516 13365 41525
rect 13323 41476 13324 41516
rect 13364 41476 13365 41516
rect 13323 41467 13365 41476
rect 13515 41516 13557 41525
rect 13515 41476 13516 41516
rect 13556 41476 13557 41516
rect 13515 41467 13557 41476
rect 13419 41432 13461 41441
rect 13419 41392 13420 41432
rect 13460 41392 13461 41432
rect 13419 41383 13461 41392
rect 13420 41298 13460 41383
rect 13228 41215 13268 41224
rect 12939 39668 12981 39677
rect 12939 39628 12940 39668
rect 12980 39628 12981 39668
rect 12939 39619 12981 39628
rect 12940 39534 12980 39619
rect 12652 38704 12788 38744
rect 12652 36056 12692 38704
rect 13036 38669 13076 39712
rect 13516 39752 13556 41467
rect 13516 39703 13556 39712
rect 13419 38744 13461 38753
rect 13419 38704 13420 38744
rect 13460 38704 13461 38744
rect 13419 38695 13461 38704
rect 13035 38660 13077 38669
rect 13035 38620 13036 38660
rect 13076 38620 13077 38660
rect 13035 38611 13077 38620
rect 13323 38240 13365 38249
rect 13323 38200 13324 38240
rect 13364 38200 13365 38240
rect 13323 38191 13365 38200
rect 12748 38156 12788 38165
rect 12748 37829 12788 38116
rect 12843 38156 12885 38165
rect 12843 38116 12844 38156
rect 12884 38116 12885 38156
rect 12843 38107 12885 38116
rect 12844 38022 12884 38107
rect 13324 37913 13364 38191
rect 13420 38165 13460 38695
rect 13419 38156 13461 38165
rect 13419 38116 13420 38156
rect 13460 38116 13461 38156
rect 13419 38107 13461 38116
rect 13323 37904 13365 37913
rect 13323 37864 13324 37904
rect 13364 37864 13365 37904
rect 13323 37855 13365 37864
rect 12747 37820 12789 37829
rect 12747 37780 12748 37820
rect 12788 37780 12789 37820
rect 12747 37771 12789 37780
rect 12843 37316 12885 37325
rect 12843 37276 12844 37316
rect 12884 37276 12885 37316
rect 12843 37267 12885 37276
rect 12747 36728 12789 36737
rect 12747 36688 12748 36728
rect 12788 36688 12789 36728
rect 12747 36679 12789 36688
rect 12748 36594 12788 36679
rect 12844 36140 12884 37267
rect 13420 36989 13460 38107
rect 13515 37400 13557 37409
rect 13515 37360 13516 37400
rect 13556 37360 13557 37400
rect 13515 37351 13557 37360
rect 13516 37266 13556 37351
rect 13419 36980 13461 36989
rect 13419 36940 13420 36980
rect 13460 36940 13461 36980
rect 13419 36931 13461 36940
rect 12940 36812 12980 36821
rect 12980 36772 13268 36812
rect 12940 36763 12980 36772
rect 13228 36728 13268 36772
rect 13228 36679 13268 36688
rect 13324 36728 13364 36737
rect 13324 36569 13364 36688
rect 13323 36560 13365 36569
rect 13323 36520 13324 36560
rect 13364 36520 13365 36560
rect 13323 36511 13365 36520
rect 13227 36476 13269 36485
rect 13227 36436 13228 36476
rect 13268 36436 13269 36476
rect 13227 36427 13269 36436
rect 12844 36100 13076 36140
rect 12652 36016 12980 36056
rect 12556 35932 12788 35972
rect 12172 35839 12212 35848
rect 12460 35888 12500 35897
rect 11980 35754 12020 35839
rect 12076 35720 12116 35729
rect 12460 35720 12500 35848
rect 12652 35877 12692 35886
rect 12652 35729 12692 35837
rect 11787 35468 11829 35477
rect 11787 35428 11788 35468
rect 11828 35428 11829 35468
rect 11787 35419 11829 35428
rect 11788 35216 11828 35244
rect 11692 35176 11788 35216
rect 11692 34973 11732 35176
rect 11788 35167 11828 35176
rect 12076 35141 12116 35680
rect 12268 35680 12500 35720
rect 12556 35720 12596 35729
rect 12172 35225 12212 35310
rect 12171 35216 12213 35225
rect 12171 35176 12172 35216
rect 12212 35176 12213 35216
rect 12171 35167 12213 35176
rect 12075 35132 12117 35141
rect 12075 35092 12076 35132
rect 12116 35092 12117 35132
rect 12075 35083 12117 35092
rect 11691 34964 11733 34973
rect 11979 34964 12021 34973
rect 11691 34924 11692 34964
rect 11732 34924 11733 34964
rect 11691 34915 11733 34924
rect 11788 34924 11980 34964
rect 12020 34924 12021 34964
rect 11691 34544 11733 34553
rect 11691 34504 11692 34544
rect 11732 34504 11733 34544
rect 11691 34495 11733 34504
rect 11692 33620 11732 34495
rect 11788 34381 11828 34924
rect 11979 34915 12021 34924
rect 12172 34964 12212 34973
rect 11980 34830 12020 34915
rect 11979 34712 12021 34721
rect 11979 34672 11980 34712
rect 12020 34672 12021 34712
rect 11979 34663 12021 34672
rect 11788 33797 11828 34341
rect 11980 34292 12020 34663
rect 12172 34376 12212 34924
rect 12268 34721 12308 35680
rect 12459 35552 12501 35561
rect 12459 35512 12460 35552
rect 12500 35512 12501 35552
rect 12459 35503 12501 35512
rect 12364 35216 12404 35225
rect 12364 34973 12404 35176
rect 12460 35216 12500 35503
rect 12460 35167 12500 35176
rect 12363 34964 12405 34973
rect 12363 34924 12364 34964
rect 12404 34924 12405 34964
rect 12363 34915 12405 34924
rect 12267 34712 12309 34721
rect 12267 34672 12268 34712
rect 12308 34672 12309 34712
rect 12267 34663 12309 34672
rect 12172 34327 12212 34336
rect 12268 34376 12308 34385
rect 11980 34243 12020 34252
rect 12268 34049 12308 34336
rect 12460 34376 12500 34385
rect 12556 34376 12596 35680
rect 12651 35720 12693 35729
rect 12651 35680 12652 35720
rect 12692 35680 12693 35720
rect 12651 35671 12693 35680
rect 12651 35468 12693 35477
rect 12651 35428 12652 35468
rect 12692 35428 12693 35468
rect 12651 35419 12693 35428
rect 12500 34336 12596 34376
rect 12652 34376 12692 35419
rect 12748 34544 12788 35932
rect 12844 35888 12884 35897
rect 12844 35048 12884 35848
rect 12844 34973 12884 35008
rect 12843 34964 12885 34973
rect 12843 34924 12844 34964
rect 12884 34924 12885 34964
rect 12843 34915 12885 34924
rect 12748 34504 12884 34544
rect 12747 34376 12789 34385
rect 12652 34336 12748 34376
rect 12788 34336 12789 34376
rect 12460 34327 12500 34336
rect 12747 34327 12789 34336
rect 12748 34242 12788 34327
rect 12844 34292 12884 34504
rect 12940 34469 12980 36016
rect 12939 34460 12981 34469
rect 12939 34420 12940 34460
rect 12980 34420 12981 34460
rect 12939 34411 12981 34420
rect 12844 34252 12980 34292
rect 12363 34208 12405 34217
rect 12363 34168 12364 34208
rect 12404 34168 12405 34208
rect 12363 34159 12405 34168
rect 12364 34074 12404 34159
rect 12459 34124 12501 34133
rect 12459 34084 12460 34124
rect 12500 34084 12501 34124
rect 12459 34075 12501 34084
rect 12267 34040 12309 34049
rect 12267 34000 12268 34040
rect 12308 34000 12309 34040
rect 12267 33991 12309 34000
rect 11787 33788 11829 33797
rect 11787 33748 11788 33788
rect 11828 33748 11829 33788
rect 11787 33739 11829 33748
rect 12363 33788 12405 33797
rect 12363 33748 12364 33788
rect 12404 33748 12405 33788
rect 12363 33739 12405 33748
rect 12076 33704 12116 33713
rect 12116 33664 12212 33704
rect 12076 33655 12116 33664
rect 11692 33580 11924 33620
rect 11500 33328 11636 33368
rect 11403 32192 11445 32201
rect 11403 32152 11404 32192
rect 11444 32152 11445 32192
rect 11403 32143 11445 32152
rect 11212 29128 11308 29168
rect 11020 28960 11156 29000
rect 10731 28916 10773 28925
rect 10731 28876 10732 28916
rect 10772 28876 10773 28916
rect 10731 28867 10773 28876
rect 10732 27656 10772 28867
rect 10732 27607 10772 27616
rect 10636 26489 10676 27532
rect 10731 27488 10773 27497
rect 10731 27448 10732 27488
rect 10772 27448 10773 27488
rect 10731 27439 10773 27448
rect 10635 26480 10677 26489
rect 10635 26440 10636 26480
rect 10676 26440 10677 26480
rect 10635 26431 10677 26440
rect 10635 23960 10677 23969
rect 10635 23920 10636 23960
rect 10676 23920 10677 23960
rect 10635 23911 10677 23920
rect 10539 20096 10581 20105
rect 10539 20056 10540 20096
rect 10580 20056 10581 20096
rect 10539 20047 10581 20056
rect 10540 19853 10580 20047
rect 10636 20021 10676 23911
rect 10732 21617 10772 27439
rect 10827 25556 10869 25565
rect 10827 25516 10828 25556
rect 10868 25516 10869 25556
rect 10827 25507 10869 25516
rect 10731 21608 10773 21617
rect 10731 21568 10732 21608
rect 10772 21568 10773 21608
rect 10731 21559 10773 21568
rect 10731 20768 10773 20777
rect 10731 20728 10732 20768
rect 10772 20728 10773 20768
rect 10731 20719 10773 20728
rect 10828 20768 10868 25507
rect 11019 23792 11061 23801
rect 11019 23752 11020 23792
rect 11060 23752 11061 23792
rect 11019 23743 11061 23752
rect 11020 23658 11060 23743
rect 11019 23372 11061 23381
rect 11019 23332 11020 23372
rect 11060 23332 11061 23372
rect 11019 23323 11061 23332
rect 10924 22280 10964 22289
rect 10924 22121 10964 22240
rect 10923 22112 10965 22121
rect 10923 22072 10924 22112
rect 10964 22072 10965 22112
rect 10923 22063 10965 22072
rect 10923 21860 10965 21869
rect 10923 21820 10924 21860
rect 10964 21820 10965 21860
rect 10923 21811 10965 21820
rect 10924 21113 10964 21811
rect 11020 21608 11060 23323
rect 11116 23129 11156 28960
rect 11212 27656 11252 29128
rect 11308 29119 11348 29128
rect 11404 28580 11444 32143
rect 11500 28757 11540 33328
rect 11596 32869 11636 32878
rect 11596 32360 11636 32829
rect 11787 32780 11829 32789
rect 11787 32740 11788 32780
rect 11828 32740 11829 32780
rect 11787 32731 11829 32740
rect 11788 32646 11828 32731
rect 11596 32311 11636 32320
rect 11692 31352 11732 31361
rect 11692 30680 11732 31312
rect 11692 30521 11732 30640
rect 11691 30512 11733 30521
rect 11691 30472 11692 30512
rect 11732 30472 11733 30512
rect 11691 30463 11733 30472
rect 11595 29840 11637 29849
rect 11595 29800 11596 29840
rect 11636 29800 11637 29840
rect 11595 29791 11637 29800
rect 11596 29261 11636 29791
rect 11595 29252 11637 29261
rect 11595 29212 11596 29252
rect 11636 29212 11637 29252
rect 11595 29203 11637 29212
rect 11499 28748 11541 28757
rect 11499 28708 11500 28748
rect 11540 28708 11541 28748
rect 11499 28699 11541 28708
rect 11308 28540 11444 28580
rect 11308 28421 11348 28540
rect 11307 28412 11349 28421
rect 11307 28372 11308 28412
rect 11348 28372 11349 28412
rect 11307 28363 11349 28372
rect 11403 28328 11445 28337
rect 11403 28288 11404 28328
rect 11444 28288 11445 28328
rect 11403 28279 11445 28288
rect 11500 28328 11540 28337
rect 11596 28328 11636 29203
rect 11788 29154 11828 29163
rect 11692 28580 11732 28589
rect 11788 28580 11828 29114
rect 11884 28673 11924 33580
rect 12172 33293 12212 33664
rect 12268 33452 12308 33461
rect 12171 33284 12213 33293
rect 12171 33244 12172 33284
rect 12212 33244 12213 33284
rect 12171 33235 12213 33244
rect 11979 33116 12021 33125
rect 11979 33076 11980 33116
rect 12020 33076 12021 33116
rect 11979 33067 12021 33076
rect 11980 32864 12020 33067
rect 11980 32360 12020 32824
rect 11980 32311 12020 32320
rect 12268 31436 12308 33412
rect 12364 32192 12404 33739
rect 12460 33620 12500 34075
rect 12747 34040 12789 34049
rect 12747 34000 12748 34040
rect 12788 34000 12789 34040
rect 12747 33991 12789 34000
rect 12555 33956 12597 33965
rect 12555 33916 12556 33956
rect 12596 33916 12597 33956
rect 12555 33907 12597 33916
rect 12460 33571 12500 33580
rect 12460 32192 12500 32201
rect 12364 32152 12460 32192
rect 12460 32143 12500 32152
rect 12556 32192 12596 33907
rect 12652 33452 12692 33461
rect 12652 33209 12692 33412
rect 12651 33200 12693 33209
rect 12651 33160 12652 33200
rect 12692 33160 12693 33200
rect 12651 33151 12693 33160
rect 12651 32444 12693 32453
rect 12651 32404 12652 32444
rect 12692 32404 12693 32444
rect 12651 32395 12693 32404
rect 12556 32143 12596 32152
rect 12652 31613 12692 32395
rect 12748 32360 12788 33991
rect 12940 33797 12980 34252
rect 12939 33788 12981 33797
rect 12939 33748 12940 33788
rect 12980 33748 12981 33788
rect 13036 33788 13076 36100
rect 13132 35216 13172 35227
rect 13132 35141 13172 35176
rect 13131 35132 13173 35141
rect 13131 35092 13132 35132
rect 13172 35092 13173 35132
rect 13131 35083 13173 35092
rect 13228 34973 13268 36427
rect 13612 35057 13652 42232
rect 13804 41941 13844 41950
rect 13804 41441 13844 41901
rect 14380 41936 14420 42484
rect 14380 41887 14420 41896
rect 14476 41936 14516 41945
rect 14476 41777 14516 41896
rect 13996 41768 14036 41777
rect 13899 41684 13941 41693
rect 13899 41644 13900 41684
rect 13940 41644 13941 41684
rect 13899 41635 13941 41644
rect 13803 41432 13845 41441
rect 13803 41392 13804 41432
rect 13844 41392 13845 41432
rect 13803 41383 13845 41392
rect 13900 40424 13940 41635
rect 13900 38912 13940 40384
rect 13996 40349 14036 41728
rect 14475 41768 14517 41777
rect 14475 41728 14476 41768
rect 14516 41728 14517 41768
rect 14475 41719 14517 41728
rect 14476 41273 14516 41719
rect 14380 41264 14420 41273
rect 14092 41224 14380 41264
rect 14092 40676 14132 41224
rect 14380 41215 14420 41224
rect 14475 41264 14517 41273
rect 14475 41224 14476 41264
rect 14516 41224 14517 41264
rect 14475 41215 14517 41224
rect 14476 41130 14516 41215
rect 14092 40627 14132 40636
rect 14380 40424 14420 40433
rect 13995 40340 14037 40349
rect 13995 40300 13996 40340
rect 14036 40300 14037 40340
rect 13995 40291 14037 40300
rect 14380 40013 14420 40384
rect 14476 40424 14516 40433
rect 14476 40265 14516 40384
rect 14475 40256 14517 40265
rect 14475 40216 14476 40256
rect 14516 40216 14517 40256
rect 14475 40207 14517 40216
rect 14379 40004 14421 40013
rect 14379 39964 14380 40004
rect 14420 39964 14421 40004
rect 14379 39955 14421 39964
rect 14188 39836 14228 39845
rect 13996 39738 14036 39747
rect 13996 39089 14036 39698
rect 14188 39173 14228 39796
rect 14187 39164 14229 39173
rect 14187 39124 14188 39164
rect 14228 39124 14229 39164
rect 14187 39115 14229 39124
rect 13995 39080 14037 39089
rect 13995 39040 13996 39080
rect 14036 39040 14037 39080
rect 13995 39031 14037 39040
rect 14380 38912 14420 38921
rect 13940 38872 14036 38912
rect 13900 38863 13940 38872
rect 13899 38660 13941 38669
rect 13899 38620 13900 38660
rect 13940 38620 13941 38660
rect 13899 38611 13941 38620
rect 13804 38226 13844 38235
rect 13708 37652 13748 37661
rect 13804 37652 13844 38186
rect 13748 37612 13844 37652
rect 13708 37603 13748 37612
rect 13803 36980 13845 36989
rect 13803 36940 13804 36980
rect 13844 36940 13845 36980
rect 13803 36931 13845 36940
rect 13707 36644 13749 36653
rect 13707 36604 13708 36644
rect 13748 36604 13749 36644
rect 13707 36595 13749 36604
rect 13804 36644 13844 36931
rect 13708 36510 13748 36595
rect 13611 35048 13653 35057
rect 13611 35008 13612 35048
rect 13652 35008 13653 35048
rect 13611 34999 13653 35008
rect 13227 34964 13269 34973
rect 13227 34924 13228 34964
rect 13268 34924 13269 34964
rect 13227 34915 13269 34924
rect 13036 33748 13172 33788
rect 12939 33739 12981 33748
rect 12844 33662 12884 33671
rect 12843 33622 12844 33629
rect 12884 33622 12885 33629
rect 12843 33620 12885 33622
rect 12843 33580 12844 33620
rect 12884 33580 12885 33620
rect 12843 33571 12885 33580
rect 12748 32311 12788 32320
rect 12651 31604 12693 31613
rect 12651 31564 12652 31604
rect 12692 31564 12693 31604
rect 12651 31555 12693 31564
rect 12220 31396 12308 31436
rect 12220 31394 12260 31396
rect 12220 31345 12260 31354
rect 12363 31184 12405 31193
rect 12363 31144 12364 31184
rect 12404 31144 12405 31184
rect 12363 31135 12405 31144
rect 12364 31050 12404 31135
rect 12364 30764 12404 30773
rect 12404 30724 12596 30764
rect 12364 30715 12404 30724
rect 12220 30638 12260 30647
rect 12220 30596 12260 30598
rect 12220 30556 12500 30596
rect 11979 30092 12021 30101
rect 11979 30052 11980 30092
rect 12020 30052 12021 30092
rect 11979 30043 12021 30052
rect 12460 30092 12500 30556
rect 12460 30043 12500 30052
rect 11980 29336 12020 30043
rect 12171 29840 12213 29849
rect 12171 29800 12172 29840
rect 12212 29800 12213 29840
rect 12171 29791 12213 29800
rect 12268 29840 12308 29849
rect 11980 29287 12020 29296
rect 11979 28748 12021 28757
rect 11979 28708 11980 28748
rect 12020 28708 12021 28748
rect 11979 28699 12021 28708
rect 11883 28664 11925 28673
rect 11883 28624 11884 28664
rect 11924 28624 11925 28664
rect 11883 28615 11925 28624
rect 11732 28540 11828 28580
rect 11692 28531 11732 28540
rect 11540 28288 11636 28328
rect 11884 28328 11924 28337
rect 11500 28279 11540 28288
rect 11212 27497 11252 27616
rect 11211 27488 11253 27497
rect 11211 27448 11212 27488
rect 11252 27448 11253 27488
rect 11211 27439 11253 27448
rect 11308 26816 11348 26825
rect 11308 26153 11348 26776
rect 11307 26144 11349 26153
rect 11307 26104 11308 26144
rect 11348 26104 11349 26144
rect 11307 26095 11349 26104
rect 11404 25304 11444 28279
rect 11884 28169 11924 28288
rect 11883 28160 11925 28169
rect 11883 28120 11884 28160
rect 11924 28120 11925 28160
rect 11883 28111 11925 28120
rect 11980 27908 12020 28699
rect 12172 28580 12212 29791
rect 12268 29261 12308 29800
rect 12363 29588 12405 29597
rect 12363 29548 12364 29588
rect 12404 29548 12405 29588
rect 12363 29539 12405 29548
rect 12267 29252 12309 29261
rect 12267 29212 12268 29252
rect 12308 29212 12309 29252
rect 12267 29203 12309 29212
rect 12364 29000 12404 29539
rect 12556 29000 12596 30724
rect 12172 28531 12212 28540
rect 12268 28960 12404 29000
rect 12460 28960 12596 29000
rect 12748 29168 12788 29177
rect 12844 29168 12884 33571
rect 12939 32528 12981 32537
rect 12939 32488 12940 32528
rect 12980 32488 12981 32528
rect 12939 32479 12981 32488
rect 12788 29128 12884 29168
rect 12171 28328 12213 28337
rect 12171 28288 12172 28328
rect 12212 28288 12213 28328
rect 12171 28279 12213 28288
rect 12172 28194 12212 28279
rect 11788 27868 12020 27908
rect 11692 27642 11732 27651
rect 11692 27152 11732 27602
rect 11500 27112 11732 27152
rect 11500 27068 11540 27112
rect 11500 27019 11540 27028
rect 11788 26312 11828 27868
rect 11884 27740 11924 27749
rect 11924 27700 12020 27740
rect 11884 27691 11924 27700
rect 11788 26272 11924 26312
rect 11787 26144 11829 26153
rect 11787 26104 11788 26144
rect 11828 26104 11829 26144
rect 11787 26095 11829 26104
rect 11595 25892 11637 25901
rect 11595 25852 11596 25892
rect 11636 25852 11637 25892
rect 11595 25843 11637 25852
rect 11596 25556 11636 25843
rect 11596 25507 11636 25516
rect 11404 25220 11444 25264
rect 11212 25180 11444 25220
rect 11212 24632 11252 25180
rect 11404 25169 11444 25180
rect 11499 25220 11541 25229
rect 11499 25180 11500 25220
rect 11540 25180 11541 25220
rect 11499 25171 11541 25180
rect 11788 25220 11828 26095
rect 11788 25171 11828 25180
rect 11404 24800 11444 24809
rect 11500 24800 11540 25171
rect 11444 24760 11540 24800
rect 11404 24751 11444 24760
rect 11212 24473 11252 24592
rect 11596 24632 11636 24641
rect 11211 24464 11253 24473
rect 11211 24424 11212 24464
rect 11252 24424 11253 24464
rect 11211 24415 11253 24424
rect 11596 24389 11636 24592
rect 11595 24380 11637 24389
rect 11595 24340 11596 24380
rect 11636 24340 11637 24380
rect 11595 24331 11637 24340
rect 11691 24128 11733 24137
rect 11691 24088 11692 24128
rect 11732 24088 11737 24128
rect 11691 24079 11737 24088
rect 11212 23792 11252 23801
rect 11212 23297 11252 23752
rect 11307 23792 11349 23801
rect 11307 23752 11308 23792
rect 11348 23752 11349 23792
rect 11307 23743 11349 23752
rect 11500 23792 11540 23801
rect 11308 23658 11348 23743
rect 11500 23465 11540 23752
rect 11596 23792 11636 23801
rect 11596 23633 11636 23752
rect 11697 23792 11737 24079
rect 11737 23752 11828 23792
rect 11697 23743 11737 23752
rect 11595 23624 11637 23633
rect 11595 23584 11596 23624
rect 11636 23584 11637 23624
rect 11595 23575 11637 23584
rect 11692 23624 11732 23633
rect 11307 23456 11349 23465
rect 11307 23416 11308 23456
rect 11348 23416 11349 23456
rect 11307 23407 11349 23416
rect 11499 23456 11541 23465
rect 11499 23416 11500 23456
rect 11540 23416 11541 23456
rect 11499 23407 11541 23416
rect 11211 23288 11253 23297
rect 11211 23248 11212 23288
rect 11252 23248 11253 23288
rect 11211 23239 11253 23248
rect 11115 23120 11157 23129
rect 11115 23080 11116 23120
rect 11156 23080 11157 23120
rect 11115 23071 11157 23080
rect 11116 22986 11156 23071
rect 11115 21860 11157 21869
rect 11115 21820 11116 21860
rect 11156 21820 11157 21860
rect 11115 21811 11157 21820
rect 11020 21559 11060 21568
rect 11116 21608 11156 21811
rect 11308 21776 11348 23407
rect 11308 21727 11348 21736
rect 11404 23120 11444 23129
rect 11116 21559 11156 21568
rect 11404 21197 11444 23080
rect 11692 23045 11732 23584
rect 11691 23036 11733 23045
rect 11691 22996 11692 23036
rect 11732 22996 11733 23036
rect 11691 22987 11733 22996
rect 11403 21188 11445 21197
rect 11403 21148 11404 21188
rect 11444 21148 11445 21188
rect 11403 21139 11445 21148
rect 10923 21104 10965 21113
rect 10923 21064 10924 21104
rect 10964 21064 10965 21104
rect 10923 21055 10965 21064
rect 11019 20936 11061 20945
rect 11019 20896 11020 20936
rect 11060 20896 11061 20936
rect 11019 20887 11061 20896
rect 10868 20728 10964 20768
rect 10828 20719 10868 20728
rect 10635 20012 10677 20021
rect 10635 19972 10636 20012
rect 10676 19972 10677 20012
rect 10635 19963 10677 19972
rect 10732 19937 10772 20719
rect 10924 20105 10964 20728
rect 11020 20189 11060 20887
rect 11404 20861 11444 21139
rect 11595 20936 11637 20945
rect 11595 20896 11596 20936
rect 11636 20896 11637 20936
rect 11595 20887 11637 20896
rect 11788 20892 11828 23752
rect 11884 22793 11924 26272
rect 11980 25472 12020 27700
rect 12075 27656 12117 27665
rect 12075 27616 12076 27656
rect 12116 27616 12117 27656
rect 12075 27607 12117 27616
rect 12076 25985 12116 27607
rect 12171 27572 12213 27581
rect 12171 27532 12172 27572
rect 12212 27532 12213 27572
rect 12171 27523 12213 27532
rect 12075 25976 12117 25985
rect 12075 25936 12076 25976
rect 12116 25936 12117 25976
rect 12075 25927 12117 25936
rect 11980 25432 12116 25472
rect 11980 25309 12020 25318
rect 11980 24809 12020 25269
rect 11979 24800 12021 24809
rect 11979 24760 11980 24800
rect 12020 24760 12021 24800
rect 11979 24751 12021 24760
rect 12076 24725 12116 25432
rect 12075 24716 12117 24725
rect 12075 24676 12076 24716
rect 12116 24676 12117 24716
rect 12075 24667 12117 24676
rect 11883 22784 11925 22793
rect 11883 22744 11884 22784
rect 11924 22744 11925 22784
rect 11883 22735 11925 22744
rect 12172 22280 12212 27523
rect 12172 21449 12212 22240
rect 12171 21440 12213 21449
rect 12171 21400 12172 21440
rect 12212 21400 12213 21440
rect 12171 21391 12213 21400
rect 12075 21104 12117 21113
rect 12075 21064 12076 21104
rect 12116 21064 12117 21104
rect 12075 21055 12117 21064
rect 11403 20852 11445 20861
rect 11403 20812 11404 20852
rect 11444 20812 11445 20852
rect 11403 20803 11445 20812
rect 11212 20768 11252 20777
rect 11212 20357 11252 20728
rect 11308 20768 11348 20777
rect 11211 20348 11253 20357
rect 11211 20308 11212 20348
rect 11252 20308 11253 20348
rect 11211 20299 11253 20308
rect 11019 20180 11061 20189
rect 11019 20140 11020 20180
rect 11060 20140 11061 20180
rect 11019 20131 11061 20140
rect 11116 20180 11156 20189
rect 11308 20180 11348 20728
rect 11500 20768 11540 20777
rect 11404 20600 11444 20609
rect 11500 20600 11540 20728
rect 11596 20768 11636 20887
rect 11753 20783 11828 20892
rect 11979 20936 12021 20945
rect 11979 20896 11980 20936
rect 12020 20896 12021 20936
rect 11979 20887 12021 20896
rect 11596 20719 11636 20728
rect 11752 20728 11753 20777
rect 11793 20743 11828 20783
rect 11980 20768 12020 20887
rect 11793 20728 11794 20743
rect 11752 20719 11794 20728
rect 11980 20719 12020 20728
rect 12076 20768 12116 21055
rect 12268 20768 12308 28960
rect 12363 28160 12405 28169
rect 12363 28120 12364 28160
rect 12404 28120 12405 28160
rect 12363 28111 12405 28120
rect 12364 28026 12404 28111
rect 12363 27236 12405 27245
rect 12363 27196 12364 27236
rect 12404 27196 12405 27236
rect 12363 27187 12405 27196
rect 12364 26573 12404 27187
rect 12460 26993 12500 28960
rect 12555 28664 12597 28673
rect 12555 28624 12556 28664
rect 12596 28624 12597 28664
rect 12555 28615 12597 28624
rect 12556 28328 12596 28615
rect 12651 28580 12693 28589
rect 12651 28540 12652 28580
rect 12692 28540 12693 28580
rect 12651 28531 12693 28540
rect 12556 27581 12596 28288
rect 12555 27572 12597 27581
rect 12555 27532 12556 27572
rect 12596 27532 12597 27572
rect 12555 27523 12597 27532
rect 12555 27404 12597 27413
rect 12555 27364 12556 27404
rect 12596 27364 12597 27404
rect 12555 27355 12597 27364
rect 12459 26984 12501 26993
rect 12459 26944 12460 26984
rect 12500 26944 12501 26984
rect 12459 26935 12501 26944
rect 12363 26564 12405 26573
rect 12363 26524 12364 26564
rect 12404 26524 12405 26564
rect 12363 26515 12405 26524
rect 12364 25136 12404 26515
rect 12460 25892 12500 25901
rect 12460 25481 12500 25852
rect 12556 25565 12596 27355
rect 12652 27245 12692 28531
rect 12651 27236 12693 27245
rect 12651 27196 12652 27236
rect 12692 27196 12693 27236
rect 12651 27187 12693 27196
rect 12748 26741 12788 29128
rect 12940 28337 12980 32479
rect 13132 31688 13172 33748
rect 13228 33125 13268 34915
rect 13707 34460 13749 34469
rect 13707 34420 13708 34460
rect 13748 34420 13749 34460
rect 13707 34411 13749 34420
rect 13419 33284 13461 33293
rect 13419 33244 13420 33284
rect 13460 33244 13461 33284
rect 13419 33235 13461 33244
rect 13227 33116 13269 33125
rect 13227 33076 13228 33116
rect 13268 33076 13269 33116
rect 13227 33067 13269 33076
rect 13420 33041 13460 33235
rect 13419 33032 13461 33041
rect 13419 32992 13420 33032
rect 13460 32992 13461 33032
rect 13419 32983 13461 32992
rect 13611 33032 13653 33041
rect 13611 32992 13612 33032
rect 13652 32992 13653 33032
rect 13611 32983 13653 32992
rect 13227 32948 13269 32957
rect 13227 32908 13228 32948
rect 13268 32908 13269 32948
rect 13227 32899 13269 32908
rect 13515 32948 13557 32957
rect 13515 32908 13516 32948
rect 13556 32908 13557 32948
rect 13515 32899 13557 32908
rect 13612 32906 13652 32983
rect 13228 32864 13268 32899
rect 13228 32813 13268 32824
rect 13419 32696 13461 32705
rect 13419 32656 13420 32696
rect 13460 32656 13461 32696
rect 13419 32647 13461 32656
rect 13420 32562 13460 32647
rect 13516 32537 13556 32899
rect 13708 32869 13748 34411
rect 13804 33377 13844 36604
rect 13803 33368 13845 33377
rect 13803 33328 13804 33368
rect 13844 33328 13845 33368
rect 13803 33319 13845 33328
rect 13612 32857 13652 32866
rect 13703 32829 13748 32869
rect 13703 32780 13743 32829
rect 13703 32740 13748 32780
rect 13708 32612 13748 32740
rect 13708 32572 13844 32612
rect 13515 32528 13557 32537
rect 13515 32488 13516 32528
rect 13556 32488 13557 32528
rect 13515 32479 13557 32488
rect 13707 32444 13749 32453
rect 13707 32404 13708 32444
rect 13748 32404 13749 32444
rect 13707 32395 13749 32404
rect 13227 32360 13269 32369
rect 13227 32320 13228 32360
rect 13268 32320 13269 32360
rect 13227 32311 13269 32320
rect 13228 32192 13268 32311
rect 13228 32143 13268 32152
rect 13323 32192 13365 32201
rect 13323 32152 13324 32192
rect 13364 32152 13365 32192
rect 13323 32143 13365 32152
rect 13708 32192 13748 32395
rect 13708 32143 13748 32152
rect 13804 32192 13844 32572
rect 13324 32058 13364 32143
rect 13132 31648 13268 31688
rect 13131 31520 13173 31529
rect 13131 31480 13132 31520
rect 13172 31480 13173 31520
rect 13131 31471 13173 31480
rect 13132 31386 13172 31471
rect 13036 31184 13076 31193
rect 13036 28673 13076 31144
rect 13228 30680 13268 31648
rect 13419 31604 13461 31613
rect 13419 31564 13420 31604
rect 13460 31564 13461 31604
rect 13419 31555 13461 31564
rect 13323 31520 13365 31529
rect 13323 31480 13324 31520
rect 13364 31480 13365 31520
rect 13323 31471 13365 31480
rect 13324 31352 13364 31471
rect 13324 31303 13364 31312
rect 13324 30680 13364 30689
rect 13228 30640 13324 30680
rect 13228 29000 13268 30640
rect 13324 30631 13364 30640
rect 13228 28960 13364 29000
rect 13035 28664 13077 28673
rect 13035 28624 13036 28664
rect 13076 28624 13077 28664
rect 13035 28615 13077 28624
rect 13227 28664 13269 28673
rect 13227 28624 13228 28664
rect 13268 28624 13269 28664
rect 13227 28615 13269 28624
rect 12939 28328 12981 28337
rect 12939 28288 12940 28328
rect 12980 28288 12981 28328
rect 12939 28279 12981 28288
rect 12844 26816 12884 26825
rect 12747 26732 12789 26741
rect 12747 26692 12748 26732
rect 12788 26692 12789 26732
rect 12747 26683 12789 26692
rect 12844 26657 12884 26776
rect 12940 26816 12980 26825
rect 12843 26648 12885 26657
rect 12843 26608 12844 26648
rect 12884 26608 12885 26648
rect 12843 26599 12885 26608
rect 12651 26396 12693 26405
rect 12651 26356 12652 26396
rect 12692 26356 12693 26396
rect 12651 26347 12693 26356
rect 12555 25556 12597 25565
rect 12555 25516 12556 25556
rect 12596 25516 12597 25556
rect 12555 25507 12597 25516
rect 12459 25472 12501 25481
rect 12459 25432 12460 25472
rect 12500 25432 12501 25472
rect 12459 25423 12501 25432
rect 12460 25304 12500 25313
rect 12652 25304 12692 26347
rect 12748 26144 12788 26153
rect 12748 25733 12788 26104
rect 12843 26144 12885 26153
rect 12843 26104 12844 26144
rect 12884 26104 12885 26144
rect 12843 26095 12885 26104
rect 12844 26010 12884 26095
rect 12747 25724 12789 25733
rect 12747 25684 12748 25724
rect 12788 25684 12789 25724
rect 12747 25675 12789 25684
rect 12940 25649 12980 26776
rect 13132 26144 13172 26153
rect 13132 25901 13172 26104
rect 13131 25892 13173 25901
rect 13131 25852 13132 25892
rect 13172 25852 13173 25892
rect 13131 25843 13173 25852
rect 12939 25640 12981 25649
rect 12939 25600 12940 25640
rect 12980 25600 12981 25640
rect 12939 25591 12981 25600
rect 13035 25388 13077 25397
rect 13035 25348 13036 25388
rect 13076 25348 13077 25388
rect 13035 25339 13077 25348
rect 12940 25304 12980 25313
rect 12500 25264 12788 25304
rect 12460 25255 12500 25264
rect 12651 25136 12693 25145
rect 12364 25096 12500 25136
rect 12363 22448 12405 22457
rect 12363 22408 12364 22448
rect 12404 22408 12405 22448
rect 12363 22399 12405 22408
rect 12364 22314 12404 22399
rect 12268 20728 12404 20768
rect 12076 20719 12116 20728
rect 12268 20600 12308 20609
rect 11500 20560 12268 20600
rect 11404 20516 11444 20560
rect 12268 20551 12308 20560
rect 11404 20476 12212 20516
rect 11499 20348 11541 20357
rect 11499 20308 11500 20348
rect 11540 20308 11541 20348
rect 11499 20299 11541 20308
rect 11979 20348 12021 20357
rect 11979 20308 11980 20348
rect 12020 20308 12021 20348
rect 11979 20299 12021 20308
rect 11500 20264 11540 20299
rect 11500 20213 11540 20224
rect 11787 20264 11829 20273
rect 11787 20224 11788 20264
rect 11828 20224 11829 20264
rect 11787 20215 11829 20224
rect 11156 20140 11348 20180
rect 11116 20131 11156 20140
rect 10923 20096 10965 20105
rect 10923 20056 10924 20096
rect 10964 20056 10965 20096
rect 10923 20047 10965 20056
rect 11308 20096 11348 20140
rect 11308 20047 11348 20056
rect 11403 20096 11445 20105
rect 11403 20056 11404 20096
rect 11444 20056 11445 20096
rect 11403 20047 11445 20056
rect 11596 20096 11636 20105
rect 10924 19962 10964 20047
rect 11115 20012 11157 20021
rect 11115 19972 11116 20012
rect 11156 19972 11157 20012
rect 11115 19963 11157 19972
rect 10731 19928 10773 19937
rect 10731 19888 10732 19928
rect 10772 19888 10773 19928
rect 10731 19879 10773 19888
rect 10539 19844 10581 19853
rect 10539 19804 10540 19844
rect 10580 19804 10581 19844
rect 10539 19795 10581 19804
rect 10731 19676 10773 19685
rect 11116 19676 11156 19963
rect 11404 19962 11444 20047
rect 11499 19928 11541 19937
rect 11499 19888 11500 19928
rect 11540 19888 11541 19928
rect 11499 19879 11541 19888
rect 10731 19636 10732 19676
rect 10772 19636 10773 19676
rect 10731 19627 10773 19636
rect 11081 19636 11156 19676
rect 10443 19592 10485 19601
rect 10443 19552 10444 19592
rect 10484 19552 10485 19592
rect 10443 19543 10485 19552
rect 10252 19508 10292 19517
rect 10060 19468 10196 19508
rect 10060 19349 10100 19393
rect 9963 19340 10005 19349
rect 9963 19300 9964 19340
rect 10004 19300 10005 19340
rect 9963 19291 10005 19300
rect 10059 19340 10101 19349
rect 10059 19300 10060 19340
rect 10100 19300 10101 19340
rect 10059 19298 10101 19300
rect 10059 19291 10060 19298
rect 9964 18929 10004 19291
rect 10100 19291 10101 19298
rect 10060 19249 10100 19258
rect 10156 19172 10196 19468
rect 10292 19468 10395 19508
rect 10252 19459 10292 19468
rect 10355 19424 10395 19468
rect 10355 19384 10676 19424
rect 10540 19256 10580 19265
rect 10060 19132 10196 19172
rect 10444 19216 10540 19256
rect 9963 18920 10005 18929
rect 9963 18880 9964 18920
rect 10004 18880 10005 18920
rect 9963 18871 10005 18880
rect 9964 18584 10004 18871
rect 9964 18535 10004 18544
rect 9867 18500 9909 18509
rect 9867 18460 9868 18500
rect 9908 18460 9909 18500
rect 9867 18451 9909 18460
rect 9771 18416 9813 18425
rect 9771 18376 9772 18416
rect 9812 18376 9813 18416
rect 9771 18367 9813 18376
rect 9675 17744 9717 17753
rect 9675 17704 9676 17744
rect 9716 17704 9717 17744
rect 9675 17695 9717 17704
rect 9772 17744 9812 18367
rect 9676 17610 9716 17695
rect 9676 17081 9716 17166
rect 9675 17072 9717 17081
rect 9675 17032 9676 17072
rect 9716 17032 9717 17072
rect 9675 17023 9717 17032
rect 9772 16904 9812 17704
rect 9963 17744 10005 17753
rect 9963 17704 9964 17744
rect 10004 17704 10005 17744
rect 9963 17695 10005 17704
rect 9964 17576 10004 17695
rect 9964 17527 10004 17536
rect 9867 17072 9909 17081
rect 9867 17032 9868 17072
rect 9908 17032 9909 17072
rect 9867 17023 9909 17032
rect 9676 16864 9812 16904
rect 9579 16484 9621 16493
rect 9579 16444 9580 16484
rect 9620 16444 9621 16484
rect 9579 16435 9621 16444
rect 9580 16232 9620 16241
rect 9580 16073 9620 16192
rect 9579 16064 9621 16073
rect 9579 16024 9580 16064
rect 9620 16024 9621 16064
rect 9579 16015 9621 16024
rect 9580 15821 9620 16015
rect 9579 15812 9621 15821
rect 9579 15772 9580 15812
rect 9620 15772 9621 15812
rect 9579 15763 9621 15772
rect 9580 14897 9620 14982
rect 9579 14888 9621 14897
rect 9579 14848 9580 14888
rect 9620 14848 9621 14888
rect 9579 14839 9621 14848
rect 9579 14720 9621 14729
rect 9579 14680 9580 14720
rect 9620 14680 9621 14720
rect 9579 14671 9621 14680
rect 9580 14586 9620 14671
rect 9676 14552 9716 16864
rect 9771 16484 9813 16493
rect 9771 16444 9772 16484
rect 9812 16444 9813 16484
rect 9771 16435 9813 16444
rect 9772 15821 9812 16435
rect 9868 16073 9908 17023
rect 10060 16493 10100 19132
rect 10156 18668 10196 18679
rect 10156 18593 10196 18628
rect 10155 18584 10197 18593
rect 10155 18544 10156 18584
rect 10196 18544 10197 18584
rect 10155 18535 10197 18544
rect 10347 18584 10389 18593
rect 10347 18544 10348 18584
rect 10388 18544 10389 18584
rect 10347 18535 10389 18544
rect 10155 18164 10197 18173
rect 10155 18124 10156 18164
rect 10196 18124 10197 18164
rect 10155 18115 10197 18124
rect 10156 17744 10196 18115
rect 10156 17695 10196 17704
rect 10348 17744 10388 18535
rect 10444 17912 10484 19216
rect 10540 19207 10580 19216
rect 10636 19256 10676 19384
rect 10636 18752 10676 19216
rect 10732 19088 10772 19627
rect 11081 19271 11121 19636
rect 11211 19592 11253 19601
rect 11211 19552 11212 19592
rect 11252 19552 11253 19592
rect 11211 19543 11253 19552
rect 10732 19039 10772 19048
rect 10828 19256 10868 19265
rect 10828 18752 10868 19216
rect 10636 18712 10772 18752
rect 10539 18584 10581 18593
rect 10539 18544 10540 18584
rect 10580 18544 10581 18584
rect 10539 18535 10581 18544
rect 10636 18584 10676 18593
rect 10540 18450 10580 18535
rect 10636 18425 10676 18544
rect 10635 18416 10677 18425
rect 10635 18376 10636 18416
rect 10676 18376 10677 18416
rect 10635 18367 10677 18376
rect 10732 17996 10772 18712
rect 10828 18703 10868 18712
rect 10924 19256 10964 19265
rect 10924 18593 10964 19216
rect 11081 18920 11121 19231
rect 11212 18929 11252 19543
rect 11211 18920 11253 18929
rect 11081 18880 11156 18920
rect 10923 18584 10965 18593
rect 10923 18544 10924 18584
rect 10964 18544 10965 18584
rect 10923 18535 10965 18544
rect 10444 17863 10484 17872
rect 10540 17956 10772 17996
rect 10348 17695 10388 17704
rect 10444 17744 10484 17753
rect 10540 17744 10580 17956
rect 10827 17912 10869 17921
rect 10827 17872 10828 17912
rect 10868 17872 10869 17912
rect 10827 17863 10869 17872
rect 10484 17704 10580 17744
rect 10636 17744 10676 17755
rect 10444 17695 10484 17704
rect 10636 17669 10676 17704
rect 10732 17744 10772 17753
rect 10828 17744 10868 17863
rect 11019 17828 11061 17837
rect 11019 17788 11020 17828
rect 11060 17788 11061 17828
rect 11019 17779 11061 17788
rect 10772 17704 10868 17744
rect 10923 17744 10965 17753
rect 10923 17704 10924 17744
rect 10964 17704 10965 17744
rect 10732 17695 10772 17704
rect 10923 17695 10965 17704
rect 11020 17744 11060 17779
rect 11116 17753 11156 18880
rect 11211 18880 11212 18920
rect 11252 18880 11348 18920
rect 11211 18871 11253 18880
rect 11211 18752 11253 18761
rect 11211 18712 11212 18752
rect 11252 18712 11253 18752
rect 11211 18703 11253 18712
rect 11116 17744 11161 17753
rect 11116 17704 11121 17744
rect 10635 17660 10677 17669
rect 10635 17620 10636 17660
rect 10676 17620 10677 17660
rect 10635 17611 10677 17620
rect 10924 17610 10964 17695
rect 11020 17693 11060 17704
rect 11121 17695 11161 17704
rect 11116 17576 11156 17585
rect 10923 17492 10965 17501
rect 10923 17452 10924 17492
rect 10964 17452 10965 17492
rect 10923 17443 10965 17452
rect 10924 17072 10964 17443
rect 10964 17032 11060 17072
rect 10924 17023 10964 17032
rect 10923 16736 10965 16745
rect 10923 16696 10924 16736
rect 10964 16696 10965 16736
rect 10923 16687 10965 16696
rect 10059 16484 10101 16493
rect 10059 16444 10060 16484
rect 10100 16444 10101 16484
rect 10059 16435 10101 16444
rect 10731 16400 10773 16409
rect 10731 16360 10732 16400
rect 10772 16360 10773 16400
rect 10731 16351 10773 16360
rect 9867 16064 9909 16073
rect 9867 16024 9868 16064
rect 9908 16024 9909 16064
rect 9867 16015 9909 16024
rect 10155 15896 10197 15905
rect 10155 15856 10156 15896
rect 10196 15856 10197 15896
rect 10155 15847 10197 15856
rect 9771 15812 9813 15821
rect 9771 15772 9772 15812
rect 9812 15772 9813 15812
rect 9771 15763 9813 15772
rect 10059 15812 10101 15821
rect 10059 15772 10060 15812
rect 10100 15772 10101 15812
rect 10059 15763 10101 15772
rect 9963 14888 10005 14897
rect 9963 14848 9964 14888
rect 10004 14848 10005 14888
rect 10060 14888 10100 15763
rect 10156 15560 10196 15847
rect 10156 15511 10196 15520
rect 10539 15560 10581 15569
rect 10539 15520 10540 15560
rect 10580 15520 10581 15560
rect 10539 15511 10581 15520
rect 10732 15560 10772 16351
rect 10827 16232 10869 16241
rect 10827 16192 10828 16232
rect 10868 16192 10869 16232
rect 10827 16183 10869 16192
rect 10828 16098 10868 16183
rect 10732 15511 10772 15520
rect 10540 15426 10580 15511
rect 10348 15308 10388 15317
rect 10060 14848 10196 14888
rect 9963 14839 10005 14848
rect 9772 14720 9812 14729
rect 9964 14720 10004 14839
rect 10060 14720 10100 14729
rect 9812 14680 9908 14720
rect 9964 14680 10060 14720
rect 9772 14671 9812 14680
rect 9676 14512 9812 14552
rect 9484 14428 9716 14468
rect 9387 14216 9429 14225
rect 9387 14176 9388 14216
rect 9428 14176 9429 14216
rect 9387 14167 9429 14176
rect 9579 14132 9621 14141
rect 9579 14092 9580 14132
rect 9620 14092 9621 14132
rect 9579 14083 9621 14092
rect 9580 13208 9620 14083
rect 9676 14048 9716 14428
rect 9676 13999 9716 14008
rect 9772 13880 9812 14512
rect 9580 12293 9620 13168
rect 9676 13840 9812 13880
rect 9676 12620 9716 13840
rect 9771 13040 9813 13049
rect 9771 13000 9772 13040
rect 9812 13000 9813 13040
rect 9771 12991 9813 13000
rect 9772 12906 9812 12991
rect 9868 12965 9908 14680
rect 9963 14552 10005 14561
rect 9963 14512 9964 14552
rect 10004 14512 10005 14552
rect 9963 14503 10005 14512
rect 9964 14418 10004 14503
rect 9963 14048 10005 14057
rect 9963 14008 9964 14048
rect 10004 14008 10005 14048
rect 9963 13999 10005 14008
rect 9964 13914 10004 13999
rect 9963 13544 10005 13553
rect 9963 13504 9964 13544
rect 10004 13504 10005 13544
rect 9963 13495 10005 13504
rect 9964 13208 10004 13495
rect 9867 12956 9909 12965
rect 9867 12916 9868 12956
rect 9908 12916 9909 12956
rect 9867 12907 9909 12916
rect 9964 12797 10004 13168
rect 9963 12788 10005 12797
rect 9963 12748 9964 12788
rect 10004 12748 10005 12788
rect 9963 12739 10005 12748
rect 9676 12580 10004 12620
rect 9579 12284 9621 12293
rect 9579 12244 9580 12284
rect 9620 12244 9621 12284
rect 9579 12235 9621 12244
rect 9580 11537 9620 12235
rect 9579 11528 9621 11537
rect 9579 11488 9580 11528
rect 9620 11488 9621 11528
rect 9579 11479 9621 11488
rect 9868 11528 9908 11537
rect 9868 11360 9908 11488
rect 9676 11320 9908 11360
rect 9291 11276 9333 11285
rect 9291 11236 9292 11276
rect 9332 11236 9333 11276
rect 9291 11227 9333 11236
rect 9387 11108 9429 11117
rect 9387 11068 9388 11108
rect 9428 11068 9429 11108
rect 9387 11059 9429 11068
rect 9196 10975 9236 10984
rect 9388 11024 9428 11059
rect 9388 10973 9428 10984
rect 9579 11024 9621 11033
rect 9579 10984 9580 11024
rect 9620 10984 9621 11024
rect 9579 10975 9621 10984
rect 9580 10890 9620 10975
rect 9292 10772 9332 10781
rect 9332 10732 9524 10772
rect 9292 10723 9332 10732
rect 9004 10480 9140 10520
rect 9100 10352 9140 10480
rect 9196 10352 9236 10361
rect 9100 10312 9196 10352
rect 9003 10268 9045 10277
rect 9003 10228 9004 10268
rect 9044 10228 9045 10268
rect 9003 10219 9045 10228
rect 9004 10100 9044 10219
rect 9004 10051 9044 10060
rect 9003 9848 9045 9857
rect 9003 9808 9004 9848
rect 9044 9808 9045 9848
rect 9003 9799 9045 9808
rect 8907 8504 8949 8513
rect 8907 8464 8908 8504
rect 8948 8464 8949 8504
rect 8907 8455 8949 8464
rect 8811 8336 8853 8345
rect 8811 8296 8812 8336
rect 8852 8296 8853 8336
rect 8811 8287 8853 8296
rect 8660 8128 8756 8168
rect 8620 8119 8660 8128
rect 8907 8000 8949 8009
rect 8907 7960 8908 8000
rect 8948 7960 8949 8000
rect 8907 7951 8949 7960
rect 8908 7866 8948 7951
rect 8715 7748 8757 7757
rect 8715 7708 8716 7748
rect 8756 7708 8757 7748
rect 8715 7699 8757 7708
rect 8716 7160 8756 7699
rect 8811 7580 8853 7589
rect 8811 7540 8812 7580
rect 8852 7540 8853 7580
rect 8811 7531 8853 7540
rect 8716 4817 8756 7120
rect 8812 7244 8852 7531
rect 8715 4808 8757 4817
rect 8715 4768 8716 4808
rect 8756 4768 8757 4808
rect 8715 4759 8757 4768
rect 8332 2500 8468 2540
rect 8524 2500 8660 2540
rect 7083 2036 7125 2045
rect 7083 1996 7084 2036
rect 7124 1996 7125 2036
rect 7083 1987 7125 1996
rect 6699 1868 6741 1877
rect 6699 1828 6700 1868
rect 6740 1828 6741 1868
rect 6699 1819 6741 1828
rect 7084 1868 7124 1877
rect 6700 1734 6740 1819
rect 7084 1373 7124 1828
rect 7083 1364 7125 1373
rect 7083 1324 7084 1364
rect 7124 1324 7125 1364
rect 7083 1315 7125 1324
rect 6507 1280 6549 1289
rect 6507 1240 6508 1280
rect 6548 1240 6549 1280
rect 6507 1231 6549 1240
rect 6795 1280 6837 1289
rect 6795 1240 6796 1280
rect 6836 1240 6837 1280
rect 6795 1231 6837 1240
rect 6508 1146 6548 1231
rect 6699 1196 6741 1205
rect 6699 1156 6700 1196
rect 6740 1156 6741 1196
rect 6699 1147 6741 1156
rect 6603 1112 6645 1121
rect 6603 1072 6604 1112
rect 6644 1072 6645 1112
rect 6603 1063 6645 1072
rect 6411 944 6453 953
rect 6411 904 6412 944
rect 6452 904 6453 944
rect 6411 895 6453 904
rect 6411 440 6453 449
rect 6411 400 6412 440
rect 6452 400 6453 440
rect 6411 391 6453 400
rect 6219 188 6261 197
rect 6219 148 6220 188
rect 6260 148 6261 188
rect 6219 139 6261 148
rect 6220 80 6260 139
rect 6412 80 6452 391
rect 6604 80 6644 1063
rect 6700 1062 6740 1147
rect 6796 80 6836 1231
rect 6892 1196 6932 1205
rect 7180 1196 7220 2500
rect 7659 2372 7701 2381
rect 7659 2332 7660 2372
rect 7700 2332 7701 2372
rect 7659 2323 7701 2332
rect 7275 2120 7317 2129
rect 7275 2080 7276 2120
rect 7316 2080 7317 2120
rect 7275 2071 7317 2080
rect 7660 2120 7700 2323
rect 7660 2071 7700 2080
rect 7276 1986 7316 2071
rect 7755 2036 7797 2045
rect 7755 1996 7756 2036
rect 7796 1996 7797 2036
rect 7755 1987 7797 1996
rect 7468 1868 7508 1877
rect 7275 1532 7317 1541
rect 7275 1492 7276 1532
rect 7316 1492 7317 1532
rect 7275 1483 7317 1492
rect 6932 1156 7220 1196
rect 6892 1147 6932 1156
rect 7084 944 7124 953
rect 7084 533 7124 904
rect 7276 776 7316 1483
rect 7468 1289 7508 1828
rect 7563 1448 7605 1457
rect 7563 1408 7564 1448
rect 7604 1408 7605 1448
rect 7563 1399 7605 1408
rect 7467 1280 7509 1289
rect 7467 1240 7468 1280
rect 7508 1240 7509 1280
rect 7467 1231 7509 1240
rect 7371 1196 7413 1205
rect 7371 1156 7372 1196
rect 7412 1156 7413 1196
rect 7371 1147 7413 1156
rect 7180 736 7316 776
rect 7083 524 7125 533
rect 7083 484 7084 524
rect 7124 484 7125 524
rect 7083 475 7125 484
rect 6987 104 7029 113
rect 6987 80 6988 104
rect 3380 64 3400 80
rect 3320 0 3400 64
rect 3512 0 3592 80
rect 3704 0 3784 80
rect 3896 0 3976 80
rect 4088 0 4168 80
rect 4280 0 4360 80
rect 4472 0 4552 80
rect 4664 0 4744 80
rect 4856 0 4936 80
rect 5048 0 5128 80
rect 5240 0 5320 80
rect 5432 0 5512 80
rect 5624 0 5704 80
rect 5816 0 5896 80
rect 6008 0 6088 80
rect 6200 0 6280 80
rect 6392 0 6472 80
rect 6584 0 6664 80
rect 6776 0 6856 80
rect 6968 64 6988 80
rect 7028 80 7029 104
rect 7180 80 7220 736
rect 7372 80 7412 1147
rect 7564 80 7604 1399
rect 7756 80 7796 1987
rect 7852 1868 7892 1877
rect 7852 953 7892 1828
rect 7947 1868 7989 1877
rect 7947 1828 7948 1868
rect 7988 1828 7989 1868
rect 7947 1819 7989 1828
rect 8139 1868 8181 1877
rect 8139 1828 8140 1868
rect 8180 1828 8181 1868
rect 8139 1819 8181 1828
rect 7851 944 7893 953
rect 7851 904 7852 944
rect 7892 904 7893 944
rect 7851 895 7893 904
rect 7948 80 7988 1819
rect 8140 1734 8180 1819
rect 8331 1700 8373 1709
rect 8331 1660 8332 1700
rect 8372 1660 8373 1700
rect 8331 1651 8373 1660
rect 8332 1566 8372 1651
rect 8428 1541 8468 2500
rect 8620 1868 8660 2500
rect 8812 2213 8852 7204
rect 8811 2204 8853 2213
rect 8811 2164 8812 2204
rect 8852 2164 8853 2204
rect 8811 2155 8853 2164
rect 9004 2045 9044 9799
rect 9196 9680 9236 10312
rect 9484 10184 9524 10732
rect 9484 10135 9524 10144
rect 9580 10184 9620 10193
rect 9676 10184 9716 11320
rect 9771 10268 9813 10277
rect 9771 10228 9772 10268
rect 9812 10228 9813 10268
rect 9771 10219 9813 10228
rect 9620 10144 9716 10184
rect 9772 10184 9812 10219
rect 9580 10135 9620 10144
rect 9772 10133 9812 10144
rect 9771 10016 9813 10025
rect 9771 9976 9772 10016
rect 9812 9976 9813 10016
rect 9771 9967 9813 9976
rect 9772 9882 9812 9967
rect 9196 9631 9236 9640
rect 9964 9521 10004 12580
rect 10060 12536 10100 14680
rect 10156 14057 10196 14848
rect 10348 14720 10388 15268
rect 10636 15308 10676 15317
rect 10348 14671 10388 14680
rect 10444 14720 10484 14729
rect 10155 14048 10197 14057
rect 10155 14008 10156 14048
rect 10196 14008 10197 14048
rect 10155 13999 10197 14008
rect 10347 12956 10389 12965
rect 10347 12916 10348 12956
rect 10388 12916 10389 12956
rect 10347 12907 10389 12916
rect 10252 12536 10292 12545
rect 10060 12496 10252 12536
rect 10252 12487 10292 12496
rect 10348 12536 10388 12907
rect 10348 12487 10388 12496
rect 10444 12368 10484 14680
rect 10636 13217 10676 15268
rect 10924 14888 10964 16687
rect 10732 14848 10964 14888
rect 10635 13208 10677 13217
rect 10635 13168 10636 13208
rect 10676 13168 10677 13208
rect 10635 13159 10677 13168
rect 10540 12704 10580 12713
rect 10540 12620 10580 12664
rect 10635 12620 10677 12629
rect 10540 12580 10636 12620
rect 10676 12580 10677 12620
rect 10635 12571 10677 12580
rect 10252 12328 10484 12368
rect 10059 12032 10101 12041
rect 10059 11992 10060 12032
rect 10100 11992 10101 12032
rect 10059 11983 10101 11992
rect 10060 11696 10100 11983
rect 10060 11647 10100 11656
rect 10156 11696 10196 11705
rect 10059 11528 10101 11537
rect 10059 11488 10060 11528
rect 10100 11488 10101 11528
rect 10059 11479 10101 11488
rect 9676 9512 9716 9521
rect 9676 9353 9716 9472
rect 9963 9512 10005 9521
rect 9963 9472 9964 9512
rect 10004 9472 10005 9512
rect 9963 9463 10005 9472
rect 9675 9344 9717 9353
rect 9675 9304 9676 9344
rect 9716 9304 9717 9344
rect 9675 9295 9717 9304
rect 9387 8840 9429 8849
rect 9387 8800 9388 8840
rect 9428 8800 9429 8840
rect 9387 8791 9429 8800
rect 9291 8756 9333 8765
rect 9291 8716 9292 8756
rect 9332 8716 9333 8756
rect 9291 8707 9333 8716
rect 9196 8672 9236 8681
rect 9196 8429 9236 8632
rect 9292 8622 9332 8707
rect 9291 8504 9333 8513
rect 9291 8464 9292 8504
rect 9332 8464 9333 8504
rect 9291 8455 9333 8464
rect 9195 8420 9237 8429
rect 9195 8380 9196 8420
rect 9236 8380 9237 8420
rect 9195 8371 9237 8380
rect 9196 6992 9236 8371
rect 9292 7160 9332 8455
rect 9292 7111 9332 7120
rect 9196 6952 9332 6992
rect 9292 4481 9332 6952
rect 9291 4472 9333 4481
rect 9291 4432 9292 4472
rect 9332 4432 9333 4472
rect 9291 4423 9333 4432
rect 9388 4304 9428 8791
rect 9579 8756 9621 8765
rect 9579 8716 9580 8756
rect 9620 8716 9621 8756
rect 9579 8707 9621 8716
rect 9483 8336 9525 8345
rect 9483 8296 9484 8336
rect 9524 8296 9525 8336
rect 9483 8287 9525 8296
rect 9100 4264 9428 4304
rect 9003 2036 9045 2045
rect 9003 1996 9004 2036
rect 9044 1996 9045 2036
rect 9003 1987 9045 1996
rect 8620 1819 8660 1828
rect 9004 1868 9044 1877
rect 9100 1868 9140 4264
rect 9484 2540 9524 8287
rect 9580 6320 9620 8707
rect 9772 8672 9812 8681
rect 9964 8672 10004 9463
rect 9812 8632 10004 8672
rect 9772 8623 9812 8632
rect 10060 8000 10100 11479
rect 10156 11117 10196 11656
rect 10252 11201 10292 12328
rect 10732 12200 10772 14848
rect 10828 14720 10868 14731
rect 10828 14645 10868 14680
rect 10923 14720 10965 14729
rect 10923 14680 10924 14720
rect 10964 14680 10965 14720
rect 10923 14671 10965 14680
rect 10827 14636 10869 14645
rect 10827 14596 10828 14636
rect 10868 14596 10869 14636
rect 10827 14587 10869 14596
rect 10924 14586 10964 14671
rect 10827 13040 10869 13049
rect 10827 13000 10828 13040
rect 10868 13000 10869 13040
rect 10827 12991 10869 13000
rect 10828 12536 10868 12991
rect 10828 12487 10868 12496
rect 10924 12536 10964 12545
rect 10540 12160 10772 12200
rect 10348 11696 10388 11705
rect 10251 11192 10293 11201
rect 10251 11152 10252 11192
rect 10292 11152 10293 11192
rect 10251 11143 10293 11152
rect 10155 11108 10197 11117
rect 10155 11068 10156 11108
rect 10196 11068 10197 11108
rect 10155 11059 10197 11068
rect 10156 10184 10196 11059
rect 10252 10445 10292 11143
rect 10251 10436 10293 10445
rect 10251 10396 10252 10436
rect 10292 10396 10293 10436
rect 10251 10387 10293 10396
rect 10156 10135 10196 10144
rect 10348 10109 10388 11656
rect 10540 11360 10580 12160
rect 10636 11957 10676 12042
rect 10635 11948 10677 11957
rect 10635 11908 10636 11948
rect 10676 11908 10677 11948
rect 10635 11899 10677 11908
rect 10636 11696 10676 11705
rect 10827 11696 10869 11705
rect 10676 11656 10772 11696
rect 10636 11647 10676 11656
rect 10540 11320 10676 11360
rect 10539 10604 10581 10613
rect 10539 10564 10540 10604
rect 10580 10564 10581 10604
rect 10539 10555 10581 10564
rect 10443 10268 10485 10277
rect 10443 10228 10444 10268
rect 10484 10228 10485 10268
rect 10443 10219 10485 10228
rect 10444 10184 10484 10219
rect 10444 10133 10484 10144
rect 10540 10184 10580 10555
rect 10540 10135 10580 10144
rect 10347 10100 10389 10109
rect 10347 10060 10348 10100
rect 10388 10060 10389 10100
rect 10347 10051 10389 10060
rect 10300 8681 10340 8690
rect 10340 8641 10388 8672
rect 10300 8632 10388 8641
rect 10348 8168 10388 8632
rect 10348 8119 10388 8128
rect 10444 8504 10484 8513
rect 10156 8000 10196 8009
rect 10060 7960 10156 8000
rect 9963 7916 10005 7925
rect 9963 7876 9964 7916
rect 10004 7876 10100 7916
rect 9963 7867 10005 7876
rect 9675 7496 9717 7505
rect 9675 7456 9676 7496
rect 9716 7456 9717 7496
rect 9675 7447 9717 7456
rect 9676 6488 9716 7447
rect 9820 7169 9860 7178
rect 9860 7129 9908 7160
rect 9820 7120 9908 7129
rect 9868 6656 9908 7120
rect 9964 7001 10004 7086
rect 9963 6992 10005 7001
rect 9963 6952 9964 6992
rect 10004 6952 10005 6992
rect 9963 6943 10005 6952
rect 9963 6824 10005 6833
rect 9963 6784 9964 6824
rect 10004 6784 10005 6824
rect 9963 6775 10005 6784
rect 9868 6607 9908 6616
rect 9676 6439 9716 6448
rect 9580 6280 9716 6320
rect 9388 2500 9524 2540
rect 9579 2540 9621 2549
rect 9579 2500 9580 2540
rect 9620 2500 9621 2540
rect 9388 2045 9428 2500
rect 9579 2491 9621 2500
rect 9387 2036 9429 2045
rect 9387 1996 9388 2036
rect 9428 1996 9429 2036
rect 9387 1987 9429 1996
rect 9580 1868 9620 2491
rect 9676 1961 9716 6280
rect 9771 4136 9813 4145
rect 9771 4096 9772 4136
rect 9812 4096 9813 4136
rect 9771 4087 9813 4096
rect 9675 1952 9717 1961
rect 9675 1912 9676 1952
rect 9716 1912 9717 1952
rect 9675 1903 9717 1912
rect 9044 1828 9140 1868
rect 9292 1828 9524 1868
rect 9004 1819 9044 1828
rect 9196 1784 9236 1793
rect 9292 1784 9332 1828
rect 9236 1744 9332 1784
rect 9196 1735 9236 1744
rect 8812 1700 8852 1709
rect 8427 1532 8469 1541
rect 8427 1492 8428 1532
rect 8468 1492 8469 1532
rect 8427 1483 8469 1492
rect 8139 1364 8181 1373
rect 8139 1324 8140 1364
rect 8180 1324 8181 1364
rect 8139 1315 8181 1324
rect 8140 80 8180 1315
rect 8331 1280 8373 1289
rect 8331 1240 8332 1280
rect 8372 1240 8373 1280
rect 8331 1231 8373 1240
rect 8235 1112 8277 1121
rect 8235 1072 8236 1112
rect 8276 1072 8277 1112
rect 8235 1063 8277 1072
rect 8236 785 8276 1063
rect 8235 776 8277 785
rect 8235 736 8236 776
rect 8276 736 8277 776
rect 8235 727 8277 736
rect 8332 80 8372 1231
rect 8523 944 8565 953
rect 8523 904 8524 944
rect 8564 904 8565 944
rect 8523 895 8565 904
rect 8715 944 8757 953
rect 8715 904 8716 944
rect 8756 904 8757 944
rect 8715 895 8757 904
rect 8524 80 8564 895
rect 8716 80 8756 895
rect 8812 785 8852 1660
rect 8907 1700 8949 1709
rect 9388 1700 9428 1709
rect 8907 1660 8908 1700
rect 8948 1660 8949 1700
rect 8907 1651 8949 1660
rect 9292 1660 9388 1700
rect 8811 776 8853 785
rect 8811 736 8812 776
rect 8852 736 8853 776
rect 8811 727 8853 736
rect 8908 80 8948 1651
rect 9195 944 9237 953
rect 9195 904 9196 944
rect 9236 904 9237 944
rect 9195 895 9237 904
rect 9196 810 9236 895
rect 9099 524 9141 533
rect 9099 484 9100 524
rect 9140 484 9141 524
rect 9099 475 9141 484
rect 9100 80 9140 475
rect 9292 80 9332 1660
rect 9388 1651 9428 1660
rect 9387 1196 9429 1205
rect 9387 1156 9388 1196
rect 9428 1156 9429 1196
rect 9387 1147 9429 1156
rect 9388 1062 9428 1147
rect 9484 860 9524 1828
rect 9580 1819 9620 1828
rect 9772 1868 9812 4087
rect 9964 2540 10004 6775
rect 9772 1819 9812 1828
rect 9868 2500 10004 2540
rect 10060 2540 10100 7876
rect 10156 7505 10196 7960
rect 10155 7496 10197 7505
rect 10155 7456 10156 7496
rect 10196 7456 10197 7496
rect 10155 7447 10197 7456
rect 10155 6992 10197 7001
rect 10155 6952 10156 6992
rect 10196 6952 10197 6992
rect 10155 6943 10197 6952
rect 10156 6404 10196 6943
rect 10156 6355 10196 6364
rect 10251 6320 10293 6329
rect 10251 6280 10252 6320
rect 10292 6280 10293 6320
rect 10251 6271 10293 6280
rect 10060 2500 10196 2540
rect 9771 1700 9813 1709
rect 9771 1660 9772 1700
rect 9812 1660 9813 1700
rect 9771 1651 9813 1660
rect 9484 820 9716 860
rect 9483 692 9525 701
rect 9483 652 9484 692
rect 9524 652 9525 692
rect 9483 643 9525 652
rect 9484 80 9524 643
rect 9676 80 9716 820
rect 9772 281 9812 1651
rect 9868 1205 9908 2500
rect 10156 1881 10196 2500
rect 10156 1832 10196 1841
rect 10252 1784 10292 6271
rect 10348 6236 10388 6245
rect 10348 2540 10388 6196
rect 10444 4145 10484 8464
rect 10443 4136 10485 4145
rect 10443 4096 10444 4136
rect 10484 4096 10485 4136
rect 10443 4087 10485 4096
rect 10636 2540 10676 11320
rect 10732 10184 10772 11656
rect 10827 11656 10828 11696
rect 10868 11656 10869 11696
rect 10827 11647 10869 11656
rect 10828 11562 10868 11647
rect 10827 11192 10869 11201
rect 10827 11152 10828 11192
rect 10868 11152 10869 11192
rect 10827 11143 10869 11152
rect 10828 11024 10868 11143
rect 10924 11033 10964 12496
rect 11020 11705 11060 17032
rect 11116 16325 11156 17536
rect 11212 16661 11252 18703
rect 11308 18416 11348 18880
rect 11404 18584 11444 18593
rect 11500 18584 11540 19879
rect 11596 19517 11636 20056
rect 11788 20096 11828 20215
rect 11828 20056 11924 20096
rect 11788 20016 11828 20056
rect 11595 19508 11637 19517
rect 11595 19468 11596 19508
rect 11636 19468 11637 19508
rect 11595 19459 11637 19468
rect 11691 19424 11733 19433
rect 11691 19384 11692 19424
rect 11732 19384 11733 19424
rect 11691 19375 11733 19384
rect 11444 18544 11540 18584
rect 11404 18535 11444 18544
rect 11308 18376 11444 18416
rect 11404 17744 11444 18376
rect 11404 17695 11444 17704
rect 11308 17072 11348 17081
rect 11500 17072 11540 18544
rect 11692 19256 11732 19375
rect 11692 17669 11732 19216
rect 11691 17660 11733 17669
rect 11691 17620 11692 17660
rect 11732 17620 11733 17660
rect 11691 17611 11733 17620
rect 11884 17249 11924 20056
rect 11883 17240 11925 17249
rect 11883 17200 11884 17240
rect 11924 17200 11925 17240
rect 11883 17191 11925 17200
rect 11500 17032 11732 17072
rect 11211 16652 11253 16661
rect 11211 16612 11212 16652
rect 11252 16612 11253 16652
rect 11211 16603 11253 16612
rect 11212 16409 11252 16603
rect 11308 16577 11348 17032
rect 11307 16568 11349 16577
rect 11307 16528 11308 16568
rect 11348 16528 11349 16568
rect 11307 16519 11349 16528
rect 11211 16400 11253 16409
rect 11211 16360 11212 16400
rect 11252 16360 11253 16400
rect 11211 16351 11253 16360
rect 11115 16316 11157 16325
rect 11115 16276 11116 16316
rect 11156 16276 11157 16316
rect 11115 16267 11157 16276
rect 11211 15896 11253 15905
rect 11211 15856 11212 15896
rect 11252 15856 11253 15896
rect 11211 15847 11253 15856
rect 11115 14636 11157 14645
rect 11115 14596 11116 14636
rect 11156 14596 11157 14636
rect 11115 14587 11157 14596
rect 11019 11696 11061 11705
rect 11019 11656 11020 11696
rect 11060 11656 11061 11696
rect 11019 11647 11061 11656
rect 11019 11108 11061 11117
rect 11019 11068 11020 11108
rect 11060 11068 11061 11108
rect 11019 11059 11061 11068
rect 10828 10975 10868 10984
rect 10923 11024 10965 11033
rect 10923 10984 10924 11024
rect 10964 10984 10965 11024
rect 10923 10975 10965 10984
rect 11020 10974 11060 11059
rect 11116 10520 11156 14587
rect 11212 14057 11252 15847
rect 11308 14813 11348 16519
rect 11595 16232 11637 16241
rect 11595 16192 11596 16232
rect 11636 16192 11637 16232
rect 11595 16183 11637 16192
rect 11596 15560 11636 16183
rect 11596 15511 11636 15520
rect 11595 14972 11637 14981
rect 11595 14932 11596 14972
rect 11636 14932 11637 14972
rect 11595 14923 11637 14932
rect 11307 14804 11349 14813
rect 11307 14764 11308 14804
rect 11348 14764 11349 14804
rect 11307 14755 11349 14764
rect 11404 14720 11444 14729
rect 11499 14720 11541 14729
rect 11444 14680 11500 14720
rect 11540 14680 11541 14720
rect 11404 14671 11444 14680
rect 11499 14671 11541 14680
rect 11403 14300 11445 14309
rect 11403 14260 11404 14300
rect 11444 14260 11445 14300
rect 11403 14251 11445 14260
rect 11404 14216 11444 14251
rect 11404 14165 11444 14176
rect 11211 14048 11253 14057
rect 11211 14008 11212 14048
rect 11252 14008 11253 14048
rect 11211 13999 11253 14008
rect 11212 13208 11252 13999
rect 11212 11873 11252 13168
rect 11403 13124 11445 13133
rect 11403 13084 11404 13124
rect 11444 13084 11445 13124
rect 11403 13075 11445 13084
rect 11404 12990 11444 13075
rect 11403 12788 11445 12797
rect 11403 12748 11404 12788
rect 11444 12748 11445 12788
rect 11403 12739 11445 12748
rect 11404 12536 11444 12739
rect 11404 12487 11444 12496
rect 11307 12452 11349 12461
rect 11307 12412 11308 12452
rect 11348 12412 11349 12452
rect 11307 12403 11349 12412
rect 11308 12125 11348 12403
rect 11500 12200 11540 14671
rect 11596 14048 11636 14923
rect 11596 13973 11636 14008
rect 11595 13964 11637 13973
rect 11595 13924 11596 13964
rect 11636 13924 11637 13964
rect 11595 13915 11637 13924
rect 11596 13376 11636 13915
rect 11596 13327 11636 13336
rect 11500 12160 11636 12200
rect 11307 12116 11349 12125
rect 11307 12076 11308 12116
rect 11348 12076 11349 12116
rect 11307 12067 11349 12076
rect 11499 12032 11541 12041
rect 11499 11992 11500 12032
rect 11540 11992 11541 12032
rect 11499 11983 11541 11992
rect 11211 11864 11253 11873
rect 11211 11824 11212 11864
rect 11252 11824 11253 11864
rect 11211 11815 11253 11824
rect 11212 11201 11252 11815
rect 11211 11192 11253 11201
rect 11211 11152 11212 11192
rect 11252 11152 11253 11192
rect 11211 11143 11253 11152
rect 11307 11108 11349 11117
rect 11307 11068 11308 11108
rect 11348 11068 11349 11108
rect 11307 11059 11349 11068
rect 11308 11024 11348 11059
rect 11308 10973 11348 10984
rect 11403 11024 11445 11033
rect 11403 10984 11404 11024
rect 11444 10984 11445 11024
rect 11403 10975 11445 10984
rect 11404 10890 11444 10975
rect 11116 10480 11348 10520
rect 10828 10352 10868 10361
rect 11211 10352 11253 10361
rect 10868 10312 11060 10352
rect 10828 10303 10868 10312
rect 11020 10184 11060 10312
rect 11211 10312 11212 10352
rect 11252 10312 11253 10352
rect 11211 10303 11253 10312
rect 10732 10144 10964 10184
rect 10732 8672 10772 10144
rect 10827 10016 10869 10025
rect 10827 9976 10828 10016
rect 10868 9976 10869 10016
rect 10924 10016 10964 10144
rect 11020 10135 11060 10144
rect 11212 10184 11252 10303
rect 11212 10135 11252 10144
rect 11116 10100 11156 10109
rect 11116 10016 11156 10060
rect 10924 9976 11156 10016
rect 10827 9967 10869 9976
rect 10732 8623 10772 8632
rect 10828 8672 10868 9967
rect 10924 9605 10964 9636
rect 10923 9596 10965 9605
rect 10923 9556 10924 9596
rect 10964 9556 10965 9596
rect 10923 9547 10965 9556
rect 10828 8623 10868 8632
rect 10924 9512 10964 9547
rect 10924 7505 10964 9472
rect 11116 9260 11156 9269
rect 11019 9008 11061 9017
rect 11019 8968 11020 9008
rect 11060 8968 11061 9008
rect 11019 8959 11061 8968
rect 11020 8504 11060 8959
rect 11020 8455 11060 8464
rect 11116 8336 11156 9220
rect 11308 8849 11348 10480
rect 11403 10184 11445 10193
rect 11403 10144 11404 10184
rect 11444 10144 11445 10184
rect 11403 10135 11445 10144
rect 11404 10050 11444 10135
rect 11307 8840 11349 8849
rect 11307 8800 11308 8840
rect 11348 8800 11349 8840
rect 11307 8791 11349 8800
rect 11211 8672 11253 8681
rect 11211 8632 11212 8672
rect 11252 8632 11253 8672
rect 11211 8623 11253 8632
rect 11212 8538 11252 8623
rect 11020 8296 11156 8336
rect 11020 8000 11060 8296
rect 11115 8168 11157 8177
rect 11115 8128 11116 8168
rect 11156 8128 11157 8168
rect 11115 8119 11157 8128
rect 11020 7951 11060 7960
rect 11116 8000 11156 8119
rect 11500 8084 11540 11983
rect 11596 11705 11636 12160
rect 11595 11696 11637 11705
rect 11595 11656 11596 11696
rect 11636 11656 11637 11696
rect 11595 11647 11637 11656
rect 11692 11117 11732 17032
rect 11787 16064 11829 16073
rect 11787 16024 11788 16064
rect 11828 16024 11829 16064
rect 11787 16015 11829 16024
rect 11788 12797 11828 16015
rect 11884 14725 11924 14734
rect 11884 14309 11924 14685
rect 11883 14300 11925 14309
rect 11883 14260 11884 14300
rect 11924 14260 11925 14300
rect 11883 14251 11925 14260
rect 11787 12788 11829 12797
rect 11787 12748 11788 12788
rect 11828 12748 11829 12788
rect 11787 12739 11829 12748
rect 11884 12536 11924 12545
rect 11980 12536 12020 20299
rect 12075 17408 12117 17417
rect 12075 17368 12076 17408
rect 12116 17368 12117 17408
rect 12075 17359 12117 17368
rect 12076 17081 12116 17359
rect 12075 17072 12117 17081
rect 12075 17032 12076 17072
rect 12116 17032 12117 17072
rect 12075 17023 12117 17032
rect 12172 15065 12212 20476
rect 12364 20357 12404 20728
rect 12363 20348 12405 20357
rect 12363 20308 12364 20348
rect 12404 20308 12405 20348
rect 12363 20299 12405 20308
rect 12460 20180 12500 25096
rect 12651 25096 12652 25136
rect 12692 25096 12693 25136
rect 12651 25087 12693 25096
rect 12652 23960 12692 25087
rect 12556 23920 12692 23960
rect 12556 23549 12596 23920
rect 12651 23792 12693 23801
rect 12651 23752 12652 23792
rect 12692 23752 12693 23792
rect 12651 23743 12693 23752
rect 12555 23540 12597 23549
rect 12555 23500 12556 23540
rect 12596 23500 12597 23540
rect 12555 23491 12597 23500
rect 12652 23120 12692 23743
rect 12652 22961 12692 23080
rect 12651 22952 12693 22961
rect 12651 22912 12652 22952
rect 12692 22912 12693 22952
rect 12651 22903 12693 22912
rect 12748 22625 12788 25264
rect 12940 24977 12980 25264
rect 13036 25254 13076 25339
rect 13228 25145 13268 28615
rect 13324 27824 13364 28960
rect 13420 28589 13460 31555
rect 13804 30008 13844 32152
rect 13612 29968 13844 30008
rect 13900 30008 13940 38611
rect 13996 38585 14036 38872
rect 14092 38828 14132 38837
rect 14380 38828 14420 38872
rect 14132 38788 14420 38828
rect 14476 38912 14516 38921
rect 14092 38779 14132 38788
rect 13995 38576 14037 38585
rect 13995 38536 13996 38576
rect 14036 38536 14132 38576
rect 13995 38527 14037 38536
rect 13996 38324 14036 38335
rect 13996 38249 14036 38284
rect 13995 38240 14037 38249
rect 13995 38200 13996 38240
rect 14036 38200 14037 38240
rect 13995 38191 14037 38200
rect 14092 36737 14132 38536
rect 14476 38324 14516 38872
rect 14380 38284 14516 38324
rect 14187 37820 14229 37829
rect 14187 37780 14188 37820
rect 14228 37780 14229 37820
rect 14187 37771 14229 37780
rect 14188 37409 14228 37771
rect 14283 37736 14325 37745
rect 14283 37696 14284 37736
rect 14324 37696 14325 37736
rect 14283 37687 14325 37696
rect 14187 37400 14229 37409
rect 14187 37360 14188 37400
rect 14228 37360 14229 37400
rect 14187 37351 14229 37360
rect 14091 36728 14133 36737
rect 14091 36688 14092 36728
rect 14132 36688 14133 36728
rect 14091 36679 14133 36688
rect 14284 36728 14324 37687
rect 14284 36679 14324 36688
rect 14092 35888 14132 36679
rect 14380 36569 14420 38284
rect 14475 38156 14517 38165
rect 14475 38116 14476 38156
rect 14516 38116 14517 38156
rect 14475 38107 14517 38116
rect 14379 36560 14421 36569
rect 14379 36520 14380 36560
rect 14420 36520 14421 36560
rect 14379 36511 14421 36520
rect 14283 36140 14325 36149
rect 14283 36100 14284 36140
rect 14324 36100 14325 36140
rect 14283 36091 14325 36100
rect 14284 36006 14324 36091
rect 14092 35225 14132 35848
rect 14091 35216 14133 35225
rect 14091 35176 14092 35216
rect 14132 35176 14133 35216
rect 14091 35167 14133 35176
rect 14379 35216 14421 35225
rect 14379 35176 14380 35216
rect 14420 35176 14421 35216
rect 14379 35167 14421 35176
rect 14380 35082 14420 35167
rect 14476 34544 14516 38107
rect 14572 37913 14612 42736
rect 14668 42727 14708 42736
rect 14667 42104 14709 42113
rect 14667 42064 14668 42104
rect 14708 42064 14709 42104
rect 14667 42055 14709 42064
rect 14668 40181 14708 42055
rect 14667 40172 14709 40181
rect 14667 40132 14668 40172
rect 14708 40132 14709 40172
rect 14667 40123 14709 40132
rect 14667 40004 14709 40013
rect 14667 39964 14668 40004
rect 14708 39964 14709 40004
rect 14667 39955 14709 39964
rect 14668 39920 14708 39955
rect 14668 39869 14708 39880
rect 14667 39080 14709 39089
rect 14667 39040 14668 39080
rect 14708 39040 14709 39080
rect 14667 39031 14709 39040
rect 14668 38417 14708 39031
rect 14667 38408 14709 38417
rect 14667 38368 14668 38408
rect 14708 38368 14709 38408
rect 14667 38359 14709 38368
rect 14667 38240 14709 38249
rect 14667 38200 14668 38240
rect 14708 38200 14709 38240
rect 14667 38191 14709 38200
rect 14668 38106 14708 38191
rect 14571 37904 14613 37913
rect 14571 37864 14572 37904
rect 14612 37864 14613 37904
rect 14571 37855 14613 37864
rect 14764 36812 14804 45088
rect 14860 44965 14900 44974
rect 14860 44633 14900 44925
rect 14859 44624 14901 44633
rect 14859 44584 14860 44624
rect 14900 44584 14901 44624
rect 14859 44575 14901 44584
rect 14956 43961 14996 46852
rect 15148 46565 15188 48700
rect 15147 46556 15189 46565
rect 15147 46516 15148 46556
rect 15188 46516 15189 46556
rect 15532 46556 15572 48784
rect 15628 46640 15668 49195
rect 15916 48740 15956 48749
rect 15916 48245 15956 48700
rect 16012 48740 16052 48749
rect 16108 48740 16148 49624
rect 16052 48700 16148 48740
rect 16012 48691 16052 48700
rect 15915 48236 15957 48245
rect 15915 48196 15916 48236
rect 15956 48196 15957 48236
rect 15915 48187 15957 48196
rect 16011 47984 16053 47993
rect 16011 47944 16012 47984
rect 16052 47944 16053 47984
rect 16011 47935 16053 47944
rect 16012 47850 16052 47935
rect 15628 46600 15764 46640
rect 15532 46516 15668 46556
rect 15147 46507 15189 46516
rect 15339 46472 15381 46481
rect 15339 46432 15340 46472
rect 15380 46432 15381 46472
rect 15339 46423 15381 46432
rect 15051 46388 15093 46397
rect 15051 46348 15052 46388
rect 15092 46348 15093 46388
rect 15051 46339 15093 46348
rect 15243 46388 15285 46397
rect 15243 46348 15244 46388
rect 15284 46348 15285 46388
rect 15243 46339 15285 46348
rect 15052 45305 15092 46339
rect 15244 45893 15284 46339
rect 15340 46313 15380 46423
rect 15339 46304 15381 46313
rect 15339 46264 15340 46304
rect 15380 46264 15381 46304
rect 15339 46255 15381 46264
rect 15243 45884 15285 45893
rect 15243 45844 15244 45884
rect 15284 45844 15285 45884
rect 15243 45835 15285 45844
rect 15628 45809 15668 46516
rect 15532 45800 15572 45809
rect 15532 45557 15572 45760
rect 15627 45800 15669 45809
rect 15627 45760 15628 45800
rect 15668 45760 15669 45800
rect 15627 45751 15669 45760
rect 15628 45666 15668 45751
rect 15531 45548 15573 45557
rect 15531 45508 15532 45548
rect 15572 45508 15573 45548
rect 15531 45499 15573 45508
rect 15243 45464 15285 45473
rect 15243 45424 15244 45464
rect 15284 45424 15285 45464
rect 15243 45415 15285 45424
rect 15244 45305 15284 45415
rect 15051 45296 15093 45305
rect 15051 45256 15052 45296
rect 15092 45256 15093 45296
rect 15051 45247 15093 45256
rect 15243 45296 15285 45305
rect 15243 45256 15244 45296
rect 15284 45256 15285 45296
rect 15243 45247 15285 45256
rect 15244 44960 15284 44969
rect 15052 44750 15092 44759
rect 15052 44540 15092 44710
rect 15052 44500 15188 44540
rect 15148 44297 15188 44500
rect 15244 44465 15284 44920
rect 15436 44960 15476 44969
rect 15340 44792 15380 44801
rect 15243 44456 15285 44465
rect 15243 44416 15244 44456
rect 15284 44416 15285 44456
rect 15243 44407 15285 44416
rect 15147 44288 15189 44297
rect 15147 44248 15148 44288
rect 15188 44248 15189 44288
rect 15147 44239 15189 44248
rect 15051 44204 15093 44213
rect 15051 44164 15052 44204
rect 15092 44164 15093 44204
rect 15051 44155 15093 44164
rect 14955 43952 14997 43961
rect 14955 43912 14956 43952
rect 14996 43912 14997 43952
rect 14955 43903 14997 43912
rect 14955 42020 14997 42029
rect 14955 41980 14956 42020
rect 14996 41980 14997 42020
rect 14955 41971 14997 41980
rect 14859 41936 14901 41945
rect 14859 41896 14860 41936
rect 14900 41896 14901 41936
rect 14859 41887 14901 41896
rect 14860 41180 14900 41887
rect 14956 41264 14996 41971
rect 14956 41215 14996 41224
rect 14860 40676 14900 41140
rect 15052 40760 15092 44155
rect 15340 43457 15380 44752
rect 15436 44297 15476 44920
rect 15435 44288 15477 44297
rect 15435 44248 15436 44288
rect 15476 44248 15477 44288
rect 15435 44239 15477 44248
rect 15339 43448 15381 43457
rect 15339 43408 15340 43448
rect 15380 43408 15381 43448
rect 15339 43399 15381 43408
rect 15724 42029 15764 46600
rect 15915 46388 15957 46397
rect 15915 46348 15916 46388
rect 15956 46348 15957 46388
rect 15915 46339 15957 46348
rect 15819 45800 15861 45809
rect 15819 45760 15820 45800
rect 15860 45760 15861 45800
rect 15819 45751 15861 45760
rect 15820 45473 15860 45751
rect 15819 45464 15861 45473
rect 15819 45424 15820 45464
rect 15860 45424 15861 45464
rect 15819 45415 15861 45424
rect 15916 44288 15956 46339
rect 16108 45977 16148 48700
rect 16204 48236 16244 50287
rect 16300 49496 16340 51547
rect 16395 51260 16437 51269
rect 16395 51220 16396 51260
rect 16436 51220 16437 51260
rect 16395 51211 16437 51220
rect 16396 50261 16436 51211
rect 16395 50252 16437 50261
rect 16395 50212 16396 50252
rect 16436 50212 16437 50252
rect 16395 50203 16437 50212
rect 16395 49916 16437 49925
rect 16395 49876 16396 49916
rect 16436 49876 16437 49916
rect 16395 49867 16437 49876
rect 16300 48917 16340 49456
rect 16396 49496 16436 49867
rect 16396 49447 16436 49456
rect 16395 49244 16437 49253
rect 16395 49204 16396 49244
rect 16436 49204 16437 49244
rect 16395 49195 16437 49204
rect 16299 48908 16341 48917
rect 16299 48868 16300 48908
rect 16340 48868 16341 48908
rect 16299 48859 16341 48868
rect 16300 48497 16340 48859
rect 16299 48488 16341 48497
rect 16299 48448 16300 48488
rect 16340 48448 16341 48488
rect 16299 48439 16341 48448
rect 16396 48404 16436 49195
rect 16492 48824 16532 48833
rect 16492 48665 16532 48784
rect 16491 48656 16533 48665
rect 16491 48616 16492 48656
rect 16532 48616 16533 48656
rect 16491 48607 16533 48616
rect 16396 48364 16532 48404
rect 16204 48187 16244 48196
rect 16395 48152 16437 48161
rect 16395 48112 16396 48152
rect 16436 48112 16437 48152
rect 16395 48103 16437 48112
rect 16203 47984 16245 47993
rect 16203 47944 16204 47984
rect 16244 47944 16245 47984
rect 16203 47935 16245 47944
rect 16396 47984 16436 48103
rect 16396 47935 16436 47944
rect 16492 47984 16532 48364
rect 16204 47312 16244 47935
rect 16299 47480 16341 47489
rect 16299 47440 16300 47480
rect 16340 47440 16341 47480
rect 16299 47431 16341 47440
rect 16396 47480 16436 47489
rect 16492 47480 16532 47944
rect 16436 47440 16532 47480
rect 16396 47431 16436 47440
rect 16204 46901 16244 47272
rect 16203 46892 16245 46901
rect 16203 46852 16204 46892
rect 16244 46852 16245 46892
rect 16203 46843 16245 46852
rect 16107 45968 16149 45977
rect 16107 45928 16108 45968
rect 16148 45928 16149 45968
rect 16107 45919 16149 45928
rect 16011 45800 16053 45809
rect 16011 45760 16012 45800
rect 16052 45760 16053 45800
rect 16011 45751 16053 45760
rect 16108 45800 16148 45919
rect 16108 45751 16148 45760
rect 16012 45666 16052 45751
rect 16107 45548 16149 45557
rect 16107 45508 16108 45548
rect 16148 45508 16149 45548
rect 16107 45499 16149 45508
rect 16108 44456 16148 45499
rect 16300 45221 16340 47431
rect 16588 47405 16628 52144
rect 16683 52100 16725 52109
rect 16683 52060 16684 52100
rect 16724 52060 16725 52100
rect 16683 52051 16725 52060
rect 16684 51848 16724 52051
rect 16780 51941 16820 53320
rect 16876 53311 16916 53320
rect 16972 53360 17012 53479
rect 16972 53311 17012 53320
rect 17067 53360 17109 53369
rect 17067 53320 17068 53360
rect 17108 53320 17109 53360
rect 17067 53311 17109 53320
rect 17164 53360 17204 53479
rect 17164 53311 17204 53320
rect 17068 53226 17108 53311
rect 17067 53108 17109 53117
rect 17067 53068 17068 53108
rect 17108 53068 17109 53108
rect 17067 53059 17109 53068
rect 16875 52856 16917 52865
rect 16875 52816 16876 52856
rect 16916 52816 16917 52856
rect 16875 52807 16917 52816
rect 16876 52520 16916 52807
rect 16971 52688 17013 52697
rect 16971 52648 16972 52688
rect 17012 52648 17013 52688
rect 16971 52639 17013 52648
rect 16876 52471 16916 52480
rect 16875 52184 16917 52193
rect 16875 52144 16876 52184
rect 16916 52144 16917 52184
rect 16875 52135 16917 52144
rect 16779 51932 16821 51941
rect 16779 51892 16780 51932
rect 16820 51892 16821 51932
rect 16779 51883 16821 51892
rect 16684 51799 16724 51808
rect 16780 51764 16820 51773
rect 16876 51764 16916 52135
rect 16820 51724 16916 51764
rect 16780 51715 16820 51724
rect 16779 51596 16821 51605
rect 16779 51556 16780 51596
rect 16820 51556 16821 51596
rect 16779 51547 16821 51556
rect 16683 51008 16725 51017
rect 16683 50968 16684 51008
rect 16724 50968 16725 51008
rect 16683 50959 16725 50968
rect 16780 51008 16820 51547
rect 16972 51008 17012 52639
rect 17068 52529 17108 53059
rect 17164 52697 17204 52782
rect 17163 52688 17205 52697
rect 17163 52648 17164 52688
rect 17204 52648 17205 52688
rect 17163 52639 17205 52648
rect 17067 52520 17109 52529
rect 17067 52480 17068 52520
rect 17108 52480 17109 52520
rect 17067 52471 17109 52480
rect 17164 52520 17204 52529
rect 17067 51764 17109 51773
rect 17067 51724 17068 51764
rect 17108 51724 17109 51764
rect 17067 51715 17109 51724
rect 16684 49748 16724 50959
rect 16684 49699 16724 49708
rect 16780 50336 16820 50968
rect 16780 48665 16820 50296
rect 16876 50968 17012 51008
rect 16779 48656 16821 48665
rect 16779 48616 16780 48656
rect 16820 48616 16821 48656
rect 16779 48607 16821 48616
rect 16683 48320 16725 48329
rect 16683 48280 16684 48320
rect 16724 48280 16725 48320
rect 16683 48271 16725 48280
rect 16684 47816 16724 48271
rect 16684 47767 16724 47776
rect 16876 47732 16916 50968
rect 16972 50840 17012 50849
rect 16972 50681 17012 50800
rect 16971 50672 17013 50681
rect 16971 50632 16972 50672
rect 17012 50632 17013 50672
rect 16971 50623 17013 50632
rect 16972 50504 17012 50513
rect 17068 50504 17108 51715
rect 17164 51521 17204 52480
rect 17260 51848 17300 53647
rect 17548 53360 17588 54151
rect 17643 54032 17685 54041
rect 17643 53992 17644 54032
rect 17684 53992 17685 54032
rect 17643 53983 17685 53992
rect 17740 54032 17780 55000
rect 17835 54991 17877 55000
rect 17836 54906 17876 54991
rect 17932 54872 17972 55336
rect 18316 55292 18356 56260
rect 18412 56251 18452 56260
rect 18411 55964 18453 55973
rect 18411 55924 18412 55964
rect 18452 55924 18453 55964
rect 18411 55915 18453 55924
rect 18412 55544 18452 55915
rect 18412 55495 18452 55504
rect 18220 55252 18356 55292
rect 18124 55049 18164 55134
rect 18123 55040 18165 55049
rect 18123 55000 18124 55040
rect 18164 55000 18165 55040
rect 18123 54991 18165 55000
rect 17932 54823 17972 54832
rect 18220 54209 18260 55252
rect 18508 55208 18548 56344
rect 18988 56335 19028 56344
rect 18808 55964 19176 55973
rect 18848 55924 18890 55964
rect 18930 55924 18972 55964
rect 19012 55924 19054 55964
rect 19094 55924 19136 55964
rect 18808 55915 19176 55924
rect 18316 55168 18548 55208
rect 18219 54200 18261 54209
rect 18219 54160 18220 54200
rect 18260 54160 18261 54200
rect 18219 54151 18261 54160
rect 17644 53898 17684 53983
rect 17740 53537 17780 53992
rect 17931 54032 17973 54041
rect 17931 53992 17932 54032
rect 17972 53992 17973 54032
rect 17931 53983 17973 53992
rect 17739 53528 17781 53537
rect 17739 53488 17740 53528
rect 17780 53488 17781 53528
rect 17739 53479 17781 53488
rect 17548 53311 17588 53320
rect 17644 53360 17684 53369
rect 17548 52865 17588 52884
rect 17547 52856 17589 52865
rect 17644 52856 17684 53320
rect 17740 53360 17780 53369
rect 17740 53033 17780 53320
rect 17836 53360 17876 53369
rect 17739 53024 17781 53033
rect 17739 52984 17740 53024
rect 17780 52984 17781 53024
rect 17739 52975 17781 52984
rect 17547 52816 17548 52856
rect 17588 52816 17684 52856
rect 17547 52807 17589 52816
rect 17836 52772 17876 53320
rect 17644 52732 17876 52772
rect 17547 52688 17589 52697
rect 17547 52648 17548 52688
rect 17588 52648 17589 52688
rect 17547 52639 17589 52648
rect 17260 51799 17300 51808
rect 17356 52520 17396 52529
rect 17356 51773 17396 52480
rect 17548 52520 17588 52639
rect 17548 52471 17588 52480
rect 17644 52520 17684 52732
rect 17932 52688 17972 53983
rect 18316 53957 18356 55168
rect 18507 55040 18549 55049
rect 18507 55000 18508 55040
rect 18548 55000 18549 55040
rect 18507 54991 18549 55000
rect 18508 54906 18548 54991
rect 18700 54872 18740 54881
rect 18508 54620 18548 54629
rect 18412 54580 18508 54620
rect 18412 54046 18452 54580
rect 18508 54571 18548 54580
rect 18412 53997 18452 54006
rect 18315 53948 18357 53957
rect 18315 53908 18316 53948
rect 18356 53908 18357 53948
rect 18315 53899 18357 53908
rect 18220 53864 18260 53873
rect 18027 53360 18069 53369
rect 18027 53320 18028 53360
rect 18068 53320 18069 53360
rect 18027 53311 18069 53320
rect 18028 52865 18068 53311
rect 18220 52949 18260 53824
rect 18700 53369 18740 54832
rect 18808 54452 19176 54461
rect 18848 54412 18890 54452
rect 18930 54412 18972 54452
rect 19012 54412 19054 54452
rect 19094 54412 19136 54452
rect 18808 54403 19176 54412
rect 18891 54032 18933 54041
rect 18891 53992 18892 54032
rect 18932 53992 18933 54032
rect 18891 53983 18933 53992
rect 18892 53898 18932 53983
rect 19276 53864 19316 56839
rect 19372 55553 19412 57091
rect 19468 56981 19508 57856
rect 19564 57401 19604 58612
rect 19755 58612 19756 58652
rect 19796 58612 19797 58652
rect 19755 58603 19797 58612
rect 19756 58518 19796 58603
rect 19660 57896 19700 57905
rect 19700 57856 19796 57896
rect 19660 57847 19700 57856
rect 19660 57644 19700 57653
rect 19563 57392 19605 57401
rect 19563 57352 19564 57392
rect 19604 57352 19605 57392
rect 19563 57343 19605 57352
rect 19660 57317 19700 57604
rect 19659 57308 19701 57317
rect 19659 57268 19660 57308
rect 19700 57268 19701 57308
rect 19659 57259 19701 57268
rect 19563 57140 19605 57149
rect 19756 57140 19796 57856
rect 19852 57812 19892 59359
rect 19947 59156 19989 59165
rect 19947 59116 19948 59156
rect 19988 59116 19989 59156
rect 19947 59107 19989 59116
rect 19948 58820 19988 59107
rect 20715 58904 20757 58913
rect 20715 58864 20716 58904
rect 20756 58864 20757 58904
rect 20715 58855 20757 58864
rect 19948 58771 19988 58780
rect 20048 58232 20416 58241
rect 20088 58192 20130 58232
rect 20170 58192 20212 58232
rect 20252 58192 20294 58232
rect 20334 58192 20376 58232
rect 20048 58183 20416 58192
rect 20716 58157 20756 58855
rect 20715 58148 20757 58157
rect 20715 58108 20716 58148
rect 20756 58108 20757 58148
rect 20715 58099 20757 58108
rect 20619 57896 20661 57905
rect 20619 57856 20620 57896
rect 20660 57856 20661 57896
rect 20619 57847 20661 57856
rect 19852 57763 19892 57772
rect 19947 57812 19989 57821
rect 19947 57772 19948 57812
rect 19988 57772 19989 57812
rect 19947 57763 19989 57772
rect 19948 57476 19988 57763
rect 20043 57728 20085 57737
rect 20043 57688 20044 57728
rect 20084 57688 20085 57728
rect 20043 57679 20085 57688
rect 20044 57594 20084 57679
rect 20235 57644 20277 57653
rect 20235 57604 20236 57644
rect 20276 57604 20277 57644
rect 20235 57595 20277 57604
rect 19948 57436 20084 57476
rect 20044 57392 20084 57436
rect 20044 57352 20180 57392
rect 19948 57233 19988 57318
rect 19947 57224 19989 57233
rect 19947 57184 19948 57224
rect 19988 57184 19989 57224
rect 19947 57175 19989 57184
rect 19563 57100 19564 57140
rect 19604 57100 19605 57140
rect 19563 57091 19605 57100
rect 19660 57100 19796 57140
rect 19564 57056 19604 57091
rect 19564 57005 19604 57016
rect 19467 56972 19509 56981
rect 19467 56932 19468 56972
rect 19508 56932 19509 56972
rect 19467 56923 19509 56932
rect 19660 56552 19700 57100
rect 20140 57070 20180 57352
rect 19947 57056 19989 57065
rect 19947 57016 19948 57056
rect 19988 57016 19989 57056
rect 20140 57021 20180 57030
rect 20236 57056 20276 57595
rect 19947 57007 19989 57016
rect 20236 57007 20276 57016
rect 19755 56972 19797 56981
rect 19755 56932 19756 56972
rect 19796 56932 19797 56972
rect 19755 56923 19797 56932
rect 19756 56838 19796 56923
rect 19948 56922 19988 57007
rect 20048 56720 20416 56729
rect 20088 56680 20130 56720
rect 20170 56680 20212 56720
rect 20252 56680 20294 56720
rect 20334 56680 20376 56720
rect 20048 56671 20416 56680
rect 19660 56503 19700 56512
rect 19468 56393 19508 56494
rect 19467 56384 19509 56393
rect 19852 56384 19892 56393
rect 19467 56335 19468 56384
rect 19508 56335 19509 56384
rect 19564 56344 19852 56384
rect 19468 55805 19508 56330
rect 19467 55796 19509 55805
rect 19467 55756 19468 55796
rect 19508 55756 19509 55796
rect 19467 55747 19509 55756
rect 19371 55544 19413 55553
rect 19371 55504 19372 55544
rect 19412 55504 19413 55544
rect 19371 55495 19413 55504
rect 19564 55049 19604 56344
rect 19852 56335 19892 56344
rect 20044 56384 20084 56393
rect 19852 56132 19892 56141
rect 19756 56092 19852 56132
rect 19660 55553 19700 55638
rect 19659 55544 19701 55553
rect 19659 55504 19660 55544
rect 19700 55504 19701 55544
rect 19659 55495 19701 55504
rect 19563 55040 19605 55049
rect 19563 55000 19564 55040
rect 19604 55000 19605 55040
rect 19563 54991 19605 55000
rect 19371 54788 19413 54797
rect 19371 54748 19372 54788
rect 19412 54748 19413 54788
rect 19371 54739 19413 54748
rect 19372 54116 19412 54739
rect 19372 54067 19412 54076
rect 19468 54032 19508 54041
rect 19276 53824 19412 53864
rect 18411 53360 18453 53369
rect 18411 53320 18412 53360
rect 18452 53320 18453 53360
rect 18411 53311 18453 53320
rect 18699 53360 18741 53369
rect 18699 53320 18700 53360
rect 18740 53320 18741 53360
rect 18699 53311 18741 53320
rect 19275 53360 19317 53369
rect 19275 53320 19276 53360
rect 19316 53320 19317 53360
rect 19275 53311 19317 53320
rect 18219 52940 18261 52949
rect 18219 52900 18220 52940
rect 18260 52900 18261 52940
rect 18219 52891 18261 52900
rect 18027 52856 18069 52865
rect 18027 52816 18028 52856
rect 18068 52816 18069 52856
rect 18027 52807 18069 52816
rect 18219 52772 18261 52781
rect 18219 52732 18220 52772
rect 18260 52732 18261 52772
rect 18219 52723 18261 52732
rect 17644 52471 17684 52480
rect 17740 52648 17972 52688
rect 17452 52436 17492 52445
rect 17355 51764 17397 51773
rect 17355 51724 17356 51764
rect 17396 51724 17397 51764
rect 17355 51715 17397 51724
rect 17259 51596 17301 51605
rect 17259 51556 17260 51596
rect 17300 51556 17301 51596
rect 17259 51547 17301 51556
rect 17163 51512 17205 51521
rect 17163 51472 17164 51512
rect 17204 51472 17205 51512
rect 17163 51463 17205 51472
rect 17012 50464 17108 50504
rect 16972 50455 17012 50464
rect 17260 50420 17300 51547
rect 17452 51185 17492 52396
rect 17740 52352 17780 52648
rect 18028 52529 18068 52614
rect 17644 52312 17780 52352
rect 17836 52520 17876 52529
rect 17547 51680 17589 51689
rect 17644 51680 17684 52312
rect 17740 51834 17780 51859
rect 17740 51773 17780 51794
rect 17739 51764 17781 51773
rect 17739 51724 17740 51764
rect 17780 51724 17781 51764
rect 17739 51715 17781 51724
rect 17547 51640 17548 51680
rect 17588 51640 17684 51680
rect 17547 51631 17589 51640
rect 17644 51596 17684 51640
rect 17644 51556 17780 51596
rect 17451 51176 17493 51185
rect 17451 51136 17452 51176
rect 17492 51136 17493 51176
rect 17451 51127 17493 51136
rect 17356 51008 17396 51017
rect 17356 50513 17396 50968
rect 17548 51008 17588 51017
rect 17452 50840 17492 50849
rect 17355 50504 17397 50513
rect 17355 50464 17356 50504
rect 17396 50464 17397 50504
rect 17355 50455 17397 50464
rect 17068 50380 17300 50420
rect 16971 50252 17013 50261
rect 16971 50212 16972 50252
rect 17012 50212 17013 50252
rect 16971 50203 17013 50212
rect 16972 49496 17012 50203
rect 16972 49447 17012 49456
rect 16971 49244 17013 49253
rect 16971 49204 16972 49244
rect 17012 49204 17013 49244
rect 16971 49195 17013 49204
rect 16972 48819 17012 49195
rect 16972 48770 17012 48779
rect 16972 47993 17012 48078
rect 16971 47984 17013 47993
rect 16971 47944 16972 47984
rect 17012 47944 17013 47984
rect 16971 47935 17013 47944
rect 17068 47816 17108 50380
rect 17355 50336 17397 50345
rect 17164 50323 17204 50332
rect 17355 50296 17356 50336
rect 17396 50296 17397 50336
rect 17355 50287 17397 50296
rect 17164 50252 17204 50283
rect 17164 50212 17300 50252
rect 17164 50084 17204 50093
rect 17164 49505 17204 50044
rect 17163 49496 17205 49505
rect 17163 49456 17164 49496
rect 17204 49456 17205 49496
rect 17163 49447 17205 49456
rect 17164 48992 17204 49001
rect 17260 48992 17300 50212
rect 17356 50202 17396 50287
rect 17452 49589 17492 50800
rect 17548 50513 17588 50968
rect 17643 51008 17685 51017
rect 17643 50968 17644 51008
rect 17684 50968 17685 51008
rect 17643 50959 17685 50968
rect 17644 50874 17684 50959
rect 17643 50756 17685 50765
rect 17643 50716 17644 50756
rect 17684 50716 17685 50756
rect 17643 50707 17685 50716
rect 17547 50504 17589 50513
rect 17547 50464 17548 50504
rect 17588 50464 17589 50504
rect 17547 50455 17589 50464
rect 17548 50336 17588 50345
rect 17644 50336 17684 50707
rect 17588 50296 17684 50336
rect 17548 50287 17588 50296
rect 17643 50168 17685 50177
rect 17643 50128 17644 50168
rect 17684 50128 17685 50168
rect 17643 50119 17685 50128
rect 17644 49673 17684 50119
rect 17643 49664 17685 49673
rect 17643 49624 17644 49664
rect 17684 49624 17685 49664
rect 17643 49615 17685 49624
rect 17451 49580 17493 49589
rect 17451 49540 17452 49580
rect 17492 49540 17493 49580
rect 17451 49531 17493 49540
rect 17547 49244 17589 49253
rect 17547 49204 17548 49244
rect 17588 49204 17589 49244
rect 17547 49195 17589 49204
rect 17355 49160 17397 49169
rect 17355 49120 17356 49160
rect 17396 49120 17397 49160
rect 17355 49111 17397 49120
rect 17204 48952 17300 48992
rect 17356 48992 17396 49111
rect 17164 48943 17204 48952
rect 17356 48943 17396 48952
rect 17452 48824 17492 48833
rect 17452 48329 17492 48784
rect 17548 48824 17588 49195
rect 17548 48775 17588 48784
rect 17644 48824 17684 49615
rect 17740 48824 17780 51556
rect 17836 51008 17876 52480
rect 18027 52520 18069 52529
rect 18027 52480 18028 52520
rect 18068 52480 18069 52520
rect 18027 52471 18069 52480
rect 18220 52445 18260 52723
rect 18412 52520 18452 53311
rect 19276 53226 19316 53311
rect 18808 52940 19176 52949
rect 18848 52900 18890 52940
rect 18930 52900 18972 52940
rect 19012 52900 19054 52940
rect 19094 52900 19136 52940
rect 18808 52891 19176 52900
rect 18699 52856 18741 52865
rect 18699 52816 18700 52856
rect 18740 52816 18741 52856
rect 18699 52807 18741 52816
rect 18452 52480 18644 52520
rect 18412 52471 18452 52480
rect 18219 52436 18261 52445
rect 18219 52396 18220 52436
rect 18260 52396 18261 52436
rect 18219 52387 18261 52396
rect 17931 52352 17973 52361
rect 17931 52312 17932 52352
rect 17972 52312 17973 52352
rect 17931 52303 17973 52312
rect 18507 52352 18549 52361
rect 18507 52312 18508 52352
rect 18548 52312 18549 52352
rect 18507 52303 18549 52312
rect 17932 52218 17972 52303
rect 17932 52016 17972 52025
rect 17972 51976 18453 52016
rect 17932 51967 17972 51976
rect 18413 51863 18453 51976
rect 18124 51848 18164 51857
rect 18164 51808 18260 51848
rect 18413 51814 18453 51823
rect 18124 51799 18164 51808
rect 18220 51689 18260 51808
rect 18315 51764 18357 51773
rect 18315 51724 18316 51764
rect 18356 51724 18357 51764
rect 18315 51715 18357 51724
rect 18219 51680 18261 51689
rect 18219 51640 18220 51680
rect 18260 51640 18261 51680
rect 18219 51631 18261 51640
rect 18124 51596 18164 51605
rect 18028 51185 18068 51270
rect 18027 51176 18069 51185
rect 18027 51136 18028 51176
rect 18068 51136 18069 51176
rect 18027 51127 18069 51136
rect 18028 51008 18068 51017
rect 18124 51008 18164 51556
rect 17836 50968 17972 51008
rect 17835 50840 17877 50849
rect 17835 50800 17836 50840
rect 17876 50800 17877 50840
rect 17835 50791 17877 50800
rect 17836 50706 17876 50791
rect 17836 48992 17876 49001
rect 17932 48992 17972 50968
rect 18068 50968 18164 51008
rect 18028 50959 18068 50968
rect 18220 50681 18260 51631
rect 18219 50672 18261 50681
rect 18219 50632 18220 50672
rect 18260 50632 18261 50672
rect 18219 50623 18261 50632
rect 18123 50168 18165 50177
rect 18123 50128 18124 50168
rect 18164 50128 18165 50168
rect 18123 50119 18165 50128
rect 18124 49589 18164 50119
rect 18123 49580 18165 49589
rect 18123 49540 18124 49580
rect 18164 49540 18165 49580
rect 18123 49531 18165 49540
rect 18027 49328 18069 49337
rect 18027 49288 18028 49328
rect 18068 49288 18069 49328
rect 18027 49279 18069 49288
rect 17876 48952 17972 48992
rect 17836 48943 17876 48952
rect 17740 48784 17876 48824
rect 17644 48775 17684 48784
rect 17547 48656 17589 48665
rect 17547 48616 17548 48656
rect 17588 48616 17589 48656
rect 17547 48607 17589 48616
rect 17451 48320 17493 48329
rect 17451 48280 17452 48320
rect 17492 48280 17493 48320
rect 17451 48271 17493 48280
rect 16780 47692 16916 47732
rect 16972 47776 17108 47816
rect 16587 47396 16629 47405
rect 16587 47356 16588 47396
rect 16628 47356 16629 47396
rect 16587 47347 16629 47356
rect 16780 47312 16820 47692
rect 16875 47396 16917 47405
rect 16875 47356 16876 47396
rect 16916 47356 16917 47396
rect 16875 47347 16917 47356
rect 16683 47060 16725 47069
rect 16683 47020 16684 47060
rect 16724 47020 16725 47060
rect 16683 47011 16725 47020
rect 16588 46472 16628 46483
rect 16588 46397 16628 46432
rect 16587 46388 16629 46397
rect 16587 46348 16588 46388
rect 16628 46348 16629 46388
rect 16587 46339 16629 46348
rect 16587 46052 16629 46061
rect 16587 46012 16588 46052
rect 16628 46012 16629 46052
rect 16587 46003 16629 46012
rect 16588 45800 16628 46003
rect 16588 45751 16628 45760
rect 16299 45212 16341 45221
rect 16299 45172 16300 45212
rect 16340 45172 16341 45212
rect 16299 45163 16341 45172
rect 16684 44960 16724 47011
rect 16780 46481 16820 47272
rect 16779 46472 16821 46481
rect 16779 46432 16780 46472
rect 16820 46432 16821 46472
rect 16779 46423 16821 46432
rect 16779 46304 16821 46313
rect 16779 46264 16780 46304
rect 16820 46264 16821 46304
rect 16779 46255 16821 46264
rect 16780 46170 16820 46255
rect 16779 45632 16821 45641
rect 16779 45592 16780 45632
rect 16820 45592 16821 45632
rect 16779 45583 16821 45592
rect 16684 44911 16724 44920
rect 16300 44792 16340 44801
rect 16108 44407 16148 44416
rect 16203 44456 16245 44465
rect 16203 44416 16204 44456
rect 16244 44416 16245 44456
rect 16203 44407 16245 44416
rect 15916 43448 15956 44248
rect 16108 43700 16148 43709
rect 16204 43700 16244 44407
rect 16148 43660 16244 43700
rect 16300 44120 16340 44752
rect 16780 44540 16820 45583
rect 16684 44500 16820 44540
rect 16684 44120 16724 44500
rect 16780 44297 16820 44382
rect 16876 44372 16916 47347
rect 16972 46472 17012 47776
rect 17068 46481 17108 46566
rect 16972 45053 17012 46432
rect 17067 46472 17109 46481
rect 17067 46432 17068 46472
rect 17108 46432 17109 46472
rect 17067 46423 17109 46432
rect 17164 46472 17204 46481
rect 17067 46304 17109 46313
rect 17067 46264 17068 46304
rect 17108 46264 17109 46304
rect 17067 46255 17109 46264
rect 17068 45809 17108 46255
rect 17067 45800 17109 45809
rect 17067 45755 17068 45800
rect 17108 45755 17109 45800
rect 17067 45751 17109 45755
rect 17068 45666 17108 45751
rect 16971 45044 17013 45053
rect 16971 45004 16972 45044
rect 17012 45004 17013 45044
rect 16971 44995 17013 45004
rect 17164 44465 17204 46432
rect 17451 46472 17493 46481
rect 17451 46432 17452 46472
rect 17492 46432 17493 46472
rect 17451 46423 17493 46432
rect 17259 46304 17301 46313
rect 17259 46264 17260 46304
rect 17300 46264 17301 46304
rect 17259 46255 17301 46264
rect 17260 46170 17300 46255
rect 17260 45884 17300 45893
rect 17300 45844 17396 45884
rect 17260 45835 17300 45844
rect 17163 44456 17205 44465
rect 17163 44416 17164 44456
rect 17204 44416 17205 44456
rect 17163 44407 17205 44416
rect 16876 44332 17012 44372
rect 16779 44288 16821 44297
rect 16779 44248 16780 44288
rect 16820 44248 16821 44288
rect 16779 44239 16821 44248
rect 16780 44120 16820 44129
rect 16684 44080 16780 44120
rect 16108 43651 16148 43660
rect 15820 43408 15916 43448
rect 15723 42020 15765 42029
rect 15723 41980 15724 42020
rect 15764 41980 15765 42020
rect 15723 41971 15765 41980
rect 15436 41936 15476 41945
rect 15436 41525 15476 41896
rect 15820 41852 15860 43408
rect 15916 43399 15956 43408
rect 16300 43280 16340 44080
rect 16780 44071 16820 44080
rect 16588 44036 16628 44045
rect 16300 42944 16340 43240
rect 16300 42895 16340 42904
rect 16492 43996 16588 44036
rect 15915 42776 15957 42785
rect 15915 42736 15916 42776
rect 15956 42736 15957 42776
rect 15915 42727 15957 42736
rect 16299 42776 16341 42785
rect 16299 42736 16300 42776
rect 16340 42736 16341 42776
rect 16299 42727 16341 42736
rect 15916 42642 15956 42727
rect 16108 42524 16148 42533
rect 16108 42020 16148 42484
rect 15964 41980 16148 42020
rect 15964 41978 16004 41980
rect 16300 41945 16340 42727
rect 16396 42608 16436 42617
rect 15964 41929 16004 41938
rect 16299 41936 16341 41945
rect 16299 41896 16300 41936
rect 16340 41896 16341 41936
rect 16299 41887 16341 41896
rect 16396 41861 16436 42568
rect 16492 42104 16532 43996
rect 16588 43987 16628 43996
rect 16587 43448 16629 43457
rect 16587 43408 16588 43448
rect 16628 43408 16629 43448
rect 16587 43399 16629 43408
rect 16780 43448 16820 43457
rect 16588 43314 16628 43399
rect 16684 43280 16724 43289
rect 16684 42869 16724 43240
rect 16780 43205 16820 43408
rect 16876 43448 16916 43457
rect 16876 43289 16916 43408
rect 16875 43280 16917 43289
rect 16875 43240 16876 43280
rect 16916 43240 16917 43280
rect 16875 43231 16917 43240
rect 16779 43196 16821 43205
rect 16779 43156 16780 43196
rect 16820 43156 16821 43196
rect 16779 43147 16821 43156
rect 16683 42860 16725 42869
rect 16683 42820 16684 42860
rect 16724 42820 16725 42860
rect 16683 42811 16725 42820
rect 16492 42064 16628 42104
rect 16491 41936 16533 41945
rect 16491 41896 16492 41936
rect 16532 41896 16533 41936
rect 16491 41887 16533 41896
rect 15724 41812 15860 41852
rect 16395 41852 16437 41861
rect 16395 41812 16396 41852
rect 16436 41812 16437 41852
rect 15627 41768 15669 41777
rect 15627 41728 15628 41768
rect 15668 41728 15669 41768
rect 15627 41719 15669 41728
rect 15435 41516 15477 41525
rect 15435 41476 15436 41516
rect 15476 41476 15477 41516
rect 15435 41467 15477 41476
rect 15436 41264 15476 41467
rect 15436 41215 15476 41224
rect 15052 40720 15188 40760
rect 14860 40636 15092 40676
rect 14955 40508 14997 40517
rect 14955 40468 14956 40508
rect 14996 40468 14997 40508
rect 14955 40459 14997 40468
rect 14859 40424 14901 40433
rect 14859 40384 14860 40424
rect 14900 40384 14901 40424
rect 14859 40375 14901 40384
rect 14860 40290 14900 40375
rect 14956 40374 14996 40459
rect 15052 40265 15092 40636
rect 15148 40508 15188 40720
rect 15148 40468 15284 40508
rect 15147 40340 15189 40349
rect 15147 40300 15148 40340
rect 15188 40300 15189 40340
rect 15147 40291 15189 40300
rect 15051 40256 15093 40265
rect 15051 40216 15052 40256
rect 15092 40216 15093 40256
rect 15051 40207 15093 40216
rect 14955 40172 14997 40181
rect 14955 40132 14956 40172
rect 14996 40132 14997 40172
rect 14955 40123 14997 40132
rect 14859 39752 14901 39761
rect 14859 39712 14860 39752
rect 14900 39712 14901 39752
rect 14859 39703 14901 39712
rect 14860 39618 14900 39703
rect 14956 38996 14996 40123
rect 15051 40088 15093 40097
rect 15051 40048 15052 40088
rect 15092 40048 15093 40088
rect 15051 40039 15093 40048
rect 14860 38912 14900 38921
rect 14860 37661 14900 38872
rect 14956 38753 14996 38956
rect 14955 38744 14997 38753
rect 14955 38704 14956 38744
rect 14996 38704 14997 38744
rect 14955 38695 14997 38704
rect 14859 37652 14901 37661
rect 14859 37612 14860 37652
rect 14900 37612 14901 37652
rect 14859 37603 14901 37612
rect 14956 36812 14996 36821
rect 14764 36772 14900 36812
rect 14764 36714 14804 36723
rect 14572 35300 14612 35309
rect 14764 35300 14804 36674
rect 14860 35300 14900 36772
rect 14956 35981 14996 36772
rect 14955 35972 14997 35981
rect 14955 35932 14956 35972
rect 14996 35932 14997 35972
rect 14955 35923 14997 35932
rect 14612 35260 14804 35300
rect 14857 35260 14900 35300
rect 14572 35251 14612 35260
rect 14857 35132 14897 35260
rect 14956 35216 14996 35225
rect 14857 35092 14900 35132
rect 14476 34504 14708 34544
rect 13996 34376 14036 34385
rect 14476 34376 14516 34385
rect 14036 34336 14132 34376
rect 13996 34327 14036 34336
rect 13995 34208 14037 34217
rect 13995 34168 13996 34208
rect 14036 34168 14037 34208
rect 13995 34159 14037 34168
rect 13996 32201 14036 34159
rect 14092 34133 14132 34336
rect 14188 34292 14228 34301
rect 14476 34292 14516 34336
rect 14228 34252 14516 34292
rect 14572 34376 14612 34385
rect 14188 34243 14228 34252
rect 14572 34217 14612 34336
rect 14571 34208 14613 34217
rect 14571 34168 14572 34208
rect 14612 34168 14613 34208
rect 14571 34159 14613 34168
rect 14091 34124 14133 34133
rect 14091 34084 14092 34124
rect 14132 34084 14133 34124
rect 14091 34075 14133 34084
rect 14091 33956 14133 33965
rect 14091 33916 14092 33956
rect 14132 33916 14133 33956
rect 14091 33907 14133 33916
rect 14092 33704 14132 33907
rect 14092 33293 14132 33664
rect 14476 33704 14516 33715
rect 14476 33629 14516 33664
rect 14475 33620 14517 33629
rect 14475 33580 14476 33620
rect 14516 33580 14517 33620
rect 14475 33571 14517 33580
rect 14283 33452 14325 33461
rect 14668 33452 14708 34504
rect 14283 33412 14284 33452
rect 14324 33412 14325 33452
rect 14283 33403 14325 33412
rect 14476 33412 14708 33452
rect 14284 33318 14324 33403
rect 14091 33284 14133 33293
rect 14091 33244 14092 33284
rect 14132 33244 14133 33284
rect 14091 33235 14133 33244
rect 13995 32192 14037 32201
rect 13995 32152 13996 32192
rect 14036 32152 14037 32192
rect 13995 32143 14037 32152
rect 14283 32192 14325 32201
rect 14283 32152 14284 32192
rect 14324 32152 14325 32192
rect 14283 32143 14325 32152
rect 14284 32058 14324 32143
rect 14379 32108 14421 32117
rect 14379 32068 14380 32108
rect 14420 32068 14421 32108
rect 14379 32059 14421 32068
rect 13900 29968 14132 30008
rect 13419 28580 13461 28589
rect 13419 28540 13420 28580
rect 13460 28540 13461 28580
rect 13419 28531 13461 28540
rect 13612 27908 13652 29968
rect 13707 29840 13749 29849
rect 13707 29800 13708 29840
rect 13748 29800 13749 29840
rect 13707 29791 13749 29800
rect 13804 29840 13844 29849
rect 13708 29706 13748 29791
rect 13804 29093 13844 29800
rect 13995 29840 14037 29849
rect 13995 29800 13996 29840
rect 14036 29800 14037 29840
rect 13995 29791 14037 29800
rect 13899 29756 13941 29765
rect 13899 29716 13900 29756
rect 13940 29716 13941 29756
rect 13899 29707 13941 29716
rect 13900 29622 13940 29707
rect 13996 29706 14036 29791
rect 14092 29504 14132 29968
rect 13900 29464 14132 29504
rect 14284 29840 14324 29849
rect 13803 29084 13845 29093
rect 13803 29044 13804 29084
rect 13844 29044 13845 29084
rect 13803 29035 13845 29044
rect 13804 28337 13844 28422
rect 13803 28328 13845 28337
rect 13803 28288 13804 28328
rect 13844 28288 13845 28328
rect 13803 28279 13845 28288
rect 13612 27868 13844 27908
rect 13324 27784 13748 27824
rect 13324 27656 13364 27667
rect 13324 27581 13364 27616
rect 13323 27572 13365 27581
rect 13323 27532 13324 27572
rect 13364 27532 13365 27572
rect 13323 27523 13365 27532
rect 13516 27404 13556 27413
rect 13324 26816 13364 26825
rect 13324 26405 13364 26776
rect 13420 26816 13460 26825
rect 13420 26489 13460 26776
rect 13516 26657 13556 27364
rect 13515 26648 13557 26657
rect 13515 26608 13516 26648
rect 13556 26608 13557 26648
rect 13515 26599 13557 26608
rect 13708 26489 13748 27784
rect 13804 26816 13844 27868
rect 13900 26984 13940 29464
rect 14091 29336 14133 29345
rect 14091 29296 14092 29336
rect 14132 29296 14133 29336
rect 14091 29287 14133 29296
rect 14188 29336 14228 29345
rect 14284 29336 14324 29800
rect 14228 29296 14324 29336
rect 14380 29840 14420 32059
rect 14188 29287 14228 29296
rect 13995 29252 14037 29261
rect 13995 29212 13996 29252
rect 14036 29212 14037 29252
rect 13995 29203 14037 29212
rect 13996 29168 14036 29203
rect 13996 29117 14036 29128
rect 14092 29000 14132 29287
rect 14092 28960 14324 29000
rect 13995 28328 14037 28337
rect 13995 28288 13996 28328
rect 14036 28288 14037 28328
rect 13995 28279 14037 28288
rect 13996 28194 14036 28279
rect 13995 27656 14037 27665
rect 13995 27616 13996 27656
rect 14036 27616 14037 27656
rect 13995 27607 14037 27616
rect 13996 27522 14036 27607
rect 13900 26944 14132 26984
rect 13900 26816 13940 26825
rect 13804 26776 13900 26816
rect 13940 26776 14036 26816
rect 13900 26767 13940 26776
rect 13899 26648 13941 26657
rect 13899 26608 13900 26648
rect 13940 26608 13941 26648
rect 13899 26599 13941 26608
rect 13803 26564 13845 26573
rect 13803 26524 13804 26564
rect 13844 26524 13845 26564
rect 13803 26515 13845 26524
rect 13419 26480 13461 26489
rect 13419 26440 13420 26480
rect 13460 26440 13461 26480
rect 13419 26431 13461 26440
rect 13707 26480 13749 26489
rect 13707 26440 13708 26480
rect 13748 26440 13749 26480
rect 13707 26431 13749 26440
rect 13323 26396 13365 26405
rect 13323 26356 13324 26396
rect 13364 26356 13365 26396
rect 13323 26347 13365 26356
rect 13420 26144 13460 26153
rect 13324 26104 13420 26144
rect 13324 25892 13364 26104
rect 13420 26095 13460 26104
rect 13611 26144 13653 26153
rect 13611 26104 13612 26144
rect 13652 26104 13653 26144
rect 13611 26095 13653 26104
rect 13804 26144 13844 26515
rect 13804 26095 13844 26104
rect 13612 26010 13652 26095
rect 13612 25892 13652 25901
rect 13324 25852 13556 25892
rect 13323 25724 13365 25733
rect 13323 25684 13324 25724
rect 13364 25684 13365 25724
rect 13323 25675 13365 25684
rect 13227 25136 13269 25145
rect 13227 25096 13228 25136
rect 13268 25096 13269 25136
rect 13227 25087 13269 25096
rect 12939 24968 12981 24977
rect 12939 24928 12940 24968
rect 12980 24928 12981 24968
rect 12939 24919 12981 24928
rect 13035 24800 13077 24809
rect 13035 24760 13036 24800
rect 13076 24760 13077 24800
rect 13035 24751 13077 24760
rect 13227 24800 13269 24809
rect 13227 24760 13228 24800
rect 13268 24760 13269 24800
rect 13227 24751 13269 24760
rect 13324 24800 13364 25675
rect 13420 25313 13460 25398
rect 13516 25397 13556 25852
rect 13515 25388 13557 25397
rect 13515 25348 13516 25388
rect 13556 25348 13557 25388
rect 13515 25339 13557 25348
rect 13419 25304 13461 25313
rect 13419 25264 13420 25304
rect 13460 25264 13461 25304
rect 13419 25255 13461 25264
rect 13516 25304 13556 25339
rect 13516 25253 13556 25264
rect 13612 25136 13652 25852
rect 13803 25388 13845 25397
rect 13803 25348 13804 25388
rect 13844 25348 13845 25388
rect 13803 25339 13845 25348
rect 13324 24751 13364 24760
rect 13420 25096 13652 25136
rect 13036 24666 13076 24751
rect 12844 24632 12884 24641
rect 12844 24473 12884 24592
rect 13228 24632 13268 24751
rect 13228 24583 13268 24592
rect 13420 24632 13460 25096
rect 13804 24800 13844 25339
rect 13900 24800 13940 26599
rect 13996 26153 14036 26776
rect 14092 26732 14132 26944
rect 14284 26816 14324 28960
rect 14380 28085 14420 29800
rect 14476 29345 14516 33412
rect 14571 33284 14613 33293
rect 14571 33244 14572 33284
rect 14612 33244 14613 33284
rect 14571 33235 14613 33244
rect 14572 32864 14612 33235
rect 14860 33032 14900 35092
rect 14956 35057 14996 35176
rect 14955 35048 14997 35057
rect 14955 35008 14956 35048
rect 14996 35008 14997 35048
rect 14955 34999 14997 35008
rect 15052 34628 15092 40039
rect 15148 37829 15188 40291
rect 15244 40181 15284 40468
rect 15436 40424 15476 40433
rect 15340 40384 15436 40424
rect 15243 40172 15285 40181
rect 15243 40132 15244 40172
rect 15284 40132 15285 40172
rect 15243 40123 15285 40132
rect 15340 38165 15380 40384
rect 15436 40375 15476 40384
rect 15531 39920 15573 39929
rect 15531 39880 15532 39920
rect 15572 39880 15573 39920
rect 15531 39871 15573 39880
rect 15436 38912 15476 38921
rect 15339 38156 15381 38165
rect 15339 38116 15340 38156
rect 15380 38116 15381 38156
rect 15339 38107 15381 38116
rect 15147 37820 15189 37829
rect 15147 37780 15148 37820
rect 15188 37780 15189 37820
rect 15147 37771 15189 37780
rect 15436 37745 15476 38872
rect 15435 37736 15477 37745
rect 15435 37696 15436 37736
rect 15476 37696 15477 37736
rect 15435 37687 15477 37696
rect 15435 37568 15477 37577
rect 15435 37528 15436 37568
rect 15476 37528 15477 37568
rect 15435 37519 15477 37528
rect 15340 37400 15380 37409
rect 15148 37360 15340 37400
rect 15148 36140 15188 37360
rect 15340 37351 15380 37360
rect 15436 37400 15476 37519
rect 15436 36737 15476 37360
rect 15244 36728 15284 36737
rect 15244 36149 15284 36688
rect 15340 36728 15380 36737
rect 15340 36569 15380 36688
rect 15435 36728 15477 36737
rect 15435 36688 15436 36728
rect 15476 36688 15477 36728
rect 15435 36679 15477 36688
rect 15339 36560 15381 36569
rect 15339 36520 15340 36560
rect 15380 36520 15381 36560
rect 15339 36511 15381 36520
rect 15148 36091 15188 36100
rect 15243 36140 15285 36149
rect 15243 36100 15244 36140
rect 15284 36100 15285 36140
rect 15243 36091 15285 36100
rect 15340 35888 15380 35897
rect 15244 35848 15340 35888
rect 15244 35393 15284 35848
rect 15340 35839 15380 35848
rect 15243 35384 15285 35393
rect 15243 35344 15244 35384
rect 15284 35344 15285 35384
rect 15243 35335 15285 35344
rect 15052 34588 15188 34628
rect 15051 34460 15093 34469
rect 15051 34420 15052 34460
rect 15092 34420 15093 34460
rect 15051 34411 15093 34420
rect 14955 34376 14997 34385
rect 14955 34336 14956 34376
rect 14996 34336 14997 34376
rect 14955 34327 14997 34336
rect 14956 33293 14996 34327
rect 15052 34326 15092 34411
rect 15148 34208 15188 34588
rect 15052 34168 15188 34208
rect 14955 33284 14997 33293
rect 14955 33244 14956 33284
rect 14996 33244 14997 33284
rect 14955 33235 14997 33244
rect 14860 32992 14996 33032
rect 14860 32885 14900 32894
rect 14572 32845 14860 32864
rect 14572 32824 14900 32845
rect 14572 31352 14612 32824
rect 14956 32780 14996 32992
rect 15052 32864 15092 34168
rect 15244 33965 15284 35335
rect 15435 35300 15477 35309
rect 15435 35260 15436 35300
rect 15476 35260 15477 35300
rect 15435 35251 15477 35260
rect 15436 34553 15476 35251
rect 15435 34544 15477 34553
rect 15435 34504 15436 34544
rect 15476 34504 15477 34544
rect 15435 34495 15477 34504
rect 15532 34376 15572 39871
rect 15628 35309 15668 41719
rect 15724 39500 15764 41812
rect 16395 41803 16437 41812
rect 16107 41768 16149 41777
rect 16300 41768 16340 41777
rect 16107 41728 16108 41768
rect 16148 41728 16149 41768
rect 16107 41719 16149 41728
rect 16204 41728 16300 41768
rect 16108 41634 16148 41719
rect 16204 41516 16244 41728
rect 16300 41719 16340 41728
rect 16012 41476 16244 41516
rect 16012 41264 16052 41476
rect 16396 41432 16436 41803
rect 16492 41802 16532 41887
rect 16108 41348 16148 41357
rect 16148 41308 16244 41348
rect 16108 41299 16148 41308
rect 15964 41254 16052 41264
rect 16004 41224 16052 41254
rect 15964 41205 16004 41214
rect 15819 40592 15861 40601
rect 15819 40552 15820 40592
rect 15860 40552 15861 40592
rect 15819 40543 15861 40552
rect 15820 39677 15860 40543
rect 16011 40508 16053 40517
rect 16011 40468 16012 40508
rect 16052 40468 16053 40508
rect 16011 40459 16053 40468
rect 15916 40433 15956 40438
rect 15915 40429 15957 40433
rect 15915 40384 15916 40429
rect 15956 40384 15957 40429
rect 15915 40375 15957 40384
rect 15916 40294 15956 40375
rect 15819 39668 15861 39677
rect 15819 39628 15820 39668
rect 15860 39628 15861 39668
rect 15819 39619 15861 39628
rect 15724 39460 15860 39500
rect 15723 38744 15765 38753
rect 15723 38704 15724 38744
rect 15764 38704 15765 38744
rect 15723 38695 15765 38704
rect 15724 37232 15764 38695
rect 15820 37913 15860 39460
rect 16012 39080 16052 40459
rect 16108 40256 16148 40265
rect 16108 39929 16148 40216
rect 16107 39920 16149 39929
rect 16107 39880 16108 39920
rect 16148 39880 16149 39920
rect 16107 39871 16149 39880
rect 16108 39752 16148 39763
rect 16108 39677 16148 39712
rect 16107 39668 16149 39677
rect 16107 39628 16108 39668
rect 16148 39628 16149 39668
rect 16107 39619 16149 39628
rect 16012 39040 16148 39080
rect 15964 38921 16004 38930
rect 16004 38881 16052 38912
rect 15964 38872 16052 38881
rect 15915 38576 15957 38585
rect 15915 38536 15916 38576
rect 15956 38536 15957 38576
rect 15915 38527 15957 38536
rect 15916 38240 15956 38527
rect 16012 38408 16052 38872
rect 16108 38828 16148 39040
rect 16108 38585 16148 38788
rect 16107 38576 16149 38585
rect 16107 38536 16108 38576
rect 16148 38536 16149 38576
rect 16107 38527 16149 38536
rect 16108 38408 16148 38417
rect 16012 38368 16108 38408
rect 16108 38359 16148 38368
rect 16204 38240 16244 41308
rect 16396 40592 16436 41392
rect 16396 39920 16436 40552
rect 16396 39871 16436 39880
rect 16300 39584 16340 39593
rect 16300 39080 16340 39544
rect 16300 38753 16340 39040
rect 16299 38744 16341 38753
rect 16299 38704 16300 38744
rect 16340 38704 16341 38744
rect 16299 38695 16341 38704
rect 16491 38744 16533 38753
rect 16491 38704 16492 38744
rect 16532 38704 16533 38744
rect 16491 38695 16533 38704
rect 16299 38576 16341 38585
rect 16299 38536 16300 38576
rect 16340 38536 16341 38576
rect 16299 38527 16341 38536
rect 15916 38191 15956 38200
rect 16012 38200 16244 38240
rect 15819 37904 15861 37913
rect 15819 37864 15820 37904
rect 15860 37864 15861 37904
rect 15819 37855 15861 37864
rect 15819 37736 15861 37745
rect 15819 37696 15820 37736
rect 15860 37696 15861 37736
rect 15819 37687 15861 37696
rect 15820 37484 15860 37687
rect 15915 37652 15957 37661
rect 15915 37612 15916 37652
rect 15956 37612 15957 37652
rect 15915 37603 15957 37612
rect 15820 37435 15860 37444
rect 15916 37484 15956 37603
rect 15724 37192 15860 37232
rect 15723 36728 15765 36737
rect 15723 36688 15724 36728
rect 15764 36688 15765 36728
rect 15723 36679 15765 36688
rect 15820 36728 15860 37192
rect 15820 36679 15860 36688
rect 15724 36594 15764 36679
rect 15916 36653 15956 37444
rect 15915 36644 15957 36653
rect 15915 36604 15916 36644
rect 15956 36604 15957 36644
rect 15915 36595 15957 36604
rect 15723 36476 15765 36485
rect 15723 36436 15724 36476
rect 15764 36436 15765 36476
rect 15723 36427 15765 36436
rect 15627 35300 15669 35309
rect 15627 35260 15628 35300
rect 15668 35260 15669 35300
rect 15627 35251 15669 35260
rect 15627 35048 15669 35057
rect 15627 35008 15628 35048
rect 15668 35008 15669 35048
rect 15627 34999 15669 35008
rect 15436 34336 15532 34376
rect 15243 33956 15285 33965
rect 15243 33916 15244 33956
rect 15284 33916 15285 33956
rect 15243 33907 15285 33916
rect 15052 32824 15188 32864
rect 14572 31277 14612 31312
rect 14668 32740 14996 32780
rect 14571 31268 14613 31277
rect 14571 31228 14572 31268
rect 14612 31228 14613 31268
rect 14571 31219 14613 31228
rect 14572 30689 14612 31219
rect 14571 30680 14613 30689
rect 14571 30640 14572 30680
rect 14612 30640 14613 30680
rect 14571 30631 14613 30640
rect 14475 29336 14517 29345
rect 14475 29296 14476 29336
rect 14516 29296 14517 29336
rect 14475 29287 14517 29296
rect 14476 29168 14516 29177
rect 14379 28076 14421 28085
rect 14379 28036 14380 28076
rect 14420 28036 14421 28076
rect 14379 28027 14421 28036
rect 14476 27917 14516 29128
rect 14475 27908 14517 27917
rect 14283 26776 14324 26816
rect 14380 27868 14476 27908
rect 14516 27868 14517 27908
rect 14380 26830 14420 27868
rect 14475 27859 14517 27868
rect 14571 27488 14613 27497
rect 14571 27448 14572 27488
rect 14612 27448 14613 27488
rect 14571 27439 14613 27448
rect 14092 26692 14228 26732
rect 14091 26564 14133 26573
rect 14091 26524 14092 26564
rect 14132 26524 14133 26564
rect 14091 26515 14133 26524
rect 13995 26144 14037 26153
rect 13995 26104 13996 26144
rect 14036 26104 14037 26144
rect 13995 26095 14037 26104
rect 13996 25313 14036 25398
rect 14092 25397 14132 26515
rect 14091 25388 14133 25397
rect 14091 25348 14092 25388
rect 14132 25348 14133 25388
rect 14091 25339 14133 25348
rect 13995 25304 14037 25313
rect 13995 25264 13996 25304
rect 14036 25264 14037 25304
rect 13995 25255 14037 25264
rect 14091 25136 14133 25145
rect 14091 25096 14092 25136
rect 14132 25096 14133 25136
rect 14091 25087 14133 25096
rect 13804 24751 13844 24760
rect 13899 24760 13940 24800
rect 13899 24716 13939 24760
rect 13899 24676 13940 24716
rect 13900 24653 13940 24676
rect 13420 24583 13460 24592
rect 13515 24632 13557 24641
rect 13515 24592 13516 24632
rect 13556 24592 13557 24632
rect 13900 24604 13940 24613
rect 13996 24632 14036 24641
rect 13515 24583 13557 24592
rect 13516 24498 13556 24583
rect 13996 24548 14036 24592
rect 14092 24632 14132 25087
rect 14092 24583 14132 24592
rect 13900 24508 14036 24548
rect 12843 24464 12885 24473
rect 12843 24424 12844 24464
rect 12884 24424 12980 24464
rect 12843 24415 12885 24424
rect 12844 23213 12884 23298
rect 12940 23288 12980 24424
rect 13515 24212 13557 24221
rect 13515 24172 13516 24212
rect 13556 24172 13557 24212
rect 13515 24163 13557 24172
rect 13227 23960 13269 23969
rect 13227 23920 13228 23960
rect 13268 23920 13269 23960
rect 13227 23911 13269 23920
rect 13228 23792 13268 23911
rect 13228 23743 13268 23752
rect 12933 23248 12980 23288
rect 12843 23204 12885 23213
rect 12843 23164 12844 23204
rect 12884 23164 12885 23204
rect 12843 23155 12885 23164
rect 12933 23120 12973 23248
rect 13131 23204 13173 23213
rect 13131 23164 13132 23204
rect 13172 23164 13173 23204
rect 13131 23155 13173 23164
rect 13132 23120 13172 23155
rect 12933 23080 12980 23120
rect 12747 22616 12789 22625
rect 12747 22576 12748 22616
rect 12788 22576 12789 22616
rect 12747 22567 12789 22576
rect 12940 22541 12980 23080
rect 13132 23069 13172 23080
rect 13228 23120 13268 23129
rect 13035 22952 13077 22961
rect 13228 22952 13268 23080
rect 13419 23120 13461 23129
rect 13419 23080 13420 23120
rect 13460 23080 13461 23120
rect 13419 23071 13461 23080
rect 13035 22912 13036 22952
rect 13076 22912 13268 22952
rect 13035 22903 13077 22912
rect 12555 22532 12597 22541
rect 12555 22492 12556 22532
rect 12596 22492 12597 22532
rect 12555 22483 12597 22492
rect 12939 22532 12981 22541
rect 12939 22492 12940 22532
rect 12980 22492 12981 22532
rect 12939 22483 12981 22492
rect 12556 21776 12596 22483
rect 12651 22364 12693 22373
rect 13036 22364 13076 22903
rect 13420 22793 13460 23071
rect 13516 22868 13556 24163
rect 13900 23885 13940 24508
rect 13995 24380 14037 24389
rect 13995 24340 13996 24380
rect 14036 24340 14037 24380
rect 13995 24331 14037 24340
rect 13611 23876 13653 23885
rect 13611 23836 13612 23876
rect 13652 23836 13653 23876
rect 13611 23827 13653 23836
rect 13899 23876 13941 23885
rect 13899 23836 13900 23876
rect 13940 23836 13941 23876
rect 13899 23827 13941 23836
rect 13612 23129 13652 23827
rect 13996 23708 14036 24331
rect 14091 24296 14133 24305
rect 14091 24256 14092 24296
rect 14132 24256 14133 24296
rect 14091 24247 14133 24256
rect 13900 23668 14036 23708
rect 13611 23120 13653 23129
rect 13611 23080 13612 23120
rect 13652 23080 13653 23120
rect 13611 23071 13653 23080
rect 13612 22986 13652 23071
rect 13708 23036 13748 23045
rect 13708 22868 13748 22996
rect 13516 22828 13748 22868
rect 13227 22784 13269 22793
rect 13227 22744 13228 22784
rect 13268 22744 13269 22784
rect 13227 22735 13269 22744
rect 13419 22784 13461 22793
rect 13419 22744 13420 22784
rect 13460 22744 13461 22784
rect 13419 22735 13461 22744
rect 13131 22616 13173 22625
rect 13131 22576 13132 22616
rect 13172 22576 13173 22616
rect 13131 22567 13173 22576
rect 12651 22324 12652 22364
rect 12692 22324 12693 22364
rect 12651 22315 12693 22324
rect 12940 22324 13076 22364
rect 12652 22280 12692 22315
rect 12748 22299 12788 22308
rect 12940 22285 12980 22324
rect 12788 22259 12980 22285
rect 13132 22280 13172 22567
rect 13228 22364 13268 22735
rect 13228 22315 13268 22324
rect 12748 22245 12980 22259
rect 12652 22229 12692 22240
rect 12940 21944 12980 22245
rect 12748 21904 12980 21944
rect 13036 22240 13132 22280
rect 12556 21736 12692 21776
rect 12555 21608 12597 21617
rect 12555 21568 12556 21608
rect 12596 21568 12597 21608
rect 12555 21559 12597 21568
rect 12556 21474 12596 21559
rect 12364 20140 12500 20180
rect 12652 20768 12692 21736
rect 12364 19433 12404 20140
rect 12363 19424 12405 19433
rect 12363 19384 12364 19424
rect 12404 19384 12405 19424
rect 12363 19375 12405 19384
rect 12555 19256 12597 19265
rect 12555 19216 12556 19256
rect 12596 19216 12597 19256
rect 12555 19207 12597 19216
rect 12267 18920 12309 18929
rect 12267 18880 12268 18920
rect 12308 18880 12309 18920
rect 12267 18871 12309 18880
rect 12171 15056 12213 15065
rect 12171 15016 12172 15056
rect 12212 15016 12213 15056
rect 12171 15007 12213 15016
rect 12075 14636 12117 14645
rect 12075 14596 12076 14636
rect 12116 14596 12117 14636
rect 12075 14587 12117 14596
rect 12076 14502 12116 14587
rect 12171 14384 12213 14393
rect 12171 14344 12172 14384
rect 12212 14344 12213 14384
rect 12171 14335 12213 14344
rect 12075 13208 12117 13217
rect 12075 13168 12076 13208
rect 12116 13168 12117 13208
rect 12075 13159 12117 13168
rect 11924 12496 12020 12536
rect 11787 12116 11829 12125
rect 11787 12076 11788 12116
rect 11828 12076 11829 12116
rect 11787 12067 11829 12076
rect 11691 11108 11733 11117
rect 11691 11068 11692 11108
rect 11732 11068 11733 11108
rect 11691 11059 11733 11068
rect 11595 11024 11637 11033
rect 11595 10984 11596 11024
rect 11636 10984 11637 11024
rect 11595 10975 11637 10984
rect 11596 10697 11636 10975
rect 11595 10688 11637 10697
rect 11595 10648 11596 10688
rect 11636 10648 11637 10688
rect 11595 10639 11637 10648
rect 11595 10436 11637 10445
rect 11595 10396 11596 10436
rect 11636 10396 11637 10436
rect 11595 10387 11637 10396
rect 11116 7951 11156 7960
rect 11404 8044 11540 8084
rect 10923 7496 10965 7505
rect 10923 7456 10924 7496
rect 10964 7456 10965 7496
rect 10923 7447 10965 7456
rect 10923 7160 10965 7169
rect 10923 7120 10924 7160
rect 10964 7120 10965 7160
rect 10923 7111 10965 7120
rect 10924 7026 10964 7111
rect 11404 2708 11444 8044
rect 11499 7916 11541 7925
rect 11499 7876 11500 7916
rect 11540 7876 11541 7916
rect 11499 7867 11541 7876
rect 11596 7916 11636 10387
rect 11692 9680 11732 11059
rect 11788 10940 11828 12067
rect 11884 11957 11924 12496
rect 12076 12452 12116 13159
rect 11980 12412 12116 12452
rect 11883 11948 11925 11957
rect 11883 11908 11884 11948
rect 11924 11908 11925 11948
rect 11883 11899 11925 11908
rect 11884 11024 11924 11033
rect 11980 11024 12020 12412
rect 12075 12284 12117 12293
rect 12075 12244 12076 12284
rect 12116 12244 12117 12284
rect 12075 12235 12117 12244
rect 12076 11696 12116 12235
rect 12172 11873 12212 14335
rect 12268 12461 12308 18871
rect 12556 18584 12596 19207
rect 12652 19097 12692 20728
rect 12651 19088 12693 19097
rect 12651 19048 12652 19088
rect 12692 19048 12693 19088
rect 12651 19039 12693 19048
rect 12652 18584 12692 18593
rect 12556 18544 12652 18584
rect 12556 18425 12596 18544
rect 12652 18535 12692 18544
rect 12555 18416 12597 18425
rect 12555 18376 12556 18416
rect 12596 18376 12597 18416
rect 12555 18367 12597 18376
rect 12556 17828 12596 18367
rect 12556 17788 12692 17828
rect 12459 17240 12501 17249
rect 12459 17200 12460 17240
rect 12500 17200 12501 17240
rect 12459 17191 12501 17200
rect 12363 15056 12405 15065
rect 12363 15016 12364 15056
rect 12404 15016 12405 15056
rect 12363 15007 12405 15016
rect 12364 13973 12404 15007
rect 12363 13964 12405 13973
rect 12363 13924 12364 13964
rect 12404 13924 12405 13964
rect 12363 13915 12405 13924
rect 12364 12522 12404 12531
rect 12267 12452 12309 12461
rect 12267 12412 12268 12452
rect 12308 12412 12309 12452
rect 12267 12403 12309 12412
rect 12268 11948 12308 11957
rect 12364 11948 12404 12482
rect 12308 11908 12404 11948
rect 12268 11899 12308 11908
rect 12171 11864 12213 11873
rect 12171 11824 12172 11864
rect 12212 11824 12213 11864
rect 12171 11815 12213 11824
rect 12363 11780 12405 11789
rect 12363 11740 12364 11780
rect 12404 11740 12405 11780
rect 12363 11731 12405 11740
rect 12076 11621 12116 11656
rect 12171 11696 12213 11705
rect 12171 11656 12172 11696
rect 12212 11656 12213 11696
rect 12171 11647 12213 11656
rect 12075 11612 12117 11621
rect 12075 11572 12076 11612
rect 12116 11572 12117 11612
rect 12075 11563 12117 11572
rect 11924 10984 12020 11024
rect 11884 10975 11924 10984
rect 11788 10856 11828 10900
rect 11788 10816 12116 10856
rect 11979 10688 12021 10697
rect 11979 10648 11980 10688
rect 12020 10648 12021 10688
rect 11979 10639 12021 10648
rect 11883 10352 11925 10361
rect 11883 10312 11884 10352
rect 11924 10312 11925 10352
rect 11883 10303 11925 10312
rect 11692 9640 11828 9680
rect 11691 9512 11733 9521
rect 11691 9472 11692 9512
rect 11732 9472 11733 9512
rect 11691 9463 11733 9472
rect 11692 9378 11732 9463
rect 11788 9008 11828 9640
rect 11692 8968 11828 9008
rect 11692 8681 11732 8968
rect 11787 8840 11829 8849
rect 11787 8800 11788 8840
rect 11828 8800 11829 8840
rect 11787 8791 11829 8800
rect 11691 8672 11733 8681
rect 11691 8632 11692 8672
rect 11732 8632 11733 8672
rect 11691 8623 11733 8632
rect 11691 8084 11733 8093
rect 11691 8044 11692 8084
rect 11732 8044 11733 8084
rect 11691 8035 11733 8044
rect 11500 6497 11540 7867
rect 11499 6488 11541 6497
rect 11499 6448 11500 6488
rect 11540 6448 11541 6488
rect 11499 6439 11541 6448
rect 11499 6320 11541 6329
rect 11499 6280 11500 6320
rect 11540 6280 11541 6320
rect 11499 6271 11541 6280
rect 11500 6186 11540 6271
rect 11596 6236 11636 7876
rect 11692 6404 11732 8035
rect 11788 7925 11828 8791
rect 11787 7916 11829 7925
rect 11787 7876 11788 7916
rect 11828 7876 11829 7916
rect 11787 7867 11829 7876
rect 11692 6355 11732 6364
rect 11596 6196 11828 6236
rect 11499 6068 11541 6077
rect 11499 6028 11500 6068
rect 11540 6028 11541 6068
rect 11499 6019 11541 6028
rect 11404 2659 11444 2668
rect 10348 2500 10484 2540
rect 10636 2500 11060 2540
rect 10156 1744 10292 1784
rect 9964 1700 10004 1709
rect 9867 1196 9909 1205
rect 9867 1156 9868 1196
rect 9908 1156 9909 1196
rect 9867 1147 9909 1156
rect 9964 869 10004 1660
rect 10059 1700 10101 1709
rect 10059 1660 10060 1700
rect 10100 1660 10101 1700
rect 10059 1651 10101 1660
rect 9963 860 10005 869
rect 9963 820 9964 860
rect 10004 820 10005 860
rect 9963 811 10005 820
rect 9867 776 9909 785
rect 9867 736 9868 776
rect 9908 736 9909 776
rect 9867 727 9909 736
rect 9771 272 9813 281
rect 9771 232 9772 272
rect 9812 232 9813 272
rect 9771 223 9813 232
rect 9868 80 9908 727
rect 10060 80 10100 1651
rect 10156 608 10196 1744
rect 10348 1700 10388 1709
rect 10252 1660 10348 1700
rect 10252 785 10292 1660
rect 10348 1651 10388 1660
rect 10347 1196 10389 1205
rect 10347 1156 10348 1196
rect 10388 1156 10389 1196
rect 10347 1147 10389 1156
rect 10348 1062 10388 1147
rect 10251 776 10293 785
rect 10251 736 10252 776
rect 10292 736 10293 776
rect 10251 727 10293 736
rect 10156 568 10292 608
rect 10252 80 10292 568
rect 10444 80 10484 2500
rect 10539 1868 10581 1877
rect 10539 1828 10540 1868
rect 10580 1828 10581 1868
rect 10539 1819 10581 1828
rect 10923 1868 10965 1877
rect 10923 1828 10924 1868
rect 10964 1828 10965 1868
rect 10923 1819 10965 1828
rect 10540 1734 10580 1819
rect 10924 1734 10964 1819
rect 10732 1700 10772 1709
rect 10732 1373 10772 1660
rect 10827 1448 10869 1457
rect 10827 1408 10828 1448
rect 10868 1408 10869 1448
rect 10827 1399 10869 1408
rect 10731 1364 10773 1373
rect 10731 1324 10732 1364
rect 10772 1324 10773 1364
rect 10731 1315 10773 1324
rect 10539 944 10581 953
rect 10539 904 10540 944
rect 10580 904 10581 944
rect 10539 895 10581 904
rect 10540 810 10580 895
rect 10635 860 10677 869
rect 10635 820 10636 860
rect 10676 820 10677 860
rect 10635 811 10677 820
rect 10636 80 10676 811
rect 10828 80 10868 1399
rect 11020 1196 11060 2500
rect 11500 1868 11540 6019
rect 11788 2540 11828 6196
rect 11884 6077 11924 10303
rect 11883 6068 11925 6077
rect 11883 6028 11884 6068
rect 11924 6028 11925 6068
rect 11883 6019 11925 6028
rect 11980 2801 12020 10639
rect 12076 8429 12116 10816
rect 12075 8420 12117 8429
rect 12075 8380 12076 8420
rect 12116 8380 12117 8420
rect 12075 8371 12117 8380
rect 12076 8000 12116 8009
rect 12172 8000 12212 11647
rect 12364 11024 12404 11731
rect 12364 10975 12404 10984
rect 12460 9521 12500 17191
rect 12556 17072 12596 17788
rect 12652 17786 12692 17788
rect 12652 17737 12692 17746
rect 12748 17576 12788 21904
rect 12940 20945 12980 21030
rect 12939 20936 12981 20945
rect 12939 20896 12940 20936
rect 12980 20896 12981 20936
rect 12939 20887 12981 20896
rect 12844 20768 12884 20777
rect 12844 20105 12884 20728
rect 12940 20768 12980 20777
rect 12843 20096 12885 20105
rect 12843 20056 12844 20096
rect 12884 20056 12885 20096
rect 12843 20047 12885 20056
rect 12843 19760 12885 19769
rect 12843 19720 12844 19760
rect 12884 19720 12885 19760
rect 12843 19711 12885 19720
rect 12844 19349 12884 19711
rect 12940 19508 12980 20728
rect 13036 20273 13076 22240
rect 13132 22231 13172 22240
rect 13131 22112 13173 22121
rect 13131 22072 13132 22112
rect 13172 22072 13173 22112
rect 13131 22063 13173 22072
rect 13132 20936 13172 22063
rect 13132 20777 13172 20896
rect 13323 20936 13365 20945
rect 13323 20896 13324 20936
rect 13364 20896 13365 20936
rect 13323 20887 13365 20896
rect 13131 20768 13173 20777
rect 13131 20728 13132 20768
rect 13172 20728 13173 20768
rect 13131 20719 13173 20728
rect 13131 20432 13173 20441
rect 13131 20392 13132 20432
rect 13172 20392 13173 20432
rect 13131 20383 13173 20392
rect 13035 20264 13077 20273
rect 13035 20224 13036 20264
rect 13076 20224 13077 20264
rect 13035 20215 13077 20224
rect 13036 20096 13076 20105
rect 13036 19769 13076 20056
rect 13035 19760 13077 19769
rect 13035 19720 13036 19760
rect 13076 19720 13077 19760
rect 13035 19711 13077 19720
rect 13132 19676 13172 20383
rect 13228 20264 13268 20273
rect 13228 20105 13268 20224
rect 13227 20096 13269 20105
rect 13227 20056 13228 20096
rect 13268 20056 13269 20096
rect 13227 20047 13269 20056
rect 13228 20045 13268 20047
rect 13132 19636 13268 19676
rect 13132 19508 13172 19517
rect 12940 19468 13132 19508
rect 13132 19459 13172 19468
rect 13228 19433 13268 19636
rect 13227 19424 13269 19433
rect 13227 19384 13228 19424
rect 13268 19384 13269 19424
rect 13227 19375 13269 19384
rect 12843 19340 12885 19349
rect 12843 19300 12844 19340
rect 12884 19300 12980 19340
rect 12843 19291 12885 19300
rect 12940 19256 12980 19300
rect 12940 19207 12980 19216
rect 13324 19256 13364 20887
rect 13419 20768 13461 20777
rect 13419 20728 13420 20768
rect 13460 20728 13461 20768
rect 13419 20719 13461 20728
rect 13420 20634 13460 20719
rect 13516 20096 13556 20105
rect 13516 19937 13556 20056
rect 13515 19928 13557 19937
rect 13515 19888 13516 19928
rect 13556 19888 13557 19928
rect 13515 19879 13557 19888
rect 13612 19760 13652 22828
rect 13708 22280 13748 22289
rect 13708 21953 13748 22240
rect 13707 21944 13749 21953
rect 13707 21904 13708 21944
rect 13748 21904 13749 21944
rect 13707 21895 13749 21904
rect 13804 21608 13844 21617
rect 13804 21365 13844 21568
rect 13803 21356 13845 21365
rect 13803 21316 13804 21356
rect 13844 21316 13845 21356
rect 13803 21307 13845 21316
rect 13804 20441 13844 21307
rect 13803 20432 13845 20441
rect 13803 20392 13804 20432
rect 13844 20392 13845 20432
rect 13803 20383 13845 20392
rect 13900 20180 13940 23668
rect 14092 21869 14132 24247
rect 14188 23297 14228 26692
rect 14283 26648 14323 26776
rect 14380 26732 14420 26790
rect 14572 26732 14612 27439
rect 14380 26692 14516 26732
rect 14283 26608 14324 26648
rect 14284 26480 14324 26608
rect 14284 26440 14420 26480
rect 14283 25220 14325 25229
rect 14283 25180 14284 25220
rect 14324 25180 14325 25220
rect 14283 25171 14325 25180
rect 14284 24632 14324 25171
rect 14284 24583 14324 24592
rect 14187 23288 14229 23297
rect 14187 23248 14188 23288
rect 14228 23248 14229 23288
rect 14187 23239 14229 23248
rect 14188 23120 14228 23129
rect 14228 23080 14324 23120
rect 14188 23071 14228 23080
rect 14188 22285 14228 22294
rect 14091 21860 14133 21869
rect 14091 21820 14092 21860
rect 14132 21820 14133 21860
rect 14188 21860 14228 22245
rect 14284 21953 14324 23080
rect 14380 22289 14420 26440
rect 14476 25145 14516 26692
rect 14572 26683 14612 26692
rect 14571 26480 14613 26489
rect 14571 26440 14572 26480
rect 14612 26440 14613 26480
rect 14571 26431 14613 26440
rect 14475 25136 14517 25145
rect 14475 25096 14476 25136
rect 14516 25096 14517 25136
rect 14475 25087 14517 25096
rect 14475 24632 14517 24641
rect 14475 24592 14476 24632
rect 14516 24592 14517 24632
rect 14475 24583 14517 24592
rect 14572 24632 14612 26431
rect 14572 24583 14612 24592
rect 14476 24498 14516 24583
rect 14668 24212 14708 32740
rect 15052 32696 15092 32705
rect 14860 32656 15052 32696
rect 14860 32192 14900 32656
rect 15052 32647 15092 32656
rect 15148 32528 15188 32824
rect 15052 32488 15188 32528
rect 14812 32182 14900 32192
rect 14852 32152 14900 32182
rect 14956 32276 14996 32285
rect 14812 32133 14852 32142
rect 14763 31520 14805 31529
rect 14763 31480 14764 31520
rect 14804 31480 14805 31520
rect 14763 31471 14805 31480
rect 14764 31386 14804 31471
rect 14763 30848 14805 30857
rect 14956 30848 14996 32236
rect 14763 30808 14764 30848
rect 14804 30808 14805 30848
rect 14763 30799 14805 30808
rect 14860 30808 14996 30848
rect 14764 30714 14804 30799
rect 14860 30185 14900 30808
rect 14956 30680 14996 30689
rect 15052 30680 15092 32488
rect 15147 32192 15189 32201
rect 15147 32152 15148 32192
rect 15188 32152 15189 32192
rect 15147 32143 15189 32152
rect 15244 32192 15284 32201
rect 14996 30640 15092 30680
rect 14859 30176 14901 30185
rect 14859 30136 14860 30176
rect 14900 30136 14901 30176
rect 14859 30127 14901 30136
rect 14859 29924 14901 29933
rect 14859 29884 14860 29924
rect 14900 29884 14901 29924
rect 14859 29875 14901 29884
rect 14764 29840 14804 29851
rect 14764 29765 14804 29800
rect 14763 29756 14805 29765
rect 14763 29716 14764 29756
rect 14804 29716 14805 29756
rect 14763 29707 14805 29716
rect 14860 29252 14900 29875
rect 14956 29345 14996 30640
rect 15051 30260 15093 30269
rect 15051 30220 15052 30260
rect 15092 30220 15093 30260
rect 15051 30211 15093 30220
rect 15052 29588 15092 30211
rect 15148 29840 15188 32143
rect 15244 31529 15284 32152
rect 15340 32192 15380 32201
rect 15243 31520 15285 31529
rect 15243 31480 15244 31520
rect 15284 31480 15285 31520
rect 15243 31471 15285 31480
rect 15340 31277 15380 32152
rect 15339 31268 15381 31277
rect 15339 31228 15340 31268
rect 15380 31228 15381 31268
rect 15339 31219 15381 31228
rect 15436 30353 15476 34336
rect 15532 34327 15572 34336
rect 15531 31352 15573 31361
rect 15531 31312 15532 31352
rect 15572 31312 15573 31352
rect 15531 31303 15573 31312
rect 15532 31218 15572 31303
rect 15531 30596 15573 30605
rect 15531 30556 15532 30596
rect 15572 30556 15573 30596
rect 15531 30547 15573 30556
rect 15435 30344 15477 30353
rect 15435 30304 15436 30344
rect 15476 30304 15477 30344
rect 15435 30295 15477 30304
rect 15340 29840 15380 29849
rect 15148 29800 15340 29840
rect 15244 29597 15284 29800
rect 15340 29791 15380 29800
rect 15339 29672 15381 29681
rect 15339 29632 15340 29672
rect 15380 29632 15381 29672
rect 15339 29623 15381 29632
rect 15243 29588 15285 29597
rect 15052 29548 15188 29588
rect 15051 29420 15093 29429
rect 15051 29380 15052 29420
rect 15092 29380 15093 29420
rect 15051 29371 15093 29380
rect 14955 29336 14997 29345
rect 14955 29296 14956 29336
rect 14996 29296 14997 29336
rect 14955 29287 14997 29296
rect 14764 29168 14804 29177
rect 14764 27245 14804 29128
rect 14763 27236 14805 27245
rect 14763 27196 14764 27236
rect 14804 27196 14805 27236
rect 14763 27187 14805 27196
rect 14860 26984 14900 29212
rect 15052 29168 15092 29371
rect 15148 29261 15188 29548
rect 15243 29548 15244 29588
rect 15284 29548 15285 29588
rect 15243 29539 15285 29548
rect 15147 29252 15189 29261
rect 15147 29212 15148 29252
rect 15188 29212 15189 29252
rect 15147 29203 15189 29212
rect 14956 29128 15092 29168
rect 14956 27161 14996 29128
rect 15051 29000 15093 29009
rect 15051 28960 15052 29000
rect 15092 28960 15093 29000
rect 15148 29000 15188 29203
rect 15340 29093 15380 29623
rect 15435 29504 15477 29513
rect 15435 29464 15436 29504
rect 15476 29464 15477 29504
rect 15435 29455 15477 29464
rect 15339 29084 15381 29093
rect 15339 29044 15340 29084
rect 15380 29044 15381 29084
rect 15339 29035 15381 29044
rect 15148 28960 15284 29000
rect 15051 28951 15093 28960
rect 14955 27152 14997 27161
rect 14955 27112 14956 27152
rect 14996 27112 14997 27152
rect 14955 27103 14997 27112
rect 14860 26944 14996 26984
rect 14764 26816 14804 26827
rect 14764 26741 14804 26776
rect 14859 26816 14901 26825
rect 14859 26776 14860 26816
rect 14900 26776 14901 26816
rect 14859 26767 14901 26776
rect 14763 26732 14805 26741
rect 14763 26692 14764 26732
rect 14804 26692 14805 26732
rect 14763 26683 14805 26692
rect 14860 26682 14900 26767
rect 14956 26489 14996 26944
rect 15052 26648 15092 28951
rect 15148 28874 15188 28883
rect 15148 26825 15188 28834
rect 15244 28337 15284 28960
rect 15243 28328 15285 28337
rect 15243 28288 15244 28328
rect 15284 28288 15285 28328
rect 15243 28279 15285 28288
rect 15244 28194 15284 28279
rect 15244 27656 15284 27667
rect 15244 27581 15284 27616
rect 15243 27572 15285 27581
rect 15243 27532 15244 27572
rect 15284 27532 15285 27572
rect 15243 27523 15285 27532
rect 15243 26900 15285 26909
rect 15243 26860 15244 26900
rect 15284 26860 15285 26900
rect 15243 26851 15285 26860
rect 15147 26816 15189 26825
rect 15147 26776 15148 26816
rect 15188 26776 15189 26816
rect 15147 26767 15189 26776
rect 15244 26766 15284 26851
rect 15052 26599 15092 26608
rect 14955 26480 14997 26489
rect 14955 26440 14956 26480
rect 14996 26440 14997 26480
rect 14955 26431 14997 26440
rect 15052 26144 15092 26153
rect 15092 26104 15188 26144
rect 15052 26095 15092 26104
rect 15148 25565 15188 26104
rect 15340 25976 15380 29035
rect 15436 28580 15476 29455
rect 15436 28531 15476 28540
rect 15435 27908 15477 27917
rect 15435 27868 15436 27908
rect 15476 27868 15477 27908
rect 15435 27859 15477 27868
rect 15436 27824 15476 27859
rect 15436 27773 15476 27784
rect 15532 27665 15572 30547
rect 15628 29336 15668 34999
rect 15724 33881 15764 36427
rect 15819 35972 15861 35981
rect 15819 35932 15820 35972
rect 15860 35932 15861 35972
rect 15819 35923 15861 35932
rect 15723 33872 15765 33881
rect 15723 33832 15724 33872
rect 15764 33832 15765 33872
rect 15723 33823 15765 33832
rect 15724 33713 15764 33823
rect 15723 33704 15765 33713
rect 15723 33664 15724 33704
rect 15764 33664 15765 33704
rect 15723 33655 15765 33664
rect 15724 33570 15764 33655
rect 15723 32360 15765 32369
rect 15723 32320 15724 32360
rect 15764 32320 15765 32360
rect 15723 32311 15765 32320
rect 15724 32192 15764 32311
rect 15724 29681 15764 32152
rect 15820 32192 15860 35923
rect 16012 35300 16052 38200
rect 16300 38156 16340 38527
rect 16396 38408 16436 38417
rect 16492 38408 16532 38695
rect 16436 38368 16532 38408
rect 16396 38359 16436 38368
rect 16395 38240 16437 38249
rect 16395 38200 16396 38240
rect 16436 38200 16437 38240
rect 16395 38191 16437 38200
rect 15916 35260 16052 35300
rect 16108 38116 16340 38156
rect 15916 34385 15956 35260
rect 15915 34376 15957 34385
rect 15915 34336 15916 34376
rect 15956 34336 15957 34376
rect 15915 34327 15957 34336
rect 16012 34381 16052 34390
rect 15916 33872 15956 33881
rect 16012 33872 16052 34341
rect 15956 33832 16052 33872
rect 15916 33823 15956 33832
rect 16108 32369 16148 38116
rect 16299 37736 16341 37745
rect 16299 37696 16300 37736
rect 16340 37696 16341 37736
rect 16299 37687 16341 37696
rect 16300 36728 16340 37687
rect 16300 36679 16340 36688
rect 16396 37400 16436 38191
rect 16491 38156 16533 38165
rect 16491 38116 16492 38156
rect 16532 38116 16533 38156
rect 16491 38107 16533 38116
rect 16396 36569 16436 37360
rect 16395 36560 16437 36569
rect 16395 36520 16396 36560
rect 16436 36520 16437 36560
rect 16395 36511 16437 36520
rect 16492 36140 16532 38107
rect 16588 37241 16628 42064
rect 16683 39752 16725 39761
rect 16683 39712 16684 39752
rect 16724 39712 16725 39752
rect 16683 39703 16725 39712
rect 16587 37232 16629 37241
rect 16587 37192 16588 37232
rect 16628 37192 16629 37232
rect 16587 37183 16629 37192
rect 16587 36812 16629 36821
rect 16587 36772 16588 36812
rect 16628 36772 16629 36812
rect 16587 36763 16629 36772
rect 16396 36100 16532 36140
rect 16396 35468 16436 36100
rect 16588 35888 16628 36763
rect 16588 35729 16628 35848
rect 16587 35720 16629 35729
rect 16587 35680 16588 35720
rect 16628 35680 16629 35720
rect 16587 35671 16629 35680
rect 16300 35428 16436 35468
rect 16203 35216 16245 35225
rect 16203 35176 16204 35216
rect 16244 35176 16245 35216
rect 16203 35167 16245 35176
rect 16204 35082 16244 35167
rect 16300 35132 16340 35428
rect 16684 35393 16724 39703
rect 16972 37820 17012 44332
rect 17164 44288 17204 44407
rect 17164 44239 17204 44248
rect 17259 44288 17301 44297
rect 17259 44248 17260 44288
rect 17300 44248 17301 44288
rect 17356 44288 17396 45844
rect 17452 45800 17492 46423
rect 17452 45557 17492 45760
rect 17451 45548 17493 45557
rect 17451 45508 17452 45548
rect 17492 45508 17493 45548
rect 17451 45499 17493 45508
rect 17452 44288 17492 44297
rect 17356 44248 17452 44288
rect 17259 44239 17301 44248
rect 17452 44239 17492 44248
rect 17260 44154 17300 44239
rect 17163 43868 17205 43877
rect 17163 43828 17164 43868
rect 17204 43828 17205 43868
rect 17163 43819 17205 43828
rect 17164 43448 17204 43819
rect 17164 43399 17204 43408
rect 17548 42785 17588 48607
rect 17739 47984 17781 47993
rect 17739 47944 17740 47984
rect 17780 47944 17781 47984
rect 17739 47935 17781 47944
rect 17643 47060 17685 47069
rect 17643 47020 17644 47060
rect 17684 47020 17685 47060
rect 17643 47011 17685 47020
rect 17644 44381 17684 47011
rect 17740 46397 17780 47935
rect 17739 46388 17781 46397
rect 17739 46348 17740 46388
rect 17780 46348 17781 46388
rect 17739 46339 17781 46348
rect 17739 46136 17781 46145
rect 17739 46096 17740 46136
rect 17780 46096 17781 46136
rect 17739 46087 17781 46096
rect 17740 45800 17780 46087
rect 17740 45751 17780 45760
rect 17739 45548 17781 45557
rect 17739 45508 17740 45548
rect 17780 45508 17781 45548
rect 17739 45499 17781 45508
rect 17740 45414 17780 45499
rect 17643 44372 17685 44381
rect 17643 44332 17644 44372
rect 17684 44332 17685 44372
rect 17643 44323 17685 44332
rect 17643 44204 17685 44213
rect 17643 44164 17644 44204
rect 17684 44164 17685 44204
rect 17643 44155 17685 44164
rect 17547 42776 17589 42785
rect 17547 42736 17548 42776
rect 17588 42736 17589 42776
rect 17547 42727 17589 42736
rect 17260 42608 17300 42617
rect 17260 41945 17300 42568
rect 17259 41936 17301 41945
rect 17259 41896 17260 41936
rect 17300 41896 17301 41936
rect 17259 41887 17301 41896
rect 17260 41096 17300 41887
rect 17163 40424 17205 40433
rect 17163 40384 17164 40424
rect 17204 40384 17205 40424
rect 17163 40375 17205 40384
rect 17164 39080 17204 40375
rect 17260 40256 17300 41056
rect 17260 39920 17300 40216
rect 17260 39871 17300 39880
rect 17451 39752 17493 39761
rect 17451 39712 17452 39752
rect 17492 39712 17493 39752
rect 17451 39703 17493 39712
rect 17356 39584 17396 39593
rect 17260 39080 17300 39089
rect 17164 39040 17260 39080
rect 17260 39031 17300 39040
rect 17259 38744 17301 38753
rect 17356 38744 17396 39544
rect 17452 38912 17492 39703
rect 17452 38863 17492 38872
rect 17259 38704 17260 38744
rect 17300 38704 17396 38744
rect 17259 38695 17301 38704
rect 16780 37780 17012 37820
rect 17260 38408 17300 38695
rect 17644 38501 17684 44155
rect 17836 44129 17876 48784
rect 18028 48819 18068 49279
rect 18028 48770 18068 48779
rect 18124 48656 18164 49531
rect 18028 48616 18164 48656
rect 18220 49496 18260 49505
rect 18316 49496 18356 51715
rect 18411 51680 18453 51689
rect 18411 51640 18412 51680
rect 18452 51640 18453 51680
rect 18411 51631 18453 51640
rect 18412 50924 18452 51631
rect 18412 50875 18452 50884
rect 18411 50336 18453 50345
rect 18411 50296 18412 50336
rect 18452 50296 18453 50336
rect 18411 50287 18453 50296
rect 18412 49748 18452 50287
rect 18412 49699 18452 49708
rect 18260 49456 18356 49496
rect 18028 47321 18068 48616
rect 18220 47993 18260 49456
rect 18411 49328 18453 49337
rect 18411 49288 18412 49328
rect 18452 49288 18453 49328
rect 18411 49279 18453 49288
rect 18412 49194 18452 49279
rect 18508 49001 18548 52303
rect 18604 51773 18644 52480
rect 18700 51941 18740 52807
rect 18795 52520 18837 52529
rect 18795 52480 18796 52520
rect 18836 52480 18837 52520
rect 18795 52471 18837 52480
rect 18699 51932 18741 51941
rect 18699 51892 18700 51932
rect 18740 51892 18741 51932
rect 18699 51883 18741 51892
rect 18700 51848 18740 51883
rect 18700 51797 18740 51808
rect 18603 51764 18645 51773
rect 18603 51724 18604 51764
rect 18644 51724 18645 51764
rect 18603 51715 18645 51724
rect 18603 51596 18645 51605
rect 18796 51596 18836 52471
rect 18603 51556 18604 51596
rect 18644 51556 18645 51596
rect 18603 51547 18645 51556
rect 18700 51556 18836 51596
rect 18604 51022 18644 51547
rect 18604 50973 18644 50982
rect 18603 49496 18645 49505
rect 18603 49456 18604 49496
rect 18644 49456 18645 49496
rect 18603 49447 18645 49456
rect 18604 49362 18644 49447
rect 18507 48992 18549 49001
rect 18507 48952 18508 48992
rect 18548 48952 18549 48992
rect 18507 48943 18549 48952
rect 18508 48824 18548 48833
rect 18508 48497 18548 48784
rect 18700 48665 18740 51556
rect 18808 51428 19176 51437
rect 18848 51388 18890 51428
rect 18930 51388 18972 51428
rect 19012 51388 19054 51428
rect 19094 51388 19136 51428
rect 18808 51379 19176 51388
rect 18891 51260 18933 51269
rect 18891 51220 18892 51260
rect 18932 51220 18933 51260
rect 18891 51211 18933 51220
rect 18796 50336 18836 50345
rect 18892 50336 18932 51211
rect 19372 51017 19412 53824
rect 19468 53537 19508 53992
rect 19467 53528 19509 53537
rect 19467 53488 19468 53528
rect 19508 53488 19509 53528
rect 19467 53479 19509 53488
rect 19659 53360 19701 53369
rect 19659 53320 19660 53360
rect 19700 53320 19701 53360
rect 19659 53311 19701 53320
rect 19660 53226 19700 53311
rect 19467 53192 19509 53201
rect 19467 53152 19468 53192
rect 19508 53152 19509 53192
rect 19467 53143 19509 53152
rect 19468 53058 19508 53143
rect 19756 53117 19796 56092
rect 19852 56083 19892 56092
rect 19851 55796 19893 55805
rect 19851 55756 19852 55796
rect 19892 55756 19893 55796
rect 19851 55747 19893 55756
rect 19852 55662 19892 55747
rect 20044 55460 20084 56344
rect 19948 55420 20084 55460
rect 20140 56384 20180 56393
rect 19851 55376 19893 55385
rect 19851 55336 19852 55376
rect 19892 55336 19893 55376
rect 19851 55327 19893 55336
rect 19852 54368 19892 55327
rect 19948 55040 19988 55420
rect 20140 55385 20180 56344
rect 20139 55376 20181 55385
rect 20139 55336 20140 55376
rect 20180 55336 20181 55376
rect 20139 55327 20181 55336
rect 20048 55208 20416 55217
rect 20088 55168 20130 55208
rect 20170 55168 20212 55208
rect 20252 55168 20294 55208
rect 20334 55168 20376 55208
rect 20048 55159 20416 55168
rect 19948 55000 20084 55040
rect 19947 54872 19989 54881
rect 19947 54832 19948 54872
rect 19988 54832 19989 54872
rect 19947 54823 19989 54832
rect 19948 54738 19988 54823
rect 19852 54328 19988 54368
rect 19851 54200 19893 54209
rect 19851 54160 19852 54200
rect 19892 54160 19893 54200
rect 19851 54151 19893 54160
rect 19852 54032 19892 54151
rect 19948 54041 19988 54328
rect 19852 53621 19892 53992
rect 19947 54032 19989 54041
rect 19947 53992 19948 54032
rect 19988 53992 19989 54032
rect 19947 53983 19989 53992
rect 20044 53864 20084 55000
rect 19948 53824 20084 53864
rect 19851 53612 19893 53621
rect 19851 53572 19852 53612
rect 19892 53572 19893 53612
rect 19851 53563 19893 53572
rect 19948 53528 19988 53824
rect 20048 53696 20416 53705
rect 20088 53656 20130 53696
rect 20170 53656 20212 53696
rect 20252 53656 20294 53696
rect 20334 53656 20376 53696
rect 20048 53647 20416 53656
rect 20140 53528 20180 53537
rect 19948 53488 20140 53528
rect 20140 53479 20180 53488
rect 19852 53360 19892 53369
rect 19660 53108 19700 53117
rect 19563 53024 19605 53033
rect 19660 53024 19700 53068
rect 19755 53108 19797 53117
rect 19755 53068 19756 53108
rect 19796 53068 19797 53108
rect 19755 53059 19797 53068
rect 19563 52984 19564 53024
rect 19604 52984 19700 53024
rect 19563 52975 19605 52984
rect 19852 52940 19892 53320
rect 19948 53360 19988 53369
rect 19948 52949 19988 53320
rect 20235 53360 20277 53369
rect 20235 53320 20236 53360
rect 20276 53320 20277 53360
rect 20235 53311 20277 53320
rect 20236 53226 20276 53311
rect 20043 53108 20085 53117
rect 20043 53068 20044 53108
rect 20084 53068 20085 53108
rect 20043 53059 20085 53068
rect 19660 52900 19892 52940
rect 19947 52940 19989 52949
rect 19947 52900 19948 52940
rect 19988 52900 19989 52940
rect 19660 52781 19700 52900
rect 19947 52891 19989 52900
rect 19659 52772 19701 52781
rect 19659 52732 19660 52772
rect 19700 52732 19701 52772
rect 19659 52723 19701 52732
rect 19851 52772 19893 52781
rect 19851 52732 19852 52772
rect 19892 52732 19893 52772
rect 19851 52723 19893 52732
rect 19659 52520 19701 52529
rect 19659 52480 19660 52520
rect 19700 52480 19701 52520
rect 19659 52471 19701 52480
rect 19852 52520 19892 52723
rect 19947 52688 19989 52697
rect 19947 52648 19948 52688
rect 19988 52648 19989 52688
rect 19947 52639 19989 52648
rect 19852 52471 19892 52480
rect 19948 52520 19988 52639
rect 19948 52471 19988 52480
rect 20044 52520 20084 53059
rect 20140 52613 20180 52660
rect 20139 52604 20181 52613
rect 20139 52555 20140 52604
rect 20180 52555 20181 52604
rect 20140 52516 20180 52525
rect 20044 52471 20084 52480
rect 19660 52386 19700 52471
rect 20048 52184 20416 52193
rect 20088 52144 20130 52184
rect 20170 52144 20212 52184
rect 20252 52144 20294 52184
rect 20334 52144 20376 52184
rect 20048 52135 20416 52144
rect 19948 51848 19988 51857
rect 19948 51269 19988 51808
rect 20139 51596 20181 51605
rect 20139 51556 20140 51596
rect 20180 51556 20181 51596
rect 20139 51547 20181 51556
rect 20140 51462 20180 51547
rect 19947 51260 19989 51269
rect 19947 51220 19948 51260
rect 19988 51220 19989 51260
rect 19947 51211 19989 51220
rect 19563 51092 19605 51101
rect 19563 51052 19564 51092
rect 19604 51052 19605 51092
rect 19563 51043 19605 51052
rect 19083 51008 19125 51017
rect 19083 50968 19084 51008
rect 19124 50968 19125 51008
rect 19083 50959 19125 50968
rect 19371 51008 19413 51017
rect 19371 50968 19372 51008
rect 19412 50968 19413 51008
rect 19371 50959 19413 50968
rect 19084 50874 19124 50959
rect 19564 50958 19604 51043
rect 19660 51008 19700 51017
rect 20044 51008 20084 51017
rect 19660 50588 19700 50968
rect 19948 50968 20044 51008
rect 19948 50681 19988 50968
rect 20044 50959 20084 50968
rect 20140 50988 20180 50997
rect 20140 50849 20180 50948
rect 20139 50840 20181 50849
rect 20139 50800 20140 50840
rect 20180 50800 20181 50840
rect 20139 50791 20181 50800
rect 19947 50672 19989 50681
rect 19947 50632 19948 50672
rect 19988 50632 19989 50672
rect 19947 50623 19989 50632
rect 20048 50672 20416 50681
rect 20088 50632 20130 50672
rect 20170 50632 20212 50672
rect 20252 50632 20294 50672
rect 20334 50632 20376 50672
rect 20048 50623 20416 50632
rect 19084 50548 19700 50588
rect 18987 50420 19029 50429
rect 18987 50380 18988 50420
rect 19028 50380 19029 50420
rect 18987 50371 19029 50380
rect 18836 50296 18932 50336
rect 18796 50177 18836 50296
rect 18988 50286 19028 50371
rect 18795 50168 18837 50177
rect 18795 50128 18796 50168
rect 18836 50128 18837 50168
rect 18795 50119 18837 50128
rect 19084 50084 19124 50548
rect 19276 50420 19316 50429
rect 19179 50336 19221 50345
rect 19179 50296 19180 50336
rect 19220 50296 19221 50336
rect 19179 50287 19221 50296
rect 19180 50202 19220 50287
rect 19276 50168 19316 50380
rect 19372 50345 19412 50430
rect 19468 50380 19796 50420
rect 19371 50336 19413 50345
rect 19371 50296 19372 50336
rect 19412 50296 19413 50336
rect 19371 50287 19413 50296
rect 19468 50336 19508 50380
rect 19756 50336 19796 50380
rect 19371 50168 19413 50177
rect 19276 50128 19372 50168
rect 19412 50128 19413 50168
rect 19371 50119 19413 50128
rect 19084 50044 19316 50084
rect 18808 49916 19176 49925
rect 18848 49876 18890 49916
rect 18930 49876 18972 49916
rect 19012 49876 19054 49916
rect 19094 49876 19136 49916
rect 18808 49867 19176 49876
rect 18891 48908 18933 48917
rect 19083 48908 19125 48917
rect 18891 48868 18892 48908
rect 18932 48868 19028 48908
rect 18891 48859 18933 48868
rect 18988 48824 19028 48868
rect 19083 48868 19084 48908
rect 19124 48868 19125 48908
rect 19083 48859 19125 48868
rect 18988 48775 19028 48784
rect 19084 48824 19124 48859
rect 19084 48773 19124 48784
rect 18699 48656 18741 48665
rect 18699 48616 18700 48656
rect 18740 48616 18741 48656
rect 18699 48607 18741 48616
rect 18507 48488 18549 48497
rect 18507 48448 18508 48488
rect 18548 48448 18549 48488
rect 18507 48439 18549 48448
rect 18603 48404 18645 48413
rect 18603 48364 18604 48404
rect 18644 48364 18645 48404
rect 18603 48355 18645 48364
rect 18808 48404 19176 48413
rect 18848 48364 18890 48404
rect 18930 48364 18972 48404
rect 19012 48364 19054 48404
rect 19094 48364 19136 48404
rect 18808 48355 19176 48364
rect 18411 48236 18453 48245
rect 18411 48196 18412 48236
rect 18452 48196 18453 48236
rect 18411 48187 18453 48196
rect 18412 48102 18452 48187
rect 18219 47984 18261 47993
rect 18219 47944 18220 47984
rect 18260 47944 18261 47984
rect 18219 47935 18261 47944
rect 18604 47984 18644 48355
rect 19276 47993 19316 50044
rect 19371 49916 19413 49925
rect 19371 49876 19372 49916
rect 19412 49876 19413 49916
rect 19371 49867 19413 49876
rect 18604 47935 18644 47944
rect 19275 47984 19317 47993
rect 19275 47944 19276 47984
rect 19316 47944 19317 47984
rect 19275 47935 19317 47944
rect 18220 47850 18260 47935
rect 18123 47732 18165 47741
rect 18123 47692 18124 47732
rect 18164 47692 18165 47732
rect 18123 47683 18165 47692
rect 18027 47312 18069 47321
rect 18027 47272 18028 47312
rect 18068 47272 18069 47312
rect 18027 47263 18069 47272
rect 18028 47178 18068 47263
rect 17931 46304 17973 46313
rect 17931 46264 17932 46304
rect 17972 46264 17973 46304
rect 17931 46255 17973 46264
rect 17932 45800 17972 46255
rect 18124 46145 18164 47683
rect 18604 47312 18644 47321
rect 18604 47069 18644 47272
rect 19275 47144 19317 47153
rect 19275 47104 19276 47144
rect 19316 47104 19317 47144
rect 19275 47095 19317 47104
rect 18220 47060 18260 47069
rect 18603 47060 18645 47069
rect 18260 47020 18548 47060
rect 18220 47011 18260 47020
rect 18508 46472 18548 47020
rect 18603 47020 18604 47060
rect 18644 47020 18645 47060
rect 18603 47011 18645 47020
rect 18808 46892 19176 46901
rect 18848 46852 18890 46892
rect 18930 46852 18972 46892
rect 19012 46852 19054 46892
rect 19094 46852 19136 46892
rect 18808 46843 19176 46852
rect 19276 46724 19316 47095
rect 18988 46684 19316 46724
rect 18604 46481 18644 46566
rect 18508 46423 18548 46432
rect 18603 46472 18645 46481
rect 18603 46432 18604 46472
rect 18644 46432 18645 46472
rect 18603 46423 18645 46432
rect 18988 46472 19028 46684
rect 19372 46640 19412 49867
rect 19468 49328 19508 50296
rect 19660 50291 19700 50300
rect 19948 50336 19988 50345
rect 19756 50287 19796 50296
rect 19852 50294 19892 50303
rect 19660 50093 19700 50251
rect 19755 50168 19797 50177
rect 19852 50168 19892 50254
rect 19755 50128 19756 50168
rect 19796 50128 19892 50168
rect 19755 50119 19797 50128
rect 19659 50084 19701 50093
rect 19659 50044 19660 50084
rect 19700 50044 19701 50084
rect 19659 50035 19701 50044
rect 19660 49925 19700 50035
rect 19659 49916 19701 49925
rect 19659 49876 19660 49916
rect 19700 49876 19701 49916
rect 19659 49867 19701 49876
rect 19851 49496 19893 49505
rect 19851 49456 19852 49496
rect 19892 49456 19893 49496
rect 19851 49447 19893 49456
rect 19852 49362 19892 49447
rect 19468 49288 19604 49328
rect 19468 48824 19508 48833
rect 19468 48749 19508 48784
rect 19564 48824 19604 49288
rect 19851 48992 19893 49001
rect 19851 48952 19852 48992
rect 19892 48952 19893 48992
rect 19948 48992 19988 50296
rect 20139 50336 20181 50345
rect 20139 50296 20140 50336
rect 20180 50296 20181 50336
rect 20139 50287 20181 50296
rect 20236 50336 20276 50347
rect 20140 50202 20180 50287
rect 20236 50261 20276 50296
rect 20620 50261 20660 57847
rect 20716 53369 20756 58099
rect 21004 57737 21044 60535
rect 21195 58232 21237 58241
rect 21195 58192 21196 58232
rect 21236 58192 21237 58232
rect 21195 58183 21237 58192
rect 21003 57728 21045 57737
rect 21003 57688 21004 57728
rect 21044 57688 21045 57728
rect 21003 57679 21045 57688
rect 20811 56216 20853 56225
rect 20811 56176 20812 56216
rect 20852 56176 20853 56216
rect 20811 56167 20853 56176
rect 20812 55889 20852 56167
rect 20811 55880 20853 55889
rect 20811 55840 20812 55880
rect 20852 55840 20853 55880
rect 20811 55831 20853 55840
rect 20715 53360 20757 53369
rect 20715 53320 20716 53360
rect 20756 53320 20757 53360
rect 20715 53311 20757 53320
rect 20812 52613 20852 55831
rect 20811 52604 20853 52613
rect 20811 52564 20812 52604
rect 20852 52564 20853 52604
rect 20811 52555 20853 52564
rect 20812 51101 20852 52555
rect 20907 51512 20949 51521
rect 20907 51472 20908 51512
rect 20948 51472 20949 51512
rect 20907 51463 20949 51472
rect 20811 51092 20853 51101
rect 20811 51052 20812 51092
rect 20852 51052 20853 51092
rect 20811 51043 20853 51052
rect 20235 50252 20277 50261
rect 20235 50212 20236 50252
rect 20276 50212 20277 50252
rect 20235 50203 20277 50212
rect 20619 50252 20661 50261
rect 20619 50212 20620 50252
rect 20660 50212 20661 50252
rect 20619 50203 20661 50212
rect 20523 50000 20565 50009
rect 20523 49960 20524 50000
rect 20564 49960 20565 50000
rect 20523 49951 20565 49960
rect 20044 49337 20084 49422
rect 20043 49328 20085 49337
rect 20043 49288 20044 49328
rect 20084 49288 20085 49328
rect 20043 49279 20085 49288
rect 20524 49169 20564 49951
rect 20619 49832 20661 49841
rect 20619 49792 20620 49832
rect 20660 49792 20661 49832
rect 20619 49783 20661 49792
rect 20048 49160 20416 49169
rect 20088 49120 20130 49160
rect 20170 49120 20212 49160
rect 20252 49120 20294 49160
rect 20334 49120 20376 49160
rect 20048 49111 20416 49120
rect 20523 49160 20565 49169
rect 20523 49120 20524 49160
rect 20564 49120 20565 49160
rect 20523 49111 20565 49120
rect 19948 48952 20180 48992
rect 19851 48943 19893 48952
rect 19467 48740 19509 48749
rect 19467 48700 19468 48740
rect 19508 48700 19509 48740
rect 19467 48691 19509 48700
rect 19468 48329 19508 48691
rect 19467 48320 19509 48329
rect 19467 48280 19468 48320
rect 19508 48280 19509 48320
rect 19467 48271 19509 48280
rect 19564 48245 19604 48784
rect 19852 48824 19892 48943
rect 19852 48775 19892 48784
rect 20044 48824 20084 48833
rect 20044 48665 20084 48784
rect 20140 48824 20180 48952
rect 20140 48775 20180 48784
rect 20620 48665 20660 49783
rect 20043 48656 20085 48665
rect 20043 48616 20044 48656
rect 20084 48616 20085 48656
rect 20043 48607 20085 48616
rect 20619 48656 20661 48665
rect 20619 48616 20620 48656
rect 20660 48616 20661 48656
rect 20619 48607 20661 48616
rect 19851 48572 19893 48581
rect 19851 48532 19852 48572
rect 19892 48532 19893 48572
rect 19851 48523 19893 48532
rect 19852 48438 19892 48523
rect 19563 48236 19605 48245
rect 19563 48196 19564 48236
rect 19604 48196 19605 48236
rect 19563 48187 19605 48196
rect 20044 48236 20084 48607
rect 20044 48187 20084 48196
rect 19563 48068 19605 48077
rect 19563 48028 19564 48068
rect 19604 48028 19605 48068
rect 19563 48019 19605 48028
rect 19084 46600 19412 46640
rect 19084 46556 19124 46600
rect 19084 46507 19124 46516
rect 18603 46304 18645 46313
rect 18603 46264 18604 46304
rect 18644 46264 18645 46304
rect 18603 46255 18645 46264
rect 18123 46136 18165 46145
rect 18123 46096 18124 46136
rect 18164 46096 18165 46136
rect 18123 46087 18165 46096
rect 18411 46136 18453 46145
rect 18411 46096 18412 46136
rect 18452 46096 18453 46136
rect 18411 46087 18453 46096
rect 17932 45751 17972 45760
rect 18028 45800 18068 45809
rect 17931 45632 17973 45641
rect 17931 45592 17932 45632
rect 17972 45592 17973 45632
rect 17931 45583 17973 45592
rect 17932 45498 17972 45583
rect 18028 45557 18068 45760
rect 18219 45800 18261 45809
rect 18219 45760 18220 45800
rect 18260 45760 18261 45800
rect 18219 45751 18261 45760
rect 18412 45800 18452 46087
rect 18412 45751 18452 45760
rect 18220 45666 18260 45751
rect 18027 45548 18069 45557
rect 18027 45508 18028 45548
rect 18068 45508 18069 45548
rect 18027 45499 18069 45508
rect 18411 45464 18453 45473
rect 18411 45424 18412 45464
rect 18452 45424 18453 45464
rect 18411 45415 18453 45424
rect 17931 45380 17973 45389
rect 17931 45340 17932 45380
rect 17972 45340 17973 45380
rect 17931 45331 17973 45340
rect 17932 44960 17972 45331
rect 18412 45128 18452 45415
rect 18412 45088 18548 45128
rect 17835 44120 17877 44129
rect 17835 44080 17836 44120
rect 17876 44080 17877 44120
rect 17835 44071 17877 44080
rect 17932 43541 17972 44920
rect 18412 44960 18452 44969
rect 18124 44792 18164 44801
rect 18124 44288 18164 44752
rect 18220 44288 18260 44297
rect 18124 44248 18220 44288
rect 18220 44239 18260 44248
rect 18316 44288 18356 44297
rect 18316 44129 18356 44248
rect 18315 44120 18357 44129
rect 18315 44080 18316 44120
rect 18356 44080 18357 44120
rect 18315 44071 18357 44080
rect 18315 43952 18357 43961
rect 18315 43912 18316 43952
rect 18356 43912 18357 43952
rect 18315 43903 18357 43912
rect 17931 43532 17973 43541
rect 17931 43492 17932 43532
rect 17972 43492 17973 43532
rect 17931 43483 17973 43492
rect 18316 43205 18356 43903
rect 18412 43700 18452 44920
rect 18508 44960 18548 45088
rect 18508 43961 18548 44920
rect 18507 43952 18549 43961
rect 18507 43912 18508 43952
rect 18548 43912 18549 43952
rect 18507 43903 18549 43912
rect 18604 43868 18644 46255
rect 18988 45800 19028 46432
rect 18700 45760 19028 45800
rect 19564 46472 19604 48019
rect 19852 47984 19892 47995
rect 19852 47909 19892 47944
rect 19947 47984 19989 47993
rect 19947 47944 19948 47984
rect 19988 47944 19989 47984
rect 19947 47935 19989 47944
rect 19851 47900 19893 47909
rect 19851 47860 19852 47900
rect 19892 47860 19893 47900
rect 19851 47851 19893 47860
rect 19852 47312 19892 47321
rect 19852 46985 19892 47272
rect 19851 46976 19893 46985
rect 19851 46936 19852 46976
rect 19892 46936 19893 46976
rect 19851 46927 19893 46936
rect 19948 46724 19988 47935
rect 20048 47648 20416 47657
rect 20088 47608 20130 47648
rect 20170 47608 20212 47648
rect 20252 47608 20294 47648
rect 20334 47608 20376 47648
rect 20048 47599 20416 47608
rect 20044 47060 20084 47069
rect 20084 47020 20180 47060
rect 20044 47011 20084 47020
rect 19852 46684 19988 46724
rect 19852 46640 19892 46684
rect 18700 45212 18740 45760
rect 18808 45380 19176 45389
rect 18848 45340 18890 45380
rect 18930 45340 18972 45380
rect 19012 45340 19054 45380
rect 19094 45340 19136 45380
rect 18808 45331 19176 45340
rect 18987 45212 19029 45221
rect 18700 45172 18836 45212
rect 18699 44456 18741 44465
rect 18699 44416 18700 44456
rect 18740 44416 18741 44456
rect 18699 44407 18741 44416
rect 18700 44288 18740 44407
rect 18700 44239 18740 44248
rect 18796 44288 18836 45172
rect 18987 45172 18988 45212
rect 19028 45172 19029 45212
rect 18987 45163 19029 45172
rect 18891 45044 18933 45053
rect 18891 45004 18892 45044
rect 18932 45004 18933 45044
rect 18891 44995 18933 45004
rect 18988 45044 19028 45163
rect 18988 44995 19028 45004
rect 18892 44910 18932 44995
rect 19468 44960 19508 44969
rect 19468 44717 19508 44920
rect 19467 44708 19509 44717
rect 19467 44668 19468 44708
rect 19508 44668 19509 44708
rect 19467 44659 19509 44668
rect 18796 44239 18836 44248
rect 19276 44288 19316 44297
rect 19564 44288 19604 46432
rect 19756 46600 19892 46640
rect 19660 45800 19700 45809
rect 19660 45557 19700 45760
rect 19659 45548 19701 45557
rect 19659 45508 19660 45548
rect 19700 45508 19701 45548
rect 19659 45499 19701 45508
rect 19756 45053 19796 46600
rect 20044 46481 20084 46567
rect 20140 46481 20180 47020
rect 20908 46649 20948 51463
rect 21196 51353 21236 58183
rect 21387 56384 21429 56393
rect 21387 56344 21388 56384
rect 21428 56344 21429 56384
rect 21387 56335 21429 56344
rect 21388 55889 21428 56335
rect 21387 55880 21429 55889
rect 21387 55840 21388 55880
rect 21428 55840 21429 55880
rect 21387 55831 21429 55840
rect 21195 51344 21237 51353
rect 21195 51304 21196 51344
rect 21236 51304 21237 51344
rect 21195 51295 21237 51304
rect 20907 46640 20949 46649
rect 20907 46600 20908 46640
rect 20948 46600 20949 46640
rect 20907 46591 20949 46600
rect 20043 46477 20085 46481
rect 20043 46432 20044 46477
rect 20084 46432 20085 46477
rect 20043 46423 20085 46432
rect 20139 46431 20180 46481
rect 20140 46304 20180 46431
rect 20235 46388 20277 46397
rect 20235 46348 20236 46388
rect 20276 46348 20277 46388
rect 20235 46339 20277 46348
rect 19948 46264 20180 46304
rect 19852 45548 19892 45557
rect 19755 45044 19797 45053
rect 19755 45004 19756 45044
rect 19796 45004 19797 45044
rect 19755 44995 19797 45004
rect 19852 44288 19892 45508
rect 19948 44974 19988 46264
rect 20236 46254 20276 46339
rect 20048 46136 20416 46145
rect 20088 46096 20130 46136
rect 20170 46096 20212 46136
rect 20252 46096 20294 46136
rect 20334 46096 20376 46136
rect 20048 46087 20416 46096
rect 19948 44925 19988 44934
rect 20140 44792 20180 44801
rect 20180 44752 20564 44792
rect 20140 44743 20180 44752
rect 20048 44624 20416 44633
rect 20088 44584 20130 44624
rect 20170 44584 20212 44624
rect 20252 44584 20294 44624
rect 20334 44584 20376 44624
rect 20048 44575 20416 44584
rect 19316 44248 19604 44288
rect 19804 44278 19892 44288
rect 19276 44239 19316 44248
rect 19844 44248 19892 44278
rect 19948 44372 19988 44381
rect 19804 44229 19844 44238
rect 19948 44213 19988 44332
rect 19947 44204 19989 44213
rect 19947 44164 19948 44204
rect 19988 44164 19989 44204
rect 19947 44155 19989 44164
rect 18808 43868 19176 43877
rect 18604 43828 18740 43868
rect 18604 43700 18644 43709
rect 18412 43660 18604 43700
rect 18604 43651 18644 43660
rect 18700 43532 18740 43828
rect 18848 43828 18890 43868
rect 18930 43828 18972 43868
rect 19012 43828 19054 43868
rect 19094 43828 19136 43868
rect 18808 43819 19176 43828
rect 18412 43492 18740 43532
rect 18412 43448 18452 43492
rect 18412 43399 18452 43408
rect 18988 43280 19028 43289
rect 18315 43196 18357 43205
rect 18315 43156 18316 43196
rect 18356 43156 18357 43196
rect 18315 43147 18357 43156
rect 18988 42608 19028 43240
rect 20048 43112 20416 43121
rect 20088 43072 20130 43112
rect 20170 43072 20212 43112
rect 20252 43072 20294 43112
rect 20334 43072 20376 43112
rect 20048 43063 20416 43072
rect 20235 42776 20277 42785
rect 20235 42736 20236 42776
rect 20276 42736 20277 42776
rect 20235 42727 20277 42736
rect 19756 42617 19796 42702
rect 20044 42692 20084 42703
rect 20044 42617 20084 42652
rect 18988 42524 19028 42568
rect 19755 42608 19797 42617
rect 19755 42568 19756 42608
rect 19796 42568 19797 42608
rect 19755 42559 19797 42568
rect 20043 42608 20085 42617
rect 20043 42568 20044 42608
rect 20084 42568 20085 42608
rect 20043 42559 20085 42568
rect 20236 42608 20276 42727
rect 20236 42559 20276 42568
rect 18700 42484 19028 42524
rect 19563 42524 19605 42533
rect 19563 42484 19564 42524
rect 19604 42484 19700 42524
rect 18123 42440 18165 42449
rect 18123 42400 18124 42440
rect 18164 42400 18165 42440
rect 18123 42391 18165 42400
rect 18124 42188 18164 42391
rect 18124 42139 18164 42148
rect 17931 42104 17973 42113
rect 17931 42064 17932 42104
rect 17972 42064 17973 42104
rect 17931 42055 17973 42064
rect 17932 42020 17972 42055
rect 17932 41969 17972 41980
rect 18123 42020 18165 42029
rect 18123 41980 18124 42020
rect 18164 41980 18165 42020
rect 18123 41971 18165 41980
rect 17739 41936 17781 41945
rect 17739 41896 17740 41936
rect 17780 41896 17781 41936
rect 17739 41887 17781 41896
rect 17740 41802 17780 41887
rect 17835 40676 17877 40685
rect 17835 40636 17836 40676
rect 17876 40636 17877 40676
rect 17835 40627 17877 40636
rect 17836 40508 17876 40627
rect 17836 40459 17876 40468
rect 18028 40592 18068 40601
rect 18028 40433 18068 40552
rect 18027 40424 18069 40433
rect 18027 40384 18028 40424
rect 18068 40384 18069 40424
rect 18027 40375 18069 40384
rect 17643 38492 17685 38501
rect 17643 38452 17644 38492
rect 17684 38452 17685 38492
rect 17643 38443 17685 38452
rect 16780 36812 16820 37780
rect 16924 37409 16964 37418
rect 16964 37369 17012 37400
rect 16924 37360 17012 37369
rect 16972 36989 17012 37360
rect 17067 37316 17109 37325
rect 17067 37276 17068 37316
rect 17108 37276 17109 37316
rect 17067 37267 17109 37276
rect 17068 37182 17108 37267
rect 17260 37232 17300 38368
rect 16971 36980 17013 36989
rect 16971 36940 16972 36980
rect 17012 36940 17013 36980
rect 16971 36931 17013 36940
rect 16971 36812 17013 36821
rect 16780 36772 16916 36812
rect 16780 36714 16820 36723
rect 16683 35384 16725 35393
rect 16683 35344 16684 35384
rect 16724 35344 16725 35384
rect 16683 35335 16725 35344
rect 16396 35300 16436 35309
rect 16396 35216 16436 35260
rect 16780 35216 16820 36674
rect 16396 35176 16820 35216
rect 16300 35092 16436 35132
rect 16204 34208 16244 34217
rect 16107 32360 16149 32369
rect 16107 32320 16108 32360
rect 16148 32320 16149 32360
rect 16107 32311 16149 32320
rect 15820 30017 15860 32152
rect 16204 31529 16244 34168
rect 16299 32192 16341 32201
rect 16299 32152 16300 32192
rect 16340 32152 16341 32192
rect 16299 32143 16341 32152
rect 16300 32058 16340 32143
rect 16396 31604 16436 35092
rect 16876 35048 16916 36772
rect 16971 36772 16972 36812
rect 17012 36772 17013 36812
rect 16971 36763 17013 36772
rect 16972 36678 17012 36763
rect 17067 36644 17109 36653
rect 17067 36604 17068 36644
rect 17108 36604 17109 36644
rect 17067 36595 17109 36604
rect 16971 36560 17013 36569
rect 16971 36520 16972 36560
rect 17012 36520 17013 36560
rect 16971 36511 17013 36520
rect 16492 35008 16916 35048
rect 16492 32201 16532 35008
rect 16683 34880 16725 34889
rect 16683 34840 16684 34880
rect 16724 34840 16725 34880
rect 16683 34831 16725 34840
rect 16684 34469 16724 34831
rect 16875 34628 16917 34637
rect 16875 34588 16876 34628
rect 16916 34588 16917 34628
rect 16875 34579 16917 34588
rect 16876 34494 16916 34579
rect 16683 34460 16725 34469
rect 16683 34420 16684 34460
rect 16724 34420 16725 34460
rect 16683 34411 16725 34420
rect 16684 34326 16724 34411
rect 16972 34385 17012 36511
rect 16971 34376 17013 34385
rect 16971 34336 16972 34376
rect 17012 34336 17013 34376
rect 16971 34327 17013 34336
rect 17068 33032 17108 36595
rect 17260 36560 17300 37192
rect 17547 36980 17589 36989
rect 17547 36940 17548 36980
rect 17588 36940 17589 36980
rect 17547 36931 17589 36940
rect 17260 35720 17300 36520
rect 17355 35888 17397 35897
rect 17355 35848 17356 35888
rect 17396 35848 17397 35888
rect 17355 35839 17397 35848
rect 17260 35057 17300 35680
rect 17356 35300 17396 35839
rect 17548 35300 17588 36931
rect 18124 36905 18164 41971
rect 18700 41945 18740 42484
rect 19563 42475 19605 42484
rect 19660 42440 19700 42484
rect 19660 42400 19796 42440
rect 18808 42356 19176 42365
rect 18848 42316 18890 42356
rect 18930 42316 18972 42356
rect 19012 42316 19054 42356
rect 19094 42316 19136 42356
rect 18808 42307 19176 42316
rect 19276 42020 19316 42029
rect 19659 42020 19701 42029
rect 19316 41980 19604 42020
rect 19276 41971 19316 41980
rect 18699 41936 18741 41945
rect 18699 41896 18700 41936
rect 18740 41896 18741 41936
rect 18699 41887 18741 41896
rect 18987 41936 19029 41945
rect 18987 41896 18988 41936
rect 19028 41896 19029 41936
rect 18987 41887 19029 41896
rect 18988 41432 19028 41887
rect 19467 41768 19509 41777
rect 19467 41728 19468 41768
rect 19508 41728 19509 41768
rect 19467 41719 19509 41728
rect 19468 41634 19508 41719
rect 18988 41383 19028 41392
rect 19275 41180 19317 41189
rect 19275 41140 19276 41180
rect 19316 41140 19317 41180
rect 19275 41131 19317 41140
rect 19276 41046 19316 41131
rect 19467 41096 19509 41105
rect 19467 41056 19468 41096
rect 19508 41056 19509 41096
rect 19467 41047 19509 41056
rect 19468 40962 19508 41047
rect 19564 40928 19604 41980
rect 19659 41980 19660 42020
rect 19700 41980 19701 42020
rect 19659 41971 19701 41980
rect 19660 41886 19700 41971
rect 19660 41180 19700 41189
rect 19756 41180 19796 42400
rect 20524 42281 20564 44752
rect 20523 42272 20565 42281
rect 20523 42232 20524 42272
rect 20564 42232 20565 42272
rect 20523 42223 20565 42232
rect 19851 42104 19893 42113
rect 19851 42064 19852 42104
rect 19892 42064 19893 42104
rect 19851 42055 19893 42064
rect 19852 41970 19892 42055
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 19851 41432 19893 41441
rect 19851 41392 19852 41432
rect 19892 41392 19893 41432
rect 19851 41383 19893 41392
rect 19852 41298 19892 41383
rect 19700 41140 19796 41180
rect 19660 41131 19700 41140
rect 19564 40888 19796 40928
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 19371 40760 19413 40769
rect 19371 40720 19372 40760
rect 19412 40720 19413 40760
rect 19371 40711 19413 40720
rect 19563 40760 19605 40769
rect 19563 40720 19564 40760
rect 19604 40720 19605 40760
rect 19563 40711 19605 40720
rect 18988 40508 19028 40517
rect 18988 39920 19028 40468
rect 19372 40508 19412 40711
rect 19564 40676 19604 40711
rect 19564 40625 19604 40636
rect 19372 40459 19412 40468
rect 19180 40256 19220 40265
rect 19180 40013 19220 40216
rect 19179 40004 19221 40013
rect 19179 39964 19180 40004
rect 19220 39964 19221 40004
rect 19179 39955 19221 39964
rect 18988 39500 19028 39880
rect 19563 39836 19605 39845
rect 19563 39796 19564 39836
rect 19604 39796 19605 39836
rect 19563 39787 19605 39796
rect 19276 39668 19316 39677
rect 19316 39628 19412 39668
rect 19276 39619 19316 39628
rect 18700 39460 19028 39500
rect 18700 38912 18740 39460
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 18700 38753 18740 38872
rect 19276 38996 19316 39005
rect 19276 38837 19316 38956
rect 19275 38828 19317 38837
rect 19275 38788 19276 38828
rect 19316 38788 19317 38828
rect 19275 38779 19317 38788
rect 18699 38744 18741 38753
rect 18699 38704 18700 38744
rect 18740 38704 18741 38744
rect 18699 38695 18741 38704
rect 18987 38744 19029 38753
rect 18987 38704 18988 38744
rect 19028 38704 19029 38744
rect 18987 38695 19029 38704
rect 18988 38408 19028 38695
rect 18988 38359 19028 38368
rect 19276 38165 19316 38250
rect 18603 38156 18645 38165
rect 18603 38116 18604 38156
rect 18644 38116 18645 38156
rect 18603 38107 18645 38116
rect 19275 38156 19317 38165
rect 19275 38116 19276 38156
rect 19316 38116 19317 38156
rect 19275 38107 19317 38116
rect 18219 38072 18261 38081
rect 18219 38032 18220 38072
rect 18260 38032 18261 38072
rect 18219 38023 18261 38032
rect 18220 37913 18260 38023
rect 18604 38022 18644 38107
rect 19084 38072 19124 38081
rect 19124 38032 19220 38072
rect 19084 38023 19124 38032
rect 18796 37988 18836 37997
rect 18700 37948 18796 37988
rect 19180 37988 19220 38032
rect 19180 37948 19316 37988
rect 18219 37904 18261 37913
rect 18219 37864 18220 37904
rect 18260 37864 18261 37904
rect 18219 37855 18261 37864
rect 18603 37904 18645 37913
rect 18603 37864 18604 37904
rect 18644 37864 18645 37904
rect 18603 37855 18645 37864
rect 18123 36896 18165 36905
rect 18123 36856 18124 36896
rect 18164 36856 18165 36896
rect 18123 36847 18165 36856
rect 18219 36812 18261 36821
rect 18219 36772 18220 36812
rect 18260 36772 18261 36812
rect 18219 36763 18261 36772
rect 18123 35972 18165 35981
rect 18123 35932 18124 35972
rect 18164 35932 18165 35972
rect 18123 35923 18165 35932
rect 17356 35260 17492 35300
rect 17259 35048 17301 35057
rect 17259 35008 17260 35048
rect 17300 35008 17301 35048
rect 17259 34999 17301 35008
rect 17260 34914 17300 34999
rect 17163 34460 17205 34469
rect 17163 34420 17164 34460
rect 17204 34420 17205 34460
rect 17163 34411 17205 34420
rect 17164 33704 17204 34411
rect 17164 33655 17204 33664
rect 17259 33284 17301 33293
rect 17259 33244 17260 33284
rect 17300 33244 17301 33284
rect 17259 33235 17301 33244
rect 16588 32992 17108 33032
rect 16491 32192 16533 32201
rect 16491 32152 16492 32192
rect 16532 32152 16533 32192
rect 16491 32143 16533 32152
rect 16300 31564 16436 31604
rect 16203 31520 16245 31529
rect 16203 31480 16204 31520
rect 16244 31480 16245 31520
rect 16203 31471 16245 31480
rect 16203 30680 16245 30689
rect 16203 30640 16204 30680
rect 16244 30640 16245 30680
rect 16300 30680 16340 31564
rect 16395 31100 16437 31109
rect 16395 31060 16396 31100
rect 16436 31060 16437 31100
rect 16395 31051 16437 31060
rect 16396 30848 16436 31051
rect 16396 30799 16436 30808
rect 16300 30640 16436 30680
rect 16203 30631 16245 30640
rect 16204 30521 16244 30631
rect 16203 30512 16245 30521
rect 16203 30472 16204 30512
rect 16244 30472 16245 30512
rect 16203 30463 16245 30472
rect 15819 30008 15861 30017
rect 15819 29968 15820 30008
rect 15860 29968 15861 30008
rect 15819 29959 15861 29968
rect 16299 30008 16341 30017
rect 16299 29968 16300 30008
rect 16340 29968 16341 30008
rect 16299 29959 16341 29968
rect 15820 29845 15860 29854
rect 15723 29672 15765 29681
rect 15723 29632 15724 29672
rect 15764 29632 15765 29672
rect 15723 29623 15765 29632
rect 15820 29513 15860 29805
rect 15915 29840 15957 29849
rect 15915 29800 15916 29840
rect 15956 29800 15957 29840
rect 15915 29791 15957 29800
rect 15819 29504 15861 29513
rect 15819 29464 15820 29504
rect 15860 29464 15861 29504
rect 15819 29455 15861 29464
rect 15916 29420 15956 29791
rect 16012 29672 16052 29681
rect 16052 29632 16244 29672
rect 16012 29623 16052 29632
rect 15916 29380 16052 29420
rect 15628 29287 15668 29296
rect 15915 29168 15957 29177
rect 15915 29128 15916 29168
rect 15956 29128 15957 29168
rect 15915 29119 15957 29128
rect 15724 29000 15764 29009
rect 15627 28664 15669 28673
rect 15627 28624 15628 28664
rect 15668 28624 15669 28664
rect 15627 28615 15669 28624
rect 15628 28496 15668 28615
rect 15628 28447 15668 28456
rect 15531 27656 15573 27665
rect 15531 27616 15532 27656
rect 15572 27616 15573 27656
rect 15531 27607 15573 27616
rect 15724 27488 15764 28960
rect 15916 28580 15956 29119
rect 15916 28531 15956 28540
rect 15819 27824 15861 27833
rect 15819 27784 15820 27824
rect 15860 27784 15861 27824
rect 15819 27775 15861 27784
rect 15435 27236 15477 27245
rect 15435 27196 15436 27236
rect 15476 27196 15477 27236
rect 15435 27187 15477 27196
rect 15436 27068 15476 27187
rect 15436 27019 15476 27028
rect 15628 26648 15668 26657
rect 15724 26648 15764 27448
rect 15820 26816 15860 27775
rect 16012 27740 16052 29380
rect 16108 28337 16148 28422
rect 16107 28328 16149 28337
rect 16107 28288 16108 28328
rect 16148 28288 16149 28328
rect 16107 28279 16149 28288
rect 16107 28160 16149 28169
rect 16107 28120 16108 28160
rect 16148 28120 16149 28160
rect 16107 28111 16149 28120
rect 16012 27691 16052 27700
rect 15916 27656 15956 27665
rect 15916 27497 15956 27616
rect 16108 27656 16148 28111
rect 16108 27607 16148 27616
rect 15915 27488 15957 27497
rect 15915 27448 15916 27488
rect 15956 27448 15957 27488
rect 15915 27439 15957 27448
rect 16204 27413 16244 29632
rect 16300 29345 16340 29959
rect 16299 29336 16341 29345
rect 16299 29296 16300 29336
rect 16340 29296 16341 29336
rect 16299 29287 16341 29296
rect 16203 27404 16245 27413
rect 16203 27364 16204 27404
rect 16244 27364 16245 27404
rect 16203 27355 16245 27364
rect 16300 26984 16340 29287
rect 16204 26944 16340 26984
rect 15820 26776 16052 26816
rect 15916 26648 15956 26657
rect 15668 26608 15916 26648
rect 15628 26144 15668 26608
rect 15916 26599 15956 26608
rect 15723 26228 15765 26237
rect 15723 26188 15724 26228
rect 15764 26188 15765 26228
rect 15723 26179 15765 26188
rect 15340 25936 15572 25976
rect 15244 25892 15284 25901
rect 15284 25852 15380 25892
rect 15244 25843 15284 25852
rect 15147 25556 15189 25565
rect 15147 25516 15148 25556
rect 15188 25516 15189 25556
rect 15147 25507 15189 25516
rect 15148 25304 15188 25507
rect 15244 25304 15284 25313
rect 15148 25264 15244 25304
rect 14860 24632 14900 24641
rect 14763 24548 14805 24557
rect 14763 24508 14764 24548
rect 14804 24508 14805 24548
rect 14763 24499 14805 24508
rect 14764 24414 14804 24499
rect 14860 24473 14900 24592
rect 14859 24464 14901 24473
rect 14859 24424 14860 24464
rect 14900 24424 14901 24464
rect 14859 24415 14901 24424
rect 15148 24380 15188 25264
rect 15244 25255 15284 25264
rect 15243 24716 15285 24725
rect 15243 24676 15244 24716
rect 15284 24676 15285 24716
rect 15243 24667 15285 24676
rect 15244 24548 15284 24667
rect 15244 24499 15284 24508
rect 15148 24340 15284 24380
rect 14668 24172 14900 24212
rect 14475 23792 14517 23801
rect 14475 23752 14476 23792
rect 14516 23752 14517 23792
rect 14475 23743 14517 23752
rect 14476 23658 14516 23743
rect 14668 23624 14708 23633
rect 14475 23288 14517 23297
rect 14475 23248 14476 23288
rect 14516 23248 14517 23288
rect 14475 23239 14517 23248
rect 14476 22541 14516 23239
rect 14668 23115 14708 23584
rect 14860 23288 14900 24172
rect 15147 23960 15189 23969
rect 15147 23920 15148 23960
rect 15188 23920 15189 23960
rect 15147 23911 15189 23920
rect 14860 23239 14900 23248
rect 14668 23066 14708 23075
rect 15148 22784 15188 23911
rect 15244 23633 15284 24340
rect 15340 23969 15380 25852
rect 15435 25220 15477 25229
rect 15435 25180 15436 25220
rect 15476 25180 15477 25220
rect 15435 25171 15477 25180
rect 15436 25086 15476 25171
rect 15435 24800 15477 24809
rect 15435 24760 15436 24800
rect 15476 24760 15477 24800
rect 15435 24751 15477 24760
rect 15436 24666 15476 24751
rect 15339 23960 15381 23969
rect 15339 23920 15340 23960
rect 15380 23920 15381 23960
rect 15339 23911 15381 23920
rect 15243 23624 15285 23633
rect 15243 23584 15244 23624
rect 15284 23584 15285 23624
rect 15243 23575 15285 23584
rect 15243 23036 15285 23045
rect 15243 22996 15244 23036
rect 15284 22996 15285 23036
rect 15243 22987 15285 22996
rect 15244 22902 15284 22987
rect 15436 22868 15476 22877
rect 15148 22744 15284 22784
rect 14475 22532 14517 22541
rect 14475 22492 14476 22532
rect 14516 22492 14517 22532
rect 14475 22483 14517 22492
rect 15147 22532 15189 22541
rect 15147 22492 15148 22532
rect 15188 22492 15189 22532
rect 15147 22483 15189 22492
rect 14572 22289 14612 22374
rect 14379 22280 14421 22289
rect 14379 22240 14380 22280
rect 14420 22240 14421 22280
rect 14379 22231 14421 22240
rect 14571 22280 14613 22289
rect 14571 22240 14572 22280
rect 14612 22240 14613 22280
rect 14571 22231 14613 22240
rect 14763 22280 14805 22289
rect 14763 22240 14764 22280
rect 14804 22240 14805 22280
rect 14763 22231 14805 22240
rect 14860 22280 14900 22289
rect 14764 22146 14804 22231
rect 14380 22112 14420 22121
rect 14668 22112 14708 22121
rect 14283 21944 14325 21953
rect 14283 21904 14284 21944
rect 14324 21904 14325 21944
rect 14283 21895 14325 21904
rect 14188 21820 14231 21860
rect 14091 21811 14133 21820
rect 14191 21776 14231 21820
rect 14188 21736 14231 21776
rect 14283 21776 14325 21785
rect 14283 21736 14284 21776
rect 14324 21736 14325 21776
rect 13996 21692 14036 21701
rect 14188 21692 14228 21736
rect 14283 21727 14325 21736
rect 14036 21652 14228 21692
rect 13996 21643 14036 21652
rect 14284 21608 14324 21727
rect 14188 21568 14324 21608
rect 13900 20140 14036 20180
rect 13707 20012 13749 20021
rect 13707 19972 13708 20012
rect 13748 19972 13749 20012
rect 13707 19963 13749 19972
rect 13516 19720 13652 19760
rect 13324 19207 13364 19216
rect 13420 19256 13460 19265
rect 12939 19088 12981 19097
rect 12939 19048 12940 19088
rect 12980 19048 12981 19088
rect 12939 19039 12981 19048
rect 13132 19088 13172 19097
rect 13420 19088 13460 19216
rect 13172 19048 13460 19088
rect 13132 19039 13172 19048
rect 12843 18332 12885 18341
rect 12843 18292 12844 18332
rect 12884 18292 12885 18332
rect 12843 18283 12885 18292
rect 12844 18198 12884 18283
rect 12843 17912 12885 17921
rect 12843 17872 12844 17912
rect 12884 17872 12885 17912
rect 12843 17863 12885 17872
rect 12844 17778 12884 17863
rect 12940 17744 12980 19039
rect 13516 19004 13556 19720
rect 13708 19349 13748 19963
rect 13707 19340 13749 19349
rect 13707 19300 13708 19340
rect 13748 19300 13749 19340
rect 13707 19291 13749 19300
rect 13612 19256 13652 19265
rect 13612 19097 13652 19216
rect 13708 19256 13748 19291
rect 13708 19206 13748 19216
rect 13809 19256 13849 19265
rect 13611 19088 13653 19097
rect 13611 19048 13612 19088
rect 13652 19048 13653 19088
rect 13611 19039 13653 19048
rect 13708 19088 13748 19097
rect 13420 18964 13556 19004
rect 13323 18920 13365 18929
rect 13323 18880 13324 18920
rect 13364 18880 13365 18920
rect 13323 18871 13365 18880
rect 13227 18584 13269 18593
rect 13227 18544 13228 18584
rect 13268 18544 13269 18584
rect 13227 18535 13269 18544
rect 13228 18257 13268 18535
rect 13227 18248 13269 18257
rect 13227 18208 13228 18248
rect 13268 18208 13269 18248
rect 13227 18199 13269 18208
rect 13324 18080 13364 18871
rect 12933 17704 12980 17744
rect 13084 18040 13364 18080
rect 13084 17755 13124 18040
rect 13324 17759 13364 17768
rect 13084 17706 13124 17715
rect 13228 17744 13268 17753
rect 12933 17660 12973 17704
rect 13228 17669 13268 17704
rect 13321 17719 13324 17759
rect 13321 17710 13364 17719
rect 13227 17660 13269 17669
rect 12933 17620 12980 17660
rect 12556 17023 12596 17032
rect 12652 17536 12788 17576
rect 12652 12797 12692 17536
rect 12940 17417 12980 17620
rect 13227 17620 13228 17660
rect 13268 17620 13269 17660
rect 13321 17660 13361 17710
rect 13321 17620 13364 17660
rect 13227 17611 13269 17620
rect 13131 17576 13173 17585
rect 13131 17536 13132 17576
rect 13172 17536 13173 17576
rect 13131 17527 13173 17536
rect 13132 17442 13172 17527
rect 12939 17408 12981 17417
rect 12939 17368 12940 17408
rect 12980 17368 12981 17408
rect 12939 17359 12981 17368
rect 13132 17165 13172 17187
rect 12748 17156 12788 17165
rect 13131 17156 13173 17165
rect 12788 17116 13076 17156
rect 12748 17107 12788 17116
rect 13036 17072 13076 17116
rect 13131 17116 13132 17156
rect 13172 17116 13173 17156
rect 13131 17107 13173 17116
rect 13132 17092 13172 17107
rect 13132 17043 13172 17052
rect 13036 17023 13076 17032
rect 13228 16988 13268 17611
rect 13132 16948 13268 16988
rect 13132 16904 13172 16948
rect 13324 16904 13364 17620
rect 12844 16864 13172 16904
rect 13228 16864 13364 16904
rect 12844 16232 12884 16864
rect 13228 16400 13268 16864
rect 13420 16736 13460 18964
rect 13708 18089 13748 19048
rect 13809 18929 13849 19216
rect 13803 18920 13849 18929
rect 13803 18880 13804 18920
rect 13844 18880 13849 18920
rect 13803 18871 13845 18880
rect 13899 18332 13941 18341
rect 13899 18292 13900 18332
rect 13940 18292 13941 18332
rect 13899 18283 13941 18292
rect 13707 18080 13749 18089
rect 13707 18040 13708 18080
rect 13748 18040 13749 18080
rect 13707 18031 13749 18040
rect 13515 17912 13557 17921
rect 13804 17912 13844 17921
rect 13515 17872 13516 17912
rect 13556 17872 13557 17912
rect 13515 17863 13557 17872
rect 13612 17872 13804 17912
rect 13516 17744 13556 17863
rect 13516 17576 13556 17704
rect 13612 17744 13652 17872
rect 13804 17863 13844 17872
rect 13900 17753 13940 18283
rect 13612 17695 13652 17704
rect 13804 17744 13844 17753
rect 13804 17660 13844 17704
rect 13899 17744 13941 17753
rect 13899 17704 13900 17744
rect 13940 17704 13941 17744
rect 13899 17695 13941 17704
rect 13708 17620 13844 17660
rect 13708 17576 13748 17620
rect 13516 17536 13748 17576
rect 13515 17408 13557 17417
rect 13515 17368 13516 17408
rect 13556 17368 13557 17408
rect 13515 17359 13557 17368
rect 13516 16997 13556 17359
rect 13707 17240 13749 17249
rect 13707 17200 13708 17240
rect 13748 17200 13749 17240
rect 13707 17191 13749 17200
rect 13515 16988 13557 16997
rect 13515 16948 13516 16988
rect 13556 16948 13557 16988
rect 13515 16939 13557 16948
rect 13612 16988 13652 16997
rect 13516 16854 13556 16939
rect 13612 16745 13652 16948
rect 13611 16736 13653 16745
rect 13420 16696 13556 16736
rect 13132 16360 13268 16400
rect 12844 16183 12884 16192
rect 12940 16232 12980 16243
rect 12940 16157 12980 16192
rect 12939 16148 12981 16157
rect 12939 16108 12940 16148
rect 12980 16108 12981 16148
rect 12939 16099 12981 16108
rect 13035 16064 13077 16073
rect 13035 16024 13036 16064
rect 13076 16024 13077 16064
rect 13035 16015 13077 16024
rect 13132 16064 13172 16360
rect 13132 16015 13172 16024
rect 13420 16232 13460 16241
rect 13036 15653 13076 16015
rect 13035 15644 13077 15653
rect 13035 15604 13036 15644
rect 13076 15604 13077 15644
rect 13035 15595 13077 15604
rect 12843 15560 12885 15569
rect 12843 15520 12844 15560
rect 12884 15520 12885 15560
rect 12843 15511 12885 15520
rect 12747 15224 12789 15233
rect 12747 15184 12748 15224
rect 12788 15184 12789 15224
rect 12747 15175 12789 15184
rect 12651 12788 12693 12797
rect 12651 12748 12652 12788
rect 12692 12748 12693 12788
rect 12651 12739 12693 12748
rect 12556 12620 12596 12629
rect 12596 12580 12692 12620
rect 12556 12571 12596 12580
rect 12555 12452 12597 12461
rect 12555 12412 12556 12452
rect 12596 12412 12597 12452
rect 12555 12403 12597 12412
rect 12556 10193 12596 12403
rect 12652 10361 12692 12580
rect 12748 11285 12788 15175
rect 12844 15149 12884 15511
rect 13420 15392 13460 16192
rect 13036 15308 13076 15317
rect 12940 15268 13036 15308
rect 12843 15140 12885 15149
rect 12843 15100 12844 15140
rect 12884 15100 12885 15140
rect 12843 15091 12885 15100
rect 12843 14048 12885 14057
rect 12843 14008 12844 14048
rect 12884 14008 12885 14048
rect 12940 14048 12980 15268
rect 13036 15259 13076 15268
rect 13420 15065 13460 15352
rect 13419 15056 13461 15065
rect 13419 15016 13420 15056
rect 13460 15016 13461 15056
rect 13419 15007 13461 15016
rect 13516 14981 13556 16696
rect 13611 16696 13612 16736
rect 13652 16696 13653 16736
rect 13611 16687 13653 16696
rect 13708 16568 13748 17191
rect 13803 17156 13845 17165
rect 13803 17116 13804 17156
rect 13844 17116 13845 17156
rect 13803 17107 13845 17116
rect 13612 16528 13748 16568
rect 13515 14972 13557 14981
rect 13515 14932 13516 14972
rect 13556 14932 13557 14972
rect 13515 14923 13557 14932
rect 13612 14813 13652 16528
rect 13707 16400 13749 16409
rect 13707 16360 13708 16400
rect 13748 16360 13749 16400
rect 13707 16351 13749 16360
rect 13708 15560 13748 16351
rect 13708 15511 13748 15520
rect 13611 14804 13653 14813
rect 13611 14764 13612 14804
rect 13652 14764 13653 14804
rect 13611 14755 13653 14764
rect 13420 14720 13460 14729
rect 13036 14680 13420 14720
rect 13036 14216 13076 14680
rect 13420 14671 13460 14680
rect 13516 14720 13556 14729
rect 13036 14167 13076 14176
rect 13420 14048 13460 14057
rect 12940 14008 13420 14048
rect 12843 13999 12885 14008
rect 13420 13999 13460 14008
rect 13516 14048 13556 14680
rect 13556 14008 13652 14048
rect 13516 13999 13556 14008
rect 12844 12461 12884 13999
rect 13131 13796 13173 13805
rect 13131 13756 13132 13796
rect 13172 13756 13173 13796
rect 13131 13747 13173 13756
rect 12940 13208 12980 13219
rect 12940 13133 12980 13168
rect 13036 13208 13076 13217
rect 13132 13208 13172 13747
rect 13516 13217 13556 13302
rect 13076 13168 13172 13208
rect 13036 13159 13076 13168
rect 12939 13124 12981 13133
rect 12939 13084 12940 13124
rect 12980 13084 12981 13124
rect 12939 13075 12981 13084
rect 12939 12620 12981 12629
rect 12939 12580 12940 12620
rect 12980 12580 12981 12620
rect 12939 12571 12981 12580
rect 12843 12452 12885 12461
rect 12843 12412 12844 12452
rect 12884 12412 12885 12452
rect 12843 12403 12885 12412
rect 12940 12041 12980 12571
rect 13035 12536 13077 12545
rect 13035 12496 13036 12536
rect 13076 12496 13077 12536
rect 13035 12487 13077 12496
rect 13036 12125 13076 12487
rect 13035 12116 13077 12125
rect 13035 12076 13036 12116
rect 13076 12076 13077 12116
rect 13035 12067 13077 12076
rect 12939 12032 12981 12041
rect 12939 11992 12940 12032
rect 12980 11992 12981 12032
rect 12939 11983 12981 11992
rect 12939 11360 12981 11369
rect 12939 11320 12940 11360
rect 12980 11320 12981 11360
rect 12939 11311 12981 11320
rect 12747 11276 12789 11285
rect 12747 11236 12748 11276
rect 12788 11236 12789 11276
rect 12747 11227 12789 11236
rect 12747 11108 12789 11117
rect 12747 11068 12748 11108
rect 12788 11068 12789 11108
rect 12747 11059 12789 11068
rect 12651 10352 12693 10361
rect 12651 10312 12652 10352
rect 12692 10312 12693 10352
rect 12651 10303 12693 10312
rect 12555 10184 12597 10193
rect 12555 10144 12556 10184
rect 12596 10144 12597 10184
rect 12555 10135 12597 10144
rect 12652 10184 12692 10193
rect 12748 10184 12788 11059
rect 12844 11010 12884 11019
rect 12844 10436 12884 10970
rect 12844 10387 12884 10396
rect 12940 10268 12980 11311
rect 13036 11285 13076 11329
rect 13035 11276 13077 11285
rect 13035 11236 13036 11276
rect 13076 11236 13077 11276
rect 13035 11234 13077 11236
rect 13035 11227 13036 11234
rect 13076 11227 13077 11234
rect 13036 11185 13076 11194
rect 13132 11192 13172 13168
rect 13420 13208 13460 13217
rect 13420 11369 13460 13168
rect 13515 13208 13557 13217
rect 13515 13168 13516 13208
rect 13556 13168 13557 13208
rect 13515 13159 13557 13168
rect 13612 13040 13652 14008
rect 13516 13000 13652 13040
rect 13419 11360 13461 11369
rect 13419 11320 13420 11360
rect 13460 11320 13461 11360
rect 13419 11311 13461 11320
rect 13132 11152 13460 11192
rect 13324 11024 13364 11033
rect 12692 10144 12788 10184
rect 12844 10228 12980 10268
rect 13132 10984 13324 11024
rect 12652 10135 12692 10144
rect 12459 9512 12501 9521
rect 12459 9472 12460 9512
rect 12500 9472 12501 9512
rect 12459 9463 12501 9472
rect 12556 9185 12596 10135
rect 12555 9176 12597 9185
rect 12555 9136 12556 9176
rect 12596 9136 12597 9176
rect 12555 9127 12597 9136
rect 12459 8672 12501 8681
rect 12116 7960 12212 8000
rect 12268 8632 12460 8672
rect 12500 8632 12501 8672
rect 12076 6833 12116 7960
rect 12172 7160 12212 7169
rect 12268 7160 12308 8632
rect 12459 8623 12501 8632
rect 12460 8538 12500 8623
rect 12652 8504 12692 8513
rect 12459 8420 12501 8429
rect 12459 8380 12460 8420
rect 12500 8380 12501 8420
rect 12459 8371 12501 8380
rect 12363 7328 12405 7337
rect 12363 7288 12364 7328
rect 12404 7288 12405 7328
rect 12363 7279 12405 7288
rect 12364 7194 12404 7279
rect 12212 7120 12308 7160
rect 12075 6824 12117 6833
rect 12075 6784 12076 6824
rect 12116 6784 12117 6824
rect 12075 6775 12117 6784
rect 12172 6497 12212 7120
rect 12171 6488 12213 6497
rect 12171 6448 12172 6488
rect 12212 6448 12213 6488
rect 12171 6439 12213 6448
rect 12075 6320 12117 6329
rect 12075 6280 12076 6320
rect 12116 6280 12117 6320
rect 12075 6271 12117 6280
rect 12076 5153 12116 6271
rect 12460 5573 12500 8371
rect 12652 8000 12692 8464
rect 12747 8084 12789 8093
rect 12747 8044 12748 8084
rect 12788 8044 12789 8084
rect 12747 8035 12789 8044
rect 12604 7990 12692 8000
rect 12644 7960 12692 7990
rect 12748 7950 12788 8035
rect 12604 7941 12644 7950
rect 12651 7328 12693 7337
rect 12651 7288 12652 7328
rect 12692 7288 12693 7328
rect 12651 7279 12693 7288
rect 12652 7160 12692 7279
rect 12652 7111 12692 7120
rect 12747 7160 12789 7169
rect 12747 7120 12748 7160
rect 12788 7120 12789 7160
rect 12747 7111 12789 7120
rect 12748 6992 12788 7111
rect 12652 6952 12788 6992
rect 12459 5564 12501 5573
rect 12459 5524 12460 5564
rect 12500 5524 12501 5564
rect 12459 5515 12501 5524
rect 12075 5144 12117 5153
rect 12075 5104 12076 5144
rect 12116 5104 12117 5144
rect 12075 5095 12117 5104
rect 11979 2792 12021 2801
rect 11979 2752 11980 2792
rect 12020 2752 12021 2792
rect 11979 2743 12021 2752
rect 11788 2500 11924 2540
rect 11500 1819 11540 1828
rect 11596 2456 11636 2465
rect 11116 1700 11156 1709
rect 11307 1700 11349 1709
rect 11156 1660 11252 1700
rect 11116 1651 11156 1660
rect 11116 1196 11156 1205
rect 11020 1156 11116 1196
rect 11116 1147 11156 1156
rect 11212 1121 11252 1660
rect 11307 1660 11308 1700
rect 11348 1660 11349 1700
rect 11307 1651 11349 1660
rect 11308 1566 11348 1651
rect 11596 1364 11636 2416
rect 11884 2381 11924 2500
rect 11883 2372 11925 2381
rect 11883 2332 11884 2372
rect 11924 2332 11925 2372
rect 11883 2323 11925 2332
rect 11691 1868 11733 1877
rect 11691 1828 11692 1868
rect 11732 1828 11733 1868
rect 11691 1819 11733 1828
rect 12075 1868 12117 1877
rect 12075 1828 12076 1868
rect 12116 1828 12117 1868
rect 12075 1819 12117 1828
rect 11692 1734 11732 1819
rect 12076 1734 12116 1819
rect 11884 1700 11924 1709
rect 11884 1373 11924 1660
rect 12268 1700 12308 1709
rect 12308 1660 12404 1700
rect 12268 1651 12308 1660
rect 11883 1364 11925 1373
rect 11596 1324 11732 1364
rect 11595 1196 11637 1205
rect 11595 1156 11596 1196
rect 11636 1156 11637 1196
rect 11595 1147 11637 1156
rect 11211 1112 11253 1121
rect 11211 1072 11212 1112
rect 11252 1072 11253 1112
rect 11211 1063 11253 1072
rect 11596 1062 11636 1147
rect 11211 944 11253 953
rect 11211 904 11212 944
rect 11252 904 11253 944
rect 11211 895 11253 904
rect 11308 944 11348 953
rect 11692 944 11732 1324
rect 11883 1324 11884 1364
rect 11924 1324 11925 1364
rect 11883 1315 11925 1324
rect 12171 1280 12213 1289
rect 12171 1240 12172 1280
rect 12212 1240 12213 1280
rect 12171 1231 12213 1240
rect 11979 1112 12021 1121
rect 11979 1072 11980 1112
rect 12020 1072 12021 1112
rect 11979 1063 12021 1072
rect 11348 904 11444 944
rect 11308 895 11348 904
rect 11019 776 11061 785
rect 11019 736 11020 776
rect 11060 736 11061 776
rect 11019 727 11061 736
rect 11020 80 11060 727
rect 11212 80 11252 895
rect 11404 80 11444 904
rect 11596 904 11732 944
rect 11788 944 11828 953
rect 11596 80 11636 904
rect 11788 80 11828 904
rect 11980 80 12020 1063
rect 12172 80 12212 1231
rect 12364 80 12404 1660
rect 12555 1028 12597 1037
rect 12555 988 12556 1028
rect 12596 988 12597 1028
rect 12555 979 12597 988
rect 12556 80 12596 979
rect 12652 785 12692 6952
rect 12748 6488 12788 6497
rect 12844 6488 12884 10228
rect 13035 10016 13077 10025
rect 13035 9976 13036 10016
rect 13076 9976 13077 10016
rect 13035 9967 13077 9976
rect 12940 9605 12980 9636
rect 12939 9596 12981 9605
rect 12939 9556 12940 9596
rect 12980 9556 12981 9596
rect 12939 9547 12981 9556
rect 12940 9512 12980 9547
rect 12940 8681 12980 9472
rect 12939 8672 12981 8681
rect 12939 8632 12940 8672
rect 12980 8632 12981 8672
rect 12939 8623 12981 8632
rect 12939 8420 12981 8429
rect 12939 8380 12940 8420
rect 12980 8380 12981 8420
rect 12939 8371 12981 8380
rect 12788 6448 12884 6488
rect 12748 6439 12788 6448
rect 12747 5060 12789 5069
rect 12747 5020 12748 5060
rect 12788 5020 12789 5060
rect 12747 5011 12789 5020
rect 12748 1868 12788 5011
rect 12940 3137 12980 8371
rect 13036 3893 13076 9967
rect 13132 9680 13172 10984
rect 13324 10975 13364 10984
rect 13420 11024 13460 11152
rect 13227 10856 13269 10865
rect 13227 10816 13228 10856
rect 13268 10816 13269 10856
rect 13227 10807 13269 10816
rect 13132 9631 13172 9640
rect 13131 7244 13173 7253
rect 13131 7204 13132 7244
rect 13172 7204 13173 7244
rect 13131 7195 13173 7204
rect 13228 7244 13268 10807
rect 13323 10772 13365 10781
rect 13323 10732 13324 10772
rect 13364 10732 13365 10772
rect 13323 10723 13365 10732
rect 13324 10184 13364 10723
rect 13324 10135 13364 10144
rect 13324 8672 13364 8681
rect 13324 8513 13364 8632
rect 13323 8504 13365 8513
rect 13323 8464 13324 8504
rect 13364 8464 13365 8504
rect 13323 8455 13365 8464
rect 13420 8177 13460 10984
rect 13516 10025 13556 13000
rect 13804 12956 13844 17107
rect 13996 14897 14036 20140
rect 14188 19517 14228 21568
rect 14380 20180 14420 22072
rect 14476 22072 14668 22112
rect 14476 21608 14516 22072
rect 14668 22063 14708 22072
rect 14667 21944 14709 21953
rect 14667 21904 14668 21944
rect 14708 21904 14709 21944
rect 14667 21895 14709 21904
rect 14571 21860 14613 21869
rect 14571 21820 14572 21860
rect 14612 21820 14613 21860
rect 14571 21811 14613 21820
rect 14476 21559 14516 21568
rect 14572 21608 14612 21811
rect 14668 21776 14708 21895
rect 14860 21776 14900 22240
rect 15051 22280 15093 22289
rect 15051 22240 15052 22280
rect 15092 22240 15093 22280
rect 15051 22231 15093 22240
rect 15148 22280 15188 22483
rect 14668 21727 14708 21736
rect 14764 21736 14900 21776
rect 14572 21559 14612 21568
rect 14764 21608 14804 21736
rect 15052 21617 15092 22231
rect 14764 21020 14804 21568
rect 14859 21608 14901 21617
rect 14859 21568 14860 21608
rect 14900 21568 14901 21608
rect 14859 21559 14901 21568
rect 15015 21608 15092 21617
rect 15055 21568 15092 21608
rect 15015 21559 15092 21568
rect 14860 21474 14900 21559
rect 14860 21020 14900 21029
rect 14764 20980 14860 21020
rect 14860 20971 14900 20980
rect 14668 20768 14708 20777
rect 14475 20684 14517 20693
rect 14475 20644 14476 20684
rect 14516 20644 14517 20684
rect 14475 20635 14517 20644
rect 14284 20140 14420 20180
rect 14187 19508 14229 19517
rect 14187 19468 14188 19508
rect 14228 19468 14229 19508
rect 14187 19459 14229 19468
rect 14091 19340 14133 19349
rect 14091 19300 14092 19340
rect 14132 19300 14133 19340
rect 14091 19291 14133 19300
rect 14092 19256 14132 19291
rect 14092 19205 14132 19216
rect 14188 19256 14228 19267
rect 14188 19181 14228 19216
rect 14187 19172 14229 19181
rect 14187 19132 14188 19172
rect 14228 19132 14229 19172
rect 14187 19123 14229 19132
rect 14284 18920 14324 20140
rect 14379 19088 14421 19097
rect 14379 19048 14380 19088
rect 14420 19048 14421 19088
rect 14379 19039 14421 19048
rect 14380 18954 14420 19039
rect 14188 18880 14324 18920
rect 14092 17744 14132 17753
rect 14092 17417 14132 17704
rect 14091 17408 14133 17417
rect 14091 17368 14092 17408
rect 14132 17368 14133 17408
rect 14091 17359 14133 17368
rect 14091 17240 14133 17249
rect 14091 17200 14092 17240
rect 14132 17200 14133 17240
rect 14091 17191 14133 17200
rect 14092 17072 14132 17191
rect 14092 15737 14132 17032
rect 14091 15728 14133 15737
rect 14091 15688 14092 15728
rect 14132 15688 14133 15728
rect 14091 15679 14133 15688
rect 14091 14972 14133 14981
rect 14091 14932 14092 14972
rect 14132 14932 14133 14972
rect 14091 14923 14133 14932
rect 13995 14888 14037 14897
rect 13995 14848 13996 14888
rect 14036 14848 14037 14888
rect 13995 14839 14037 14848
rect 13900 14720 13940 14729
rect 13900 13964 13940 14680
rect 13996 14720 14036 14729
rect 14092 14720 14132 14923
rect 14036 14680 14132 14720
rect 13996 14671 14036 14680
rect 13900 13721 13940 13924
rect 13996 13964 14036 13973
rect 13899 13712 13941 13721
rect 13899 13672 13900 13712
rect 13940 13672 13941 13712
rect 13899 13663 13941 13672
rect 13996 13376 14036 13924
rect 13612 12916 13844 12956
rect 13900 13336 14036 13376
rect 13515 10016 13557 10025
rect 13515 9976 13516 10016
rect 13556 9976 13557 10016
rect 13515 9967 13557 9976
rect 13612 9857 13652 12916
rect 13707 12788 13749 12797
rect 13707 12748 13708 12788
rect 13748 12748 13749 12788
rect 13707 12739 13749 12748
rect 13611 9848 13653 9857
rect 13611 9808 13612 9848
rect 13652 9808 13653 9848
rect 13611 9799 13653 9808
rect 13708 9680 13748 12739
rect 13900 11864 13940 13336
rect 13995 13208 14037 13217
rect 13995 13168 13996 13208
rect 14036 13168 14037 13208
rect 13995 13159 14037 13168
rect 13996 13074 14036 13159
rect 13995 12704 14037 12713
rect 13995 12664 13996 12704
rect 14036 12664 14037 12704
rect 13995 12655 14037 12664
rect 13804 11824 13940 11864
rect 13804 11285 13844 11824
rect 13900 11696 13940 11705
rect 13996 11696 14036 12655
rect 13940 11656 14036 11696
rect 13900 11453 13940 11656
rect 13899 11444 13941 11453
rect 13899 11404 13900 11444
rect 13940 11404 13941 11444
rect 13899 11395 13941 11404
rect 14188 11360 14228 18880
rect 14476 18836 14516 20635
rect 14668 20096 14708 20728
rect 14956 20264 14996 20273
rect 15052 20264 15092 21559
rect 15148 20768 15188 22240
rect 15244 21860 15284 22744
rect 15436 22289 15476 22828
rect 15435 22280 15477 22289
rect 15435 22240 15436 22280
rect 15476 22240 15477 22280
rect 15435 22231 15477 22240
rect 15339 22112 15381 22121
rect 15339 22072 15340 22112
rect 15380 22072 15381 22112
rect 15339 22063 15381 22072
rect 15340 21978 15380 22063
rect 15532 21944 15572 25936
rect 15628 25136 15668 26104
rect 15628 24464 15668 25096
rect 15724 24809 15764 26179
rect 15819 25892 15861 25901
rect 15819 25852 15820 25892
rect 15860 25852 15861 25892
rect 15819 25843 15861 25852
rect 15723 24800 15765 24809
rect 15723 24760 15724 24800
rect 15764 24760 15765 24800
rect 15723 24751 15765 24760
rect 15723 24632 15765 24641
rect 15723 24592 15724 24632
rect 15764 24592 15765 24632
rect 15723 24583 15765 24592
rect 15628 23624 15668 24424
rect 15628 22952 15668 23584
rect 15628 22121 15668 22912
rect 15724 23792 15764 24583
rect 15820 24053 15860 25843
rect 16012 25304 16052 26776
rect 15916 25264 16012 25304
rect 15916 24809 15956 25264
rect 16012 25255 16052 25264
rect 16011 25136 16053 25145
rect 16011 25096 16012 25136
rect 16052 25096 16053 25136
rect 16011 25087 16053 25096
rect 15915 24800 15957 24809
rect 15915 24760 15916 24800
rect 15956 24760 15957 24800
rect 15915 24751 15957 24760
rect 16012 24632 16052 25087
rect 16107 24884 16149 24893
rect 16107 24844 16108 24884
rect 16148 24844 16149 24884
rect 16107 24835 16149 24844
rect 15916 24592 16012 24632
rect 15819 24044 15861 24053
rect 15819 24004 15820 24044
rect 15860 24004 15861 24044
rect 15819 23995 15861 24004
rect 15916 23969 15956 24592
rect 16012 24583 16052 24592
rect 16108 24632 16148 24835
rect 16108 24583 16148 24592
rect 16204 24548 16244 26944
rect 16300 26816 16340 26825
rect 16300 25145 16340 26776
rect 16396 26657 16436 30640
rect 16492 30269 16532 32143
rect 16491 30260 16533 30269
rect 16491 30220 16492 30260
rect 16532 30220 16533 30260
rect 16491 30211 16533 30220
rect 16588 29933 16628 32992
rect 17068 32948 17108 32992
rect 17164 32948 17204 32957
rect 17068 32908 17164 32948
rect 17164 32899 17204 32908
rect 17260 32948 17300 33235
rect 17355 33032 17397 33041
rect 17355 32992 17356 33032
rect 17396 32992 17397 33032
rect 17355 32983 17397 32992
rect 17260 32899 17300 32908
rect 16684 32864 16724 32873
rect 16684 32276 16724 32824
rect 16780 32864 16820 32873
rect 16780 32705 16820 32824
rect 17356 32780 17396 32983
rect 17164 32740 17396 32780
rect 16779 32696 16821 32705
rect 16779 32656 16780 32696
rect 16820 32656 16821 32696
rect 16779 32647 16821 32656
rect 16780 32453 16820 32647
rect 16779 32444 16821 32453
rect 16779 32404 16780 32444
rect 16820 32404 16821 32444
rect 16779 32395 16821 32404
rect 17164 32360 17204 32740
rect 17164 32311 17204 32320
rect 16972 32276 17012 32285
rect 16684 32236 16916 32276
rect 16780 32178 16820 32187
rect 16780 31604 16820 32138
rect 16684 31564 16820 31604
rect 16684 31109 16724 31564
rect 16876 31520 16916 32236
rect 17012 32236 17108 32276
rect 16972 32227 17012 32236
rect 16972 31520 17012 31529
rect 16876 31480 16972 31520
rect 16972 31471 17012 31480
rect 16780 31352 16820 31361
rect 16820 31312 16916 31352
rect 16780 31303 16820 31312
rect 16779 31184 16821 31193
rect 16779 31144 16780 31184
rect 16820 31144 16821 31184
rect 16779 31135 16821 31144
rect 16683 31100 16725 31109
rect 16683 31060 16684 31100
rect 16724 31060 16725 31100
rect 16683 31051 16725 31060
rect 16780 30596 16820 31135
rect 16876 30689 16916 31312
rect 16875 30680 16917 30689
rect 16875 30640 16876 30680
rect 16916 30640 16917 30680
rect 16875 30631 16917 30640
rect 16780 30547 16820 30556
rect 16972 30428 17012 30437
rect 16684 30388 16972 30428
rect 17068 30428 17108 32236
rect 17355 32192 17397 32201
rect 17355 32152 17356 32192
rect 17396 32152 17397 32192
rect 17355 32143 17397 32152
rect 17356 31697 17396 32143
rect 17355 31688 17397 31697
rect 17355 31648 17356 31688
rect 17396 31648 17397 31688
rect 17355 31639 17397 31648
rect 17452 31520 17492 35260
rect 17548 35251 17588 35260
rect 17644 35888 17684 35897
rect 17547 34544 17589 34553
rect 17547 34504 17548 34544
rect 17588 34504 17589 34544
rect 17644 34544 17684 35848
rect 17739 35888 17781 35897
rect 17739 35848 17740 35888
rect 17780 35848 17781 35888
rect 17739 35839 17781 35848
rect 17740 35754 17780 35839
rect 18124 35838 18164 35923
rect 18220 35888 18260 36763
rect 17739 35384 17781 35393
rect 17739 35344 17740 35384
rect 17780 35344 17781 35384
rect 17739 35335 17781 35344
rect 17740 35216 17780 35335
rect 17740 35167 17780 35176
rect 17644 34504 17780 34544
rect 17547 34495 17589 34504
rect 17548 34376 17588 34495
rect 17548 34327 17588 34336
rect 17644 34376 17684 34385
rect 17644 34217 17684 34336
rect 17643 34208 17685 34217
rect 17643 34168 17644 34208
rect 17684 34168 17685 34208
rect 17643 34159 17685 34168
rect 17547 34124 17589 34133
rect 17547 34084 17548 34124
rect 17588 34084 17589 34124
rect 17547 34075 17589 34084
rect 17548 32705 17588 34075
rect 17740 33881 17780 34504
rect 18028 34376 18068 34385
rect 18028 34133 18068 34336
rect 18123 34376 18165 34385
rect 18123 34336 18124 34376
rect 18164 34336 18165 34376
rect 18123 34327 18165 34336
rect 18027 34124 18069 34133
rect 18027 34084 18028 34124
rect 18068 34084 18069 34124
rect 18027 34075 18069 34084
rect 17739 33872 17781 33881
rect 17739 33832 17740 33872
rect 17780 33832 17781 33872
rect 17739 33823 17781 33832
rect 17740 32864 17780 32873
rect 17644 32824 17740 32864
rect 17547 32696 17589 32705
rect 17547 32656 17548 32696
rect 17588 32656 17589 32696
rect 17547 32647 17589 32656
rect 17356 31480 17492 31520
rect 17163 31436 17205 31445
rect 17163 31396 17164 31436
rect 17204 31396 17205 31436
rect 17163 31387 17205 31396
rect 17164 30596 17204 31387
rect 17260 31352 17300 31361
rect 17260 30857 17300 31312
rect 17356 31352 17396 31480
rect 17356 31025 17396 31312
rect 17451 31352 17493 31361
rect 17451 31312 17452 31352
rect 17492 31312 17493 31352
rect 17451 31303 17493 31312
rect 17355 31016 17397 31025
rect 17355 30976 17356 31016
rect 17396 30976 17397 31016
rect 17355 30967 17397 30976
rect 17259 30848 17301 30857
rect 17259 30808 17260 30848
rect 17300 30808 17301 30848
rect 17259 30799 17301 30808
rect 17356 30848 17396 30857
rect 17452 30848 17492 31303
rect 17396 30808 17492 30848
rect 17356 30799 17396 30808
rect 17164 30547 17204 30556
rect 17068 30388 17300 30428
rect 16587 29924 16629 29933
rect 16587 29884 16588 29924
rect 16628 29884 16629 29924
rect 16587 29875 16629 29884
rect 16587 29672 16629 29681
rect 16587 29632 16588 29672
rect 16628 29632 16629 29672
rect 16587 29623 16629 29632
rect 16491 29168 16533 29177
rect 16491 29128 16492 29168
rect 16532 29128 16533 29168
rect 16491 29119 16533 29128
rect 16588 29168 16628 29623
rect 16588 29119 16628 29128
rect 16492 29034 16532 29119
rect 16587 28244 16629 28253
rect 16587 28204 16588 28244
rect 16628 28204 16629 28244
rect 16587 28195 16629 28204
rect 16588 27824 16628 28195
rect 16684 28001 16724 30388
rect 16972 30379 17012 30388
rect 17067 30260 17109 30269
rect 17067 30220 17068 30260
rect 17108 30220 17109 30260
rect 17067 30211 17109 30220
rect 16780 29924 16820 29933
rect 16820 29884 16916 29924
rect 16780 29875 16820 29884
rect 16779 29756 16821 29765
rect 16779 29716 16780 29756
rect 16820 29716 16821 29756
rect 16779 29707 16821 29716
rect 16683 27992 16725 28001
rect 16683 27952 16684 27992
rect 16724 27952 16725 27992
rect 16683 27943 16725 27952
rect 16588 27775 16628 27784
rect 16683 27824 16725 27833
rect 16683 27784 16684 27824
rect 16724 27784 16725 27824
rect 16780 27824 16820 29707
rect 16876 28169 16916 29884
rect 17068 29756 17108 30211
rect 17163 30092 17205 30101
rect 17163 30052 17164 30092
rect 17204 30052 17205 30092
rect 17163 30043 17205 30052
rect 17164 29924 17204 30043
rect 17164 29875 17204 29884
rect 17068 29716 17204 29756
rect 16972 29672 17012 29681
rect 17012 29632 17108 29672
rect 16972 29623 17012 29632
rect 17068 29261 17108 29632
rect 17067 29252 17109 29261
rect 17067 29212 17068 29252
rect 17108 29212 17109 29252
rect 17067 29203 17109 29212
rect 16972 29093 17012 29178
rect 16971 29084 17013 29093
rect 16971 29044 16972 29084
rect 17012 29044 17013 29084
rect 16971 29035 17013 29044
rect 17068 29084 17108 29095
rect 17068 28925 17108 29044
rect 17067 28916 17109 28925
rect 17067 28876 17068 28916
rect 17108 28876 17109 28916
rect 17067 28867 17109 28876
rect 16875 28160 16917 28169
rect 16875 28120 16876 28160
rect 16916 28120 16917 28160
rect 16875 28111 16917 28120
rect 16780 27784 16916 27824
rect 16683 27775 16725 27784
rect 16684 27656 16724 27775
rect 16492 27645 16532 27654
rect 16684 27607 16724 27616
rect 16780 27656 16820 27665
rect 16395 26648 16437 26657
rect 16395 26608 16396 26648
rect 16436 26608 16437 26648
rect 16395 26599 16437 26608
rect 16492 26573 16532 27605
rect 16587 27236 16629 27245
rect 16587 27196 16588 27236
rect 16628 27196 16629 27236
rect 16587 27187 16629 27196
rect 16588 26816 16628 27187
rect 16588 26767 16628 26776
rect 16683 26816 16725 26825
rect 16683 26776 16684 26816
rect 16724 26776 16725 26816
rect 16683 26767 16725 26776
rect 16684 26682 16724 26767
rect 16491 26564 16533 26573
rect 16491 26524 16492 26564
rect 16532 26524 16533 26564
rect 16491 26515 16533 26524
rect 16683 26564 16725 26573
rect 16683 26524 16684 26564
rect 16724 26524 16725 26564
rect 16683 26515 16725 26524
rect 16395 25808 16437 25817
rect 16395 25768 16396 25808
rect 16436 25768 16437 25808
rect 16395 25759 16437 25768
rect 16299 25136 16341 25145
rect 16299 25096 16300 25136
rect 16340 25096 16341 25136
rect 16299 25087 16341 25096
rect 16204 24508 16340 24548
rect 16011 24380 16053 24389
rect 16011 24340 16012 24380
rect 16052 24340 16053 24380
rect 16011 24331 16053 24340
rect 15915 23960 15957 23969
rect 15915 23920 15916 23960
rect 15956 23920 15957 23960
rect 15915 23911 15957 23920
rect 15916 23834 15956 23843
rect 15916 23792 15956 23794
rect 15724 23752 15956 23792
rect 15724 22541 15764 23752
rect 16012 23540 16052 24331
rect 16107 24044 16149 24053
rect 16107 24004 16108 24044
rect 16148 24004 16149 24044
rect 16107 23995 16149 24004
rect 15916 23500 16052 23540
rect 15916 23120 15956 23500
rect 15916 23071 15956 23080
rect 16012 23120 16052 23129
rect 16108 23120 16148 23995
rect 16052 23080 16148 23120
rect 16203 23120 16245 23129
rect 16203 23080 16204 23120
rect 16244 23080 16245 23120
rect 16012 23071 16052 23080
rect 16203 23071 16245 23080
rect 16204 22986 16244 23071
rect 16204 22868 16244 22877
rect 15820 22828 16204 22868
rect 15723 22532 15765 22541
rect 15723 22492 15724 22532
rect 15764 22492 15765 22532
rect 15723 22483 15765 22492
rect 15723 22364 15765 22373
rect 15723 22324 15724 22364
rect 15764 22324 15765 22364
rect 15723 22315 15765 22324
rect 15627 22112 15669 22121
rect 15627 22072 15628 22112
rect 15668 22072 15669 22112
rect 15627 22063 15669 22072
rect 15532 21904 15668 21944
rect 15244 21820 15572 21860
rect 15339 21692 15381 21701
rect 15339 21652 15340 21692
rect 15380 21652 15381 21692
rect 15339 21643 15381 21652
rect 15243 21608 15285 21617
rect 15243 21568 15244 21608
rect 15284 21568 15285 21608
rect 15243 21559 15285 21568
rect 15340 21608 15380 21643
rect 15244 21474 15284 21559
rect 15340 21557 15380 21568
rect 15532 21608 15572 21820
rect 15532 21559 15572 21568
rect 15435 21524 15477 21533
rect 15435 21484 15436 21524
rect 15476 21484 15477 21524
rect 15435 21475 15477 21484
rect 15339 20936 15381 20945
rect 15339 20896 15340 20936
rect 15380 20896 15381 20936
rect 15339 20887 15381 20896
rect 15340 20768 15380 20887
rect 15148 20728 15284 20768
rect 15147 20600 15189 20609
rect 15147 20560 15148 20600
rect 15188 20560 15189 20600
rect 15147 20551 15189 20560
rect 15148 20466 15188 20551
rect 14996 20224 15092 20264
rect 14956 20215 14996 20224
rect 15244 20180 15284 20728
rect 15340 20525 15380 20728
rect 15436 20768 15476 21475
rect 15628 21356 15668 21904
rect 15724 21533 15764 22315
rect 15723 21524 15765 21533
rect 15723 21484 15724 21524
rect 15764 21484 15765 21524
rect 15820 21524 15860 22828
rect 16204 22819 16244 22828
rect 16011 22700 16053 22709
rect 16011 22660 16012 22700
rect 16052 22660 16053 22700
rect 16011 22651 16053 22660
rect 16012 22289 16052 22651
rect 16107 22364 16149 22373
rect 16107 22324 16108 22364
rect 16148 22324 16149 22364
rect 16107 22315 16149 22324
rect 16007 22280 16052 22289
rect 16047 22240 16052 22280
rect 16108 22280 16148 22315
rect 16007 22231 16047 22240
rect 16108 22229 16148 22240
rect 16204 22280 16244 22289
rect 16011 22112 16053 22121
rect 16011 22072 16012 22112
rect 16052 22072 16053 22112
rect 16011 22063 16053 22072
rect 16108 22112 16148 22121
rect 15820 21484 15956 21524
rect 15723 21475 15765 21484
rect 15628 21316 15764 21356
rect 15627 21188 15669 21197
rect 15627 21148 15628 21188
rect 15668 21148 15669 21188
rect 15627 21139 15669 21148
rect 15436 20719 15476 20728
rect 15628 20768 15668 21139
rect 15628 20719 15668 20728
rect 15339 20516 15381 20525
rect 15339 20476 15340 20516
rect 15380 20476 15381 20516
rect 15339 20467 15381 20476
rect 15627 20516 15669 20525
rect 15627 20476 15628 20516
rect 15668 20476 15669 20516
rect 15627 20467 15669 20476
rect 15244 20140 15572 20180
rect 14764 20096 14804 20124
rect 14668 20056 14764 20096
rect 14668 18929 14708 20056
rect 14764 20047 14804 20056
rect 14859 19508 14901 19517
rect 14859 19468 14860 19508
rect 14900 19468 14901 19508
rect 14859 19459 14901 19468
rect 14763 19340 14805 19349
rect 14763 19300 14764 19340
rect 14804 19300 14805 19340
rect 14763 19291 14805 19300
rect 14667 18920 14709 18929
rect 14667 18880 14668 18920
rect 14708 18880 14709 18920
rect 14667 18871 14709 18880
rect 14284 18796 14516 18836
rect 14284 17744 14324 18796
rect 14667 18752 14709 18761
rect 14667 18712 14668 18752
rect 14708 18712 14709 18752
rect 14667 18703 14709 18712
rect 14668 18618 14708 18703
rect 14476 18584 14516 18593
rect 14516 18544 14612 18584
rect 14476 18535 14516 18544
rect 14572 18425 14612 18544
rect 14764 18500 14804 19291
rect 14668 18460 14804 18500
rect 14571 18416 14613 18425
rect 14571 18376 14572 18416
rect 14612 18376 14613 18416
rect 14571 18367 14613 18376
rect 14475 18332 14517 18341
rect 14475 18292 14476 18332
rect 14516 18292 14517 18332
rect 14475 18283 14517 18292
rect 14379 18248 14421 18257
rect 14379 18208 14380 18248
rect 14420 18208 14421 18248
rect 14379 18199 14421 18208
rect 14284 17695 14324 17704
rect 14283 14888 14325 14897
rect 14283 14848 14284 14888
rect 14324 14848 14325 14888
rect 14283 14839 14325 14848
rect 14284 12713 14324 14839
rect 14380 14720 14420 18199
rect 14476 16904 14516 18283
rect 14668 17249 14708 18460
rect 14860 18416 14900 19459
rect 15339 19424 15381 19433
rect 15339 19384 15340 19424
rect 15380 19384 15381 19424
rect 15339 19375 15381 19384
rect 14955 18752 14997 18761
rect 14955 18712 14956 18752
rect 14996 18712 14997 18752
rect 14955 18703 14997 18712
rect 14956 18584 14996 18703
rect 15051 18668 15093 18677
rect 15051 18628 15052 18668
rect 15092 18628 15093 18668
rect 15051 18619 15093 18628
rect 14956 18535 14996 18544
rect 15052 18584 15092 18619
rect 15052 18533 15092 18544
rect 15051 18416 15093 18425
rect 14860 18376 14996 18416
rect 14667 17240 14709 17249
rect 14667 17200 14668 17240
rect 14708 17200 14709 17240
rect 14667 17191 14709 17200
rect 14764 17165 14804 17250
rect 14763 17156 14805 17165
rect 14763 17116 14764 17156
rect 14804 17116 14805 17156
rect 14763 17107 14805 17116
rect 14620 17030 14660 17039
rect 14620 16988 14660 16990
rect 14620 16948 14900 16988
rect 14476 16864 14612 16904
rect 14476 14720 14516 14729
rect 14380 14680 14476 14720
rect 14476 14561 14516 14680
rect 14475 14552 14517 14561
rect 14475 14512 14476 14552
rect 14516 14512 14517 14552
rect 14475 14503 14517 14512
rect 14476 14048 14516 14503
rect 14476 13999 14516 14008
rect 14379 13208 14421 13217
rect 14379 13168 14380 13208
rect 14420 13168 14421 13208
rect 14379 13159 14421 13168
rect 14476 13213 14516 13222
rect 14283 12704 14325 12713
rect 14283 12664 14284 12704
rect 14324 12664 14325 12704
rect 14283 12655 14325 12664
rect 14284 12536 14324 12547
rect 14284 12461 14324 12496
rect 14283 12452 14325 12461
rect 14283 12412 14284 12452
rect 14324 12412 14325 12452
rect 14283 12403 14325 12412
rect 14284 11705 14324 12403
rect 14283 11696 14325 11705
rect 14283 11656 14284 11696
rect 14324 11656 14325 11696
rect 14283 11647 14325 11656
rect 14380 11444 14420 13159
rect 14476 12704 14516 13173
rect 14572 12872 14612 16864
rect 14763 16736 14805 16745
rect 14763 16696 14764 16736
rect 14804 16696 14805 16736
rect 14763 16687 14805 16696
rect 14667 16400 14709 16409
rect 14667 16360 14668 16400
rect 14708 16360 14709 16400
rect 14667 16351 14709 16360
rect 14668 16232 14708 16351
rect 14668 16183 14708 16192
rect 14667 16064 14709 16073
rect 14667 16024 14668 16064
rect 14708 16024 14709 16064
rect 14667 16015 14709 16024
rect 14668 13721 14708 16015
rect 14667 13712 14709 13721
rect 14667 13672 14668 13712
rect 14708 13672 14709 13712
rect 14667 13663 14709 13672
rect 14667 13124 14709 13133
rect 14667 13084 14668 13124
rect 14708 13084 14709 13124
rect 14667 13075 14709 13084
rect 14668 12990 14708 13075
rect 14572 12832 14708 12872
rect 14476 12655 14516 12664
rect 14571 11612 14613 11621
rect 14571 11572 14572 11612
rect 14612 11572 14613 11612
rect 14571 11563 14613 11572
rect 14375 11404 14420 11444
rect 14188 11320 14324 11360
rect 13803 11276 13845 11285
rect 13803 11236 13804 11276
rect 13844 11236 13845 11276
rect 13803 11227 13845 11236
rect 14284 11234 14324 11320
rect 13804 11024 13844 11227
rect 13995 11192 14037 11201
rect 13995 11152 13996 11192
rect 14036 11152 14037 11192
rect 13995 11143 14037 11152
rect 14188 11194 14324 11234
rect 14375 11234 14415 11404
rect 14375 11194 14420 11234
rect 13899 11108 13941 11117
rect 13899 11068 13900 11108
rect 13940 11068 13941 11108
rect 13899 11059 13941 11068
rect 13804 10975 13844 10984
rect 13900 10940 13940 11059
rect 13900 10865 13940 10900
rect 13899 10856 13941 10865
rect 13899 10816 13900 10856
rect 13940 10816 13941 10856
rect 13899 10807 13941 10816
rect 13803 9764 13845 9773
rect 13803 9724 13804 9764
rect 13844 9724 13845 9764
rect 13803 9715 13845 9724
rect 13516 9640 13748 9680
rect 13419 8168 13461 8177
rect 13419 8128 13420 8168
rect 13460 8128 13461 8168
rect 13419 8119 13461 8128
rect 13419 8000 13461 8009
rect 13419 7960 13420 8000
rect 13460 7960 13461 8000
rect 13419 7951 13461 7960
rect 13420 7866 13460 7951
rect 13132 7110 13172 7195
rect 13228 7085 13268 7204
rect 13516 7169 13556 9640
rect 13612 9512 13652 9523
rect 13612 9437 13652 9472
rect 13707 9512 13749 9521
rect 13707 9472 13708 9512
rect 13748 9472 13749 9512
rect 13707 9463 13749 9472
rect 13804 9512 13844 9715
rect 13804 9463 13844 9472
rect 13900 9512 13940 9521
rect 13611 9428 13653 9437
rect 13611 9388 13612 9428
rect 13652 9388 13653 9428
rect 13611 9379 13653 9388
rect 13708 9378 13748 9463
rect 13611 8588 13653 8597
rect 13611 8548 13612 8588
rect 13652 8548 13653 8588
rect 13611 8539 13653 8548
rect 13612 8009 13652 8539
rect 13900 8177 13940 9472
rect 13996 8597 14036 11143
rect 14091 11108 14133 11117
rect 14091 11068 14092 11108
rect 14132 11068 14133 11108
rect 14091 11059 14133 11068
rect 13995 8588 14037 8597
rect 13995 8548 13996 8588
rect 14036 8548 14037 8588
rect 13995 8539 14037 8548
rect 13899 8168 13941 8177
rect 13899 8128 13900 8168
rect 13940 8128 13941 8168
rect 13899 8119 13941 8128
rect 13611 8000 13653 8009
rect 13611 7960 13612 8000
rect 13652 7960 13653 8000
rect 13611 7951 13653 7960
rect 13707 7328 13749 7337
rect 13707 7288 13708 7328
rect 13748 7288 13749 7328
rect 13707 7279 13749 7288
rect 13515 7160 13557 7169
rect 13515 7120 13516 7160
rect 13556 7120 13557 7160
rect 13515 7111 13557 7120
rect 13708 7160 13748 7279
rect 13708 7111 13748 7120
rect 13227 7076 13269 7085
rect 13227 7036 13228 7076
rect 13268 7036 13269 7076
rect 13227 7027 13269 7036
rect 13323 6992 13365 7001
rect 13323 6952 13324 6992
rect 13364 6952 13365 6992
rect 13323 6943 13365 6952
rect 13035 3884 13077 3893
rect 13035 3844 13036 3884
rect 13076 3844 13077 3884
rect 13035 3835 13077 3844
rect 12939 3128 12981 3137
rect 12939 3088 12940 3128
rect 12980 3088 12981 3128
rect 12939 3079 12981 3088
rect 12748 1819 12788 1828
rect 13324 1868 13364 6943
rect 14092 6917 14132 11059
rect 14188 7328 14228 11194
rect 14380 11024 14420 11194
rect 14420 10984 14516 11024
rect 14380 10975 14420 10984
rect 14379 10016 14421 10025
rect 14379 9976 14380 10016
rect 14420 9976 14421 10016
rect 14379 9967 14421 9976
rect 14284 9521 14324 9606
rect 14283 9512 14325 9521
rect 14283 9472 14284 9512
rect 14324 9472 14325 9512
rect 14283 9463 14325 9472
rect 14380 9512 14420 9967
rect 14476 9680 14516 10984
rect 14572 10184 14612 11563
rect 14668 10949 14708 12832
rect 14764 11360 14804 16687
rect 14860 16484 14900 16948
rect 14860 16435 14900 16444
rect 14956 16073 14996 18376
rect 15051 18376 15052 18416
rect 15092 18376 15093 18416
rect 15051 18367 15093 18376
rect 15052 16997 15092 18367
rect 15243 17744 15285 17753
rect 15243 17704 15244 17744
rect 15284 17704 15285 17744
rect 15340 17744 15380 19375
rect 15532 18584 15572 20140
rect 15532 18535 15572 18544
rect 15436 18500 15476 18509
rect 15436 18173 15476 18460
rect 15435 18164 15477 18173
rect 15435 18124 15436 18164
rect 15476 18124 15477 18164
rect 15435 18115 15477 18124
rect 15628 18005 15668 20467
rect 15627 17996 15669 18005
rect 15627 17956 15628 17996
rect 15668 17956 15669 17996
rect 15627 17947 15669 17956
rect 15532 17744 15572 17753
rect 15724 17744 15764 21316
rect 15820 20096 15860 20105
rect 15820 19508 15860 20056
rect 15916 19685 15956 21484
rect 16012 21449 16052 22063
rect 16011 21440 16053 21449
rect 16011 21400 16012 21440
rect 16052 21400 16053 21440
rect 16011 21391 16053 21400
rect 15915 19676 15957 19685
rect 15915 19636 15916 19676
rect 15956 19636 15957 19676
rect 15915 19627 15957 19636
rect 15820 19468 15956 19508
rect 15819 19256 15861 19265
rect 15819 19216 15820 19256
rect 15860 19216 15861 19256
rect 15819 19207 15861 19216
rect 15340 17704 15532 17744
rect 15243 17695 15285 17704
rect 15147 17072 15189 17081
rect 15147 17032 15148 17072
rect 15188 17032 15189 17072
rect 15147 17023 15189 17032
rect 15051 16988 15093 16997
rect 15051 16948 15052 16988
rect 15092 16948 15093 16988
rect 15051 16939 15093 16948
rect 15052 16409 15092 16939
rect 15148 16938 15188 17023
rect 15051 16400 15093 16409
rect 15051 16360 15052 16400
rect 15092 16360 15093 16400
rect 15051 16351 15093 16360
rect 15244 16316 15284 17695
rect 15532 16745 15572 17704
rect 15628 17704 15764 17744
rect 15531 16736 15573 16745
rect 15531 16696 15532 16736
rect 15572 16696 15573 16736
rect 15531 16687 15573 16696
rect 15339 16568 15381 16577
rect 15339 16528 15340 16568
rect 15380 16528 15381 16568
rect 15339 16519 15381 16528
rect 15244 16267 15284 16276
rect 14955 16064 14997 16073
rect 14955 16024 14956 16064
rect 14996 16024 14997 16064
rect 14955 16015 14997 16024
rect 14955 15560 14997 15569
rect 14955 15520 14956 15560
rect 14996 15520 14997 15560
rect 15340 15560 15380 16519
rect 15435 16400 15477 16409
rect 15628 16400 15668 17704
rect 15435 16360 15436 16400
rect 15476 16360 15477 16400
rect 15435 16351 15477 16360
rect 15532 16360 15668 16400
rect 15724 17576 15764 17585
rect 15436 16266 15476 16351
rect 15532 15728 15572 16360
rect 15627 16232 15669 16241
rect 15627 16192 15628 16232
rect 15668 16192 15669 16232
rect 15627 16183 15669 16192
rect 15628 16098 15668 16183
rect 15532 15688 15668 15728
rect 15532 15560 15572 15569
rect 15340 15520 15532 15560
rect 14955 15511 14997 15520
rect 15532 15511 15572 15520
rect 14956 15426 14996 15511
rect 15148 15308 15188 15317
rect 14860 15268 15148 15308
rect 14860 14636 14900 15268
rect 15148 15259 15188 15268
rect 15004 14729 15044 14738
rect 15532 14720 15572 14729
rect 15044 14689 15284 14720
rect 15004 14680 15284 14689
rect 15244 14636 15284 14680
rect 15436 14680 15532 14720
rect 15340 14636 15380 14645
rect 14860 14596 14996 14636
rect 15244 14596 15340 14636
rect 14956 14043 14996 14596
rect 15340 14587 15380 14596
rect 15147 14552 15189 14561
rect 15147 14512 15148 14552
rect 15188 14512 15189 14552
rect 15147 14503 15189 14512
rect 15148 14418 15188 14503
rect 14956 13994 14996 14003
rect 15148 14132 15188 14141
rect 15148 12713 15188 14092
rect 15436 14057 15476 14680
rect 15532 14671 15572 14680
rect 15531 14132 15573 14141
rect 15531 14092 15532 14132
rect 15572 14092 15573 14132
rect 15531 14083 15573 14092
rect 15435 14048 15477 14057
rect 15435 14008 15436 14048
rect 15476 14008 15477 14048
rect 15435 13999 15477 14008
rect 15243 13208 15285 13217
rect 15243 13168 15244 13208
rect 15284 13168 15285 13208
rect 15243 13159 15285 13168
rect 15532 13208 15572 14083
rect 15244 13074 15284 13159
rect 15532 13133 15572 13168
rect 15628 13208 15668 15688
rect 15724 14048 15764 17536
rect 15820 17081 15860 19207
rect 15916 18593 15956 19468
rect 15915 18584 15957 18593
rect 15915 18544 15916 18584
rect 15956 18544 15957 18584
rect 15915 18535 15957 18544
rect 16012 18584 16052 18593
rect 16012 18341 16052 18544
rect 16011 18332 16053 18341
rect 16011 18292 16012 18332
rect 16052 18292 16053 18332
rect 16011 18283 16053 18292
rect 15915 17996 15957 18005
rect 15915 17956 15916 17996
rect 15956 17956 15957 17996
rect 15915 17947 15957 17956
rect 15819 17072 15861 17081
rect 15819 17032 15820 17072
rect 15860 17032 15861 17072
rect 15819 17023 15861 17032
rect 15819 16736 15861 16745
rect 15819 16696 15820 16736
rect 15860 16696 15861 16736
rect 15819 16687 15861 16696
rect 15820 15569 15860 16687
rect 15819 15560 15861 15569
rect 15819 15520 15820 15560
rect 15860 15520 15861 15560
rect 15819 15511 15861 15520
rect 15916 14645 15956 17947
rect 16011 17912 16053 17921
rect 16011 17872 16012 17912
rect 16052 17872 16053 17912
rect 16011 17863 16053 17872
rect 15915 14636 15957 14645
rect 15915 14596 15916 14636
rect 15956 14596 15957 14636
rect 15915 14587 15957 14596
rect 15916 14309 15956 14587
rect 16012 14393 16052 17863
rect 16108 15485 16148 22072
rect 16204 20609 16244 22240
rect 16203 20600 16245 20609
rect 16203 20560 16204 20600
rect 16244 20560 16245 20600
rect 16203 20551 16245 20560
rect 16203 20348 16245 20357
rect 16203 20308 16204 20348
rect 16244 20308 16245 20348
rect 16203 20299 16245 20308
rect 16204 19265 16244 20299
rect 16203 19256 16245 19265
rect 16203 19216 16204 19256
rect 16244 19216 16245 19256
rect 16203 19207 16245 19216
rect 16203 18668 16245 18677
rect 16203 18628 16204 18668
rect 16244 18628 16245 18668
rect 16203 18619 16245 18628
rect 16204 17828 16244 18619
rect 16204 17779 16244 17788
rect 16107 15476 16149 15485
rect 16107 15436 16108 15476
rect 16148 15436 16149 15476
rect 16107 15427 16149 15436
rect 16011 14384 16053 14393
rect 16011 14344 16012 14384
rect 16052 14344 16053 14384
rect 16011 14335 16053 14344
rect 15915 14300 15957 14309
rect 15915 14260 15916 14300
rect 15956 14260 15957 14300
rect 15915 14251 15957 14260
rect 16300 14141 16340 24508
rect 16396 23885 16436 25759
rect 16491 24632 16533 24641
rect 16491 24592 16492 24632
rect 16532 24592 16533 24632
rect 16491 24583 16533 24592
rect 16492 24498 16532 24583
rect 16588 24548 16628 24557
rect 16588 24221 16628 24508
rect 16587 24212 16629 24221
rect 16587 24172 16588 24212
rect 16628 24172 16629 24212
rect 16587 24163 16629 24172
rect 16587 23960 16629 23969
rect 16587 23920 16588 23960
rect 16628 23920 16629 23960
rect 16587 23911 16629 23920
rect 16395 23876 16437 23885
rect 16395 23836 16396 23876
rect 16436 23836 16437 23876
rect 16395 23827 16437 23836
rect 16396 23456 16436 23827
rect 16396 23416 16532 23456
rect 16395 23288 16437 23297
rect 16395 23248 16396 23288
rect 16436 23248 16437 23288
rect 16395 23239 16437 23248
rect 16396 22709 16436 23239
rect 16492 23045 16532 23416
rect 16588 23120 16628 23911
rect 16588 23071 16628 23080
rect 16491 23036 16533 23045
rect 16491 22996 16492 23036
rect 16532 22996 16533 23036
rect 16491 22987 16533 22996
rect 16684 22952 16724 26515
rect 16780 25220 16820 27616
rect 16876 26825 16916 27784
rect 17067 27572 17109 27581
rect 17067 27532 17068 27572
rect 17108 27532 17109 27572
rect 17067 27523 17109 27532
rect 17068 27438 17108 27523
rect 16972 26984 17012 26993
rect 16875 26816 16917 26825
rect 16875 26776 16876 26816
rect 16916 26776 16917 26816
rect 16875 26767 16917 26776
rect 16875 26648 16917 26657
rect 16875 26608 16876 26648
rect 16916 26608 16917 26648
rect 16875 26599 16917 26608
rect 16876 26312 16916 26599
rect 16972 26489 17012 26944
rect 16971 26480 17013 26489
rect 16971 26440 16972 26480
rect 17012 26440 17013 26480
rect 16971 26431 17013 26440
rect 17068 26321 17108 26406
rect 17067 26312 17109 26321
rect 16876 26272 17012 26312
rect 16876 26144 16916 26153
rect 16876 26069 16916 26104
rect 16875 26060 16917 26069
rect 16875 26020 16876 26060
rect 16916 26020 16917 26060
rect 16875 26011 16917 26020
rect 16876 25733 16916 26011
rect 16875 25724 16917 25733
rect 16875 25684 16876 25724
rect 16916 25684 16917 25724
rect 16875 25675 16917 25684
rect 16780 25180 16916 25220
rect 16779 25052 16821 25061
rect 16779 25012 16780 25052
rect 16820 25012 16821 25052
rect 16779 25003 16821 25012
rect 16588 22912 16724 22952
rect 16395 22700 16437 22709
rect 16395 22660 16396 22700
rect 16436 22660 16437 22700
rect 16395 22651 16437 22660
rect 16396 22280 16436 22289
rect 16396 21617 16436 22240
rect 16492 22280 16532 22289
rect 16492 21701 16532 22240
rect 16491 21692 16533 21701
rect 16491 21652 16492 21692
rect 16532 21652 16533 21692
rect 16491 21643 16533 21652
rect 16395 21608 16437 21617
rect 16395 21568 16396 21608
rect 16436 21568 16437 21608
rect 16395 21559 16437 21568
rect 16492 18570 16532 18579
rect 16396 17576 16436 17585
rect 16396 17249 16436 17536
rect 16395 17240 16437 17249
rect 16395 17200 16396 17240
rect 16436 17200 16437 17240
rect 16492 17240 16532 18530
rect 16588 17996 16628 22912
rect 16683 22364 16725 22373
rect 16683 22324 16684 22364
rect 16724 22324 16725 22364
rect 16683 22315 16725 22324
rect 16684 22280 16724 22315
rect 16684 22229 16724 22240
rect 16780 22112 16820 25003
rect 16876 23297 16916 25180
rect 16875 23288 16917 23297
rect 16875 23248 16876 23288
rect 16916 23248 16917 23288
rect 16875 23239 16917 23248
rect 16876 23120 16916 23131
rect 16876 23045 16916 23080
rect 16972 23120 17012 26272
rect 17067 26272 17068 26312
rect 17108 26272 17109 26312
rect 17067 26263 17109 26272
rect 17067 26144 17109 26153
rect 17067 26104 17068 26144
rect 17108 26104 17109 26144
rect 17067 26095 17109 26104
rect 17068 24632 17108 26095
rect 17068 24583 17108 24592
rect 17164 23960 17204 29716
rect 17260 28421 17300 30388
rect 17547 30092 17589 30101
rect 17644 30092 17684 32824
rect 17740 32815 17780 32824
rect 18027 32864 18069 32873
rect 18027 32824 18028 32864
rect 18068 32824 18069 32864
rect 18027 32815 18069 32824
rect 17739 31436 17781 31445
rect 17739 31396 17740 31436
rect 17780 31396 17781 31436
rect 17739 31387 17781 31396
rect 17740 30269 17780 31387
rect 17836 31352 17876 31363
rect 17836 31277 17876 31312
rect 17835 31268 17877 31277
rect 17835 31228 17836 31268
rect 17876 31228 17877 31268
rect 17835 31219 17877 31228
rect 17836 30689 17876 30774
rect 17835 30680 17877 30689
rect 17835 30640 17836 30680
rect 17876 30640 17877 30680
rect 17835 30631 17877 30640
rect 17931 30512 17973 30521
rect 17931 30472 17932 30512
rect 17972 30472 17973 30512
rect 17931 30463 17973 30472
rect 17835 30428 17877 30437
rect 17835 30388 17836 30428
rect 17876 30388 17877 30428
rect 17835 30379 17877 30388
rect 17739 30260 17781 30269
rect 17739 30220 17740 30260
rect 17780 30220 17781 30260
rect 17739 30211 17781 30220
rect 17547 30052 17548 30092
rect 17588 30052 17684 30092
rect 17547 30043 17589 30052
rect 17355 29672 17397 29681
rect 17355 29632 17356 29672
rect 17396 29632 17397 29672
rect 17355 29623 17397 29632
rect 17356 29538 17396 29623
rect 17548 29429 17588 30043
rect 17644 29840 17684 29849
rect 17547 29420 17589 29429
rect 17547 29380 17548 29420
rect 17588 29380 17589 29420
rect 17547 29371 17589 29380
rect 17548 29168 17588 29371
rect 17548 29119 17588 29128
rect 17644 29000 17684 29800
rect 17739 29840 17781 29849
rect 17739 29800 17740 29840
rect 17780 29800 17781 29840
rect 17739 29791 17781 29800
rect 17740 29706 17780 29791
rect 17836 29093 17876 30379
rect 17932 29177 17972 30463
rect 18028 29345 18068 32815
rect 18124 32528 18164 34327
rect 18220 33797 18260 35848
rect 18604 35888 18644 37855
rect 18700 37745 18740 37948
rect 18796 37939 18836 37948
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 18699 37736 18741 37745
rect 18699 37696 18700 37736
rect 18740 37696 18741 37736
rect 18699 37687 18741 37696
rect 19276 37652 19316 37948
rect 19084 37612 19316 37652
rect 19084 37568 19124 37612
rect 19084 36896 19124 37528
rect 19275 37484 19317 37493
rect 19275 37444 19276 37484
rect 19316 37444 19317 37484
rect 19275 37435 19317 37444
rect 19276 37350 19316 37435
rect 19372 37157 19412 39628
rect 19467 39500 19509 39509
rect 19467 39460 19468 39500
rect 19508 39460 19509 39500
rect 19467 39451 19509 39460
rect 19468 39366 19508 39451
rect 19467 38744 19509 38753
rect 19467 38704 19468 38744
rect 19508 38704 19509 38744
rect 19467 38695 19509 38704
rect 19468 38610 19508 38695
rect 19467 38408 19509 38417
rect 19467 38368 19468 38408
rect 19508 38368 19509 38408
rect 19467 38359 19509 38368
rect 19468 38274 19508 38359
rect 19564 38156 19604 39787
rect 19659 39668 19701 39677
rect 19659 39628 19660 39668
rect 19700 39628 19701 39668
rect 19659 39619 19701 39628
rect 19660 39534 19700 39619
rect 19659 38996 19701 39005
rect 19659 38956 19660 38996
rect 19700 38956 19701 38996
rect 19659 38947 19701 38956
rect 19660 38862 19700 38947
rect 19660 38156 19700 38165
rect 19564 38116 19660 38156
rect 19660 38107 19700 38116
rect 19660 37484 19700 37493
rect 19660 37325 19700 37444
rect 19756 37400 19796 40888
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 20043 39920 20085 39929
rect 20043 39880 20044 39920
rect 20084 39880 20085 39920
rect 20043 39871 20085 39880
rect 19851 39752 19893 39761
rect 19851 39712 19852 39752
rect 19892 39712 19893 39752
rect 19851 39703 19893 39712
rect 19852 39584 19892 39703
rect 19852 39535 19892 39544
rect 19851 39080 19893 39089
rect 19851 39040 19852 39080
rect 19892 39040 19893 39080
rect 19851 39031 19893 39040
rect 19852 38946 19892 39031
rect 20044 38996 20084 39871
rect 20044 38947 20084 38956
rect 20236 38744 20276 38753
rect 20276 38704 21428 38744
rect 20236 38695 20276 38704
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 20043 38156 20085 38165
rect 20043 38116 20044 38156
rect 20084 38116 20085 38156
rect 20043 38107 20085 38116
rect 20044 38022 20084 38107
rect 20235 38072 20277 38081
rect 20235 38032 20236 38072
rect 20276 38032 20277 38072
rect 20235 38023 20277 38032
rect 19851 37988 19893 37997
rect 19851 37948 19852 37988
rect 19892 37948 19893 37988
rect 19851 37939 19893 37948
rect 19852 37854 19892 37939
rect 20236 37938 20276 38023
rect 20043 37484 20085 37493
rect 20043 37444 20044 37484
rect 20084 37444 20085 37484
rect 20043 37435 20085 37444
rect 19756 37360 19988 37400
rect 19659 37316 19701 37325
rect 19659 37276 19660 37316
rect 19700 37276 19701 37316
rect 19659 37267 19701 37276
rect 19468 37232 19508 37241
rect 19371 37148 19413 37157
rect 19371 37108 19372 37148
rect 19412 37108 19413 37148
rect 19371 37099 19413 37108
rect 19084 36847 19124 36856
rect 19468 36317 19508 37192
rect 19852 37232 19892 37241
rect 19852 37148 19892 37192
rect 19660 37108 19892 37148
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 19467 36308 19509 36317
rect 19467 36268 19468 36308
rect 19508 36268 19509 36308
rect 19467 36259 19509 36268
rect 18987 36140 19029 36149
rect 19660 36140 19700 37108
rect 19755 36980 19797 36989
rect 19755 36940 19756 36980
rect 19796 36940 19797 36980
rect 19755 36931 19797 36940
rect 18987 36100 18988 36140
rect 19028 36100 19029 36140
rect 18987 36091 19029 36100
rect 19276 36100 19700 36140
rect 19756 36140 19796 36931
rect 19948 36233 19988 37360
rect 20044 37350 20084 37435
rect 20235 37400 20277 37409
rect 20235 37360 20236 37400
rect 20276 37360 20277 37400
rect 20235 37351 20277 37360
rect 20236 37232 20276 37351
rect 20236 37183 20276 37192
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 20139 36728 20181 36737
rect 20139 36688 20140 36728
rect 20180 36688 20181 36728
rect 20139 36679 20181 36688
rect 19947 36224 19989 36233
rect 19947 36184 19948 36224
rect 19988 36184 19989 36224
rect 19947 36175 19989 36184
rect 18700 35888 18740 35897
rect 18604 35848 18700 35888
rect 18315 35300 18357 35309
rect 18315 35260 18316 35300
rect 18356 35260 18357 35300
rect 18315 35251 18357 35260
rect 18219 33788 18261 33797
rect 18219 33748 18220 33788
rect 18260 33748 18261 33788
rect 18219 33739 18261 33748
rect 18219 33452 18261 33461
rect 18219 33412 18220 33452
rect 18260 33412 18261 33452
rect 18219 33403 18261 33412
rect 18220 32878 18260 33403
rect 18220 32829 18260 32838
rect 18316 32705 18356 35251
rect 18604 34376 18644 35848
rect 18700 35839 18740 35848
rect 18988 35216 19028 36091
rect 19180 35893 19220 35902
rect 19180 35393 19220 35853
rect 19179 35384 19221 35393
rect 19179 35344 19180 35384
rect 19220 35344 19221 35384
rect 19179 35335 19221 35344
rect 18988 35141 19028 35176
rect 18987 35132 19029 35141
rect 18987 35092 18988 35132
rect 19028 35092 19029 35132
rect 18987 35083 19029 35092
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 18508 34336 18604 34376
rect 19132 34385 19172 34394
rect 19276 34376 19316 36100
rect 19756 36091 19796 36100
rect 20140 36140 20180 36679
rect 20140 36091 20180 36100
rect 20043 36056 20085 36065
rect 20043 36016 20044 36056
rect 20084 36016 20085 36056
rect 20043 36007 20085 36016
rect 19563 35972 19605 35981
rect 19563 35932 19564 35972
rect 19604 35932 19605 35972
rect 19563 35923 19605 35932
rect 19948 35972 19988 35981
rect 19564 35838 19604 35923
rect 19851 35804 19893 35813
rect 19948 35804 19988 35932
rect 19851 35764 19852 35804
rect 19892 35764 19988 35804
rect 19851 35755 19893 35764
rect 19372 35720 19412 35729
rect 19755 35720 19797 35729
rect 20044 35720 20084 36007
rect 19412 35680 19604 35720
rect 19372 35671 19412 35680
rect 19468 35132 19508 35141
rect 19372 35092 19468 35132
rect 19372 34553 19412 35092
rect 19468 35083 19508 35092
rect 19467 34712 19509 34721
rect 19467 34672 19468 34712
rect 19508 34672 19509 34712
rect 19467 34663 19509 34672
rect 19371 34544 19413 34553
rect 19371 34504 19372 34544
rect 19412 34504 19413 34544
rect 19371 34495 19413 34504
rect 19468 34460 19508 34663
rect 19564 34460 19604 35680
rect 19755 35680 19756 35720
rect 19796 35680 19797 35720
rect 19755 35671 19797 35680
rect 19948 35680 20084 35720
rect 19659 35048 19701 35057
rect 19659 35008 19660 35048
rect 19700 35008 19701 35048
rect 19659 34999 19701 35008
rect 19660 34914 19700 34999
rect 19660 34628 19700 34637
rect 19756 34628 19796 35671
rect 19851 35636 19893 35645
rect 19851 35596 19852 35636
rect 19892 35596 19893 35636
rect 19851 35587 19893 35596
rect 19852 35132 19892 35587
rect 19852 35083 19892 35092
rect 19948 35048 19988 35680
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 20523 35384 20565 35393
rect 20523 35344 20524 35384
rect 20564 35344 20565 35384
rect 20523 35335 20565 35344
rect 20044 35048 20084 35057
rect 19948 35008 20044 35048
rect 20044 34999 20084 35008
rect 19700 34588 19796 34628
rect 19660 34579 19700 34588
rect 19852 34460 19892 34469
rect 19564 34420 19852 34460
rect 19468 34411 19508 34420
rect 19852 34411 19892 34420
rect 19172 34345 19220 34376
rect 19132 34336 19220 34345
rect 19276 34336 19412 34376
rect 18411 33704 18453 33713
rect 18411 33664 18412 33704
rect 18452 33664 18453 33704
rect 18411 33655 18453 33664
rect 18412 33570 18452 33655
rect 18411 32780 18453 32789
rect 18411 32740 18412 32780
rect 18452 32740 18453 32780
rect 18411 32731 18453 32740
rect 18315 32696 18357 32705
rect 18315 32656 18316 32696
rect 18356 32656 18357 32696
rect 18315 32647 18357 32656
rect 18412 32646 18452 32731
rect 18124 32488 18452 32528
rect 18316 31352 18356 31361
rect 18123 31268 18165 31277
rect 18123 31228 18124 31268
rect 18164 31228 18165 31268
rect 18123 31219 18165 31228
rect 18124 30437 18164 31219
rect 18123 30428 18165 30437
rect 18123 30388 18124 30428
rect 18164 30388 18260 30428
rect 18123 30379 18165 30388
rect 18220 29924 18260 30388
rect 18316 30101 18356 31312
rect 18315 30092 18357 30101
rect 18315 30052 18316 30092
rect 18356 30052 18357 30092
rect 18315 30043 18357 30052
rect 18412 29924 18452 32488
rect 18220 29875 18260 29884
rect 18316 29884 18452 29924
rect 18124 29840 18164 29849
rect 18124 29756 18164 29800
rect 18124 29716 18260 29756
rect 18123 29504 18165 29513
rect 18123 29464 18124 29504
rect 18164 29464 18165 29504
rect 18123 29455 18165 29464
rect 18027 29336 18069 29345
rect 18027 29296 18028 29336
rect 18068 29296 18069 29336
rect 18027 29287 18069 29296
rect 17931 29168 17973 29177
rect 17931 29128 17932 29168
rect 17972 29128 17973 29168
rect 17931 29119 17973 29128
rect 18028 29154 18068 29163
rect 17835 29084 17877 29093
rect 17835 29044 17836 29084
rect 17876 29044 17877 29084
rect 17835 29035 17877 29044
rect 17452 28960 17684 29000
rect 17355 28664 17397 28673
rect 17355 28624 17356 28664
rect 17396 28624 17397 28664
rect 17355 28615 17397 28624
rect 17259 28412 17301 28421
rect 17259 28372 17260 28412
rect 17300 28372 17301 28412
rect 17259 28363 17301 28372
rect 17356 28328 17396 28615
rect 17356 28279 17396 28288
rect 17355 28160 17397 28169
rect 17355 28120 17356 28160
rect 17396 28120 17397 28160
rect 17355 28111 17397 28120
rect 17356 27740 17396 28111
rect 17452 27908 17492 28960
rect 17547 28328 17589 28337
rect 17547 28288 17548 28328
rect 17588 28288 17589 28328
rect 17547 28279 17589 28288
rect 17548 28194 17588 28279
rect 17452 27868 17588 27908
rect 17452 27740 17492 27749
rect 17356 27700 17452 27740
rect 17452 27691 17492 27700
rect 17260 27404 17300 27413
rect 17260 27161 17300 27364
rect 17259 27152 17301 27161
rect 17259 27112 17260 27152
rect 17300 27112 17301 27152
rect 17259 27103 17301 27112
rect 17451 27152 17493 27161
rect 17451 27112 17452 27152
rect 17492 27112 17493 27152
rect 17451 27103 17493 27112
rect 17355 26900 17397 26909
rect 17355 26860 17356 26900
rect 17396 26860 17397 26900
rect 17355 26851 17397 26860
rect 17260 26816 17300 26825
rect 17260 26321 17300 26776
rect 17356 26816 17396 26851
rect 17259 26312 17301 26321
rect 17259 26272 17260 26312
rect 17300 26272 17301 26312
rect 17259 26263 17301 26272
rect 17260 26144 17300 26153
rect 17260 25985 17300 26104
rect 17259 25976 17301 25985
rect 17259 25936 17260 25976
rect 17300 25936 17301 25976
rect 17259 25927 17301 25936
rect 17356 25808 17396 26776
rect 17260 25768 17396 25808
rect 17260 25481 17300 25768
rect 17452 25724 17492 27103
rect 17356 25684 17492 25724
rect 17259 25472 17301 25481
rect 17259 25432 17260 25472
rect 17300 25432 17301 25472
rect 17259 25423 17301 25432
rect 17356 25313 17396 25684
rect 17452 25556 17492 25565
rect 17548 25556 17588 27868
rect 17492 25516 17588 25556
rect 17644 27642 17684 27651
rect 17452 25507 17492 25516
rect 17644 25481 17684 27602
rect 17740 26816 17780 26825
rect 17740 26573 17780 26776
rect 17836 26816 17876 29035
rect 17931 28916 17973 28925
rect 17931 28876 17932 28916
rect 17972 28876 17973 28916
rect 17931 28867 17973 28876
rect 17739 26564 17781 26573
rect 17739 26524 17740 26564
rect 17780 26524 17781 26564
rect 17739 26515 17781 26524
rect 17739 25640 17781 25649
rect 17739 25600 17740 25640
rect 17780 25600 17781 25640
rect 17739 25591 17781 25600
rect 17643 25472 17685 25481
rect 17643 25432 17644 25472
rect 17684 25432 17685 25472
rect 17643 25423 17685 25432
rect 17451 25388 17493 25397
rect 17451 25348 17452 25388
rect 17492 25348 17493 25388
rect 17451 25339 17493 25348
rect 17252 25304 17300 25313
rect 17252 25264 17253 25304
rect 17252 25255 17300 25264
rect 17355 25304 17397 25313
rect 17355 25264 17356 25304
rect 17396 25264 17397 25304
rect 17355 25255 17397 25264
rect 17253 25176 17293 25255
rect 17355 24464 17397 24473
rect 17355 24424 17356 24464
rect 17396 24424 17397 24464
rect 17355 24415 17397 24424
rect 17356 23969 17396 24415
rect 17355 23960 17397 23969
rect 17164 23920 17300 23960
rect 17164 23792 17204 23801
rect 17164 23633 17204 23752
rect 17163 23624 17205 23633
rect 17163 23584 17164 23624
rect 17204 23584 17205 23624
rect 17163 23575 17205 23584
rect 17260 23120 17300 23920
rect 17355 23920 17356 23960
rect 17396 23920 17397 23960
rect 17355 23911 17397 23920
rect 17356 23826 17396 23911
rect 17452 23624 17492 25339
rect 17644 25304 17684 25313
rect 17740 25304 17780 25591
rect 17684 25264 17780 25304
rect 17644 25255 17684 25264
rect 17547 25220 17589 25229
rect 17547 25180 17548 25220
rect 17588 25180 17589 25220
rect 17547 25171 17589 25180
rect 17548 24627 17588 25171
rect 17548 24578 17588 24587
rect 17740 24716 17780 24725
rect 17547 23960 17589 23969
rect 17547 23920 17548 23960
rect 17588 23920 17589 23960
rect 17547 23911 17589 23920
rect 17548 23792 17588 23911
rect 17548 23743 17588 23752
rect 17740 23792 17780 24676
rect 17740 23743 17780 23752
rect 17644 23624 17684 23633
rect 17452 23584 17588 23624
rect 17451 23204 17493 23213
rect 17451 23164 17452 23204
rect 17492 23164 17493 23204
rect 17451 23155 17493 23164
rect 17452 23120 17492 23155
rect 17260 23080 17396 23120
rect 16875 23036 16917 23045
rect 16875 22996 16876 23036
rect 16916 22996 16917 23036
rect 16875 22987 16917 22996
rect 16684 22072 16820 22112
rect 16684 20861 16724 22072
rect 16972 21953 17012 23080
rect 17259 22952 17301 22961
rect 17259 22912 17260 22952
rect 17300 22912 17301 22952
rect 17259 22903 17301 22912
rect 17260 22818 17300 22903
rect 16971 21944 17013 21953
rect 16971 21904 16972 21944
rect 17012 21904 17013 21944
rect 16971 21895 17013 21904
rect 17067 21692 17109 21701
rect 17067 21652 17068 21692
rect 17108 21652 17109 21692
rect 17067 21643 17109 21652
rect 16780 21608 16820 21617
rect 16683 20852 16725 20861
rect 16683 20812 16684 20852
rect 16724 20812 16725 20852
rect 16683 20803 16725 20812
rect 16780 20768 16820 21568
rect 16875 21608 16917 21617
rect 16875 21568 16876 21608
rect 16916 21568 16917 21608
rect 16875 21559 16917 21568
rect 16876 21188 16916 21559
rect 16972 21365 17012 21450
rect 17068 21440 17108 21643
rect 17164 21617 17204 21702
rect 17163 21608 17205 21617
rect 17163 21568 17164 21608
rect 17204 21568 17205 21608
rect 17163 21559 17205 21568
rect 17260 21608 17300 21619
rect 17260 21533 17300 21568
rect 17259 21524 17301 21533
rect 17259 21484 17260 21524
rect 17300 21484 17301 21524
rect 17259 21475 17301 21484
rect 17164 21440 17204 21449
rect 17068 21400 17164 21440
rect 17164 21391 17204 21400
rect 16971 21356 17013 21365
rect 16971 21316 16972 21356
rect 17012 21316 17013 21356
rect 16971 21307 17013 21316
rect 17163 21272 17205 21281
rect 17163 21232 17164 21272
rect 17204 21232 17205 21272
rect 17163 21223 17205 21232
rect 16876 21148 17108 21188
rect 17068 21020 17108 21148
rect 17068 20971 17108 20980
rect 16876 20768 16916 20777
rect 16780 20728 16876 20768
rect 16916 20728 17012 20768
rect 16876 20719 16916 20728
rect 16972 20684 17012 20728
rect 16972 20644 17108 20684
rect 16875 20600 16917 20609
rect 16875 20560 16876 20600
rect 16916 20560 16917 20600
rect 16875 20551 16917 20560
rect 16683 18668 16725 18677
rect 16683 18628 16684 18668
rect 16724 18628 16725 18668
rect 16683 18619 16725 18628
rect 16684 18534 16724 18619
rect 16779 18248 16821 18257
rect 16779 18208 16780 18248
rect 16820 18208 16821 18248
rect 16779 18199 16821 18208
rect 16780 17996 16820 18199
rect 16588 17956 16724 17996
rect 16587 17828 16629 17837
rect 16587 17788 16588 17828
rect 16628 17788 16629 17828
rect 16587 17779 16629 17788
rect 16588 17694 16628 17779
rect 16588 17240 16628 17249
rect 16492 17200 16588 17240
rect 16395 17191 16437 17200
rect 16588 17191 16628 17200
rect 16396 17072 16436 17083
rect 16396 16997 16436 17032
rect 16395 16988 16437 16997
rect 16395 16948 16396 16988
rect 16436 16948 16437 16988
rect 16395 16939 16437 16948
rect 16684 16400 16724 17956
rect 16780 17947 16820 17956
rect 16876 16400 16916 20551
rect 17068 20096 17108 20644
rect 16971 20012 17013 20021
rect 16971 19972 16972 20012
rect 17012 19972 17013 20012
rect 16971 19963 17013 19972
rect 16972 18752 17012 19963
rect 17068 19769 17108 20056
rect 17067 19760 17109 19769
rect 17067 19720 17068 19760
rect 17108 19720 17109 19760
rect 17067 19711 17109 19720
rect 17068 19256 17108 19711
rect 17068 19181 17108 19216
rect 17067 19172 17109 19181
rect 17067 19132 17068 19172
rect 17108 19132 17109 19172
rect 17067 19123 17109 19132
rect 17164 18752 17204 21223
rect 17259 20852 17301 20861
rect 17259 20812 17260 20852
rect 17300 20812 17301 20852
rect 17259 20803 17301 20812
rect 17260 20718 17300 20803
rect 17356 20609 17396 23080
rect 17452 23069 17492 23080
rect 17548 22952 17588 23584
rect 17644 23129 17684 23584
rect 17643 23120 17685 23129
rect 17643 23080 17644 23120
rect 17684 23080 17685 23120
rect 17643 23071 17685 23080
rect 17452 22912 17588 22952
rect 17452 21608 17492 22912
rect 17452 21559 17492 21568
rect 17643 21608 17685 21617
rect 17643 21568 17644 21608
rect 17684 21568 17685 21608
rect 17643 21559 17685 21568
rect 17451 21020 17493 21029
rect 17451 20980 17452 21020
rect 17492 20980 17493 21020
rect 17451 20971 17493 20980
rect 17452 20886 17492 20971
rect 17644 20936 17684 21559
rect 17644 20887 17684 20896
rect 17355 20600 17397 20609
rect 17355 20560 17356 20600
rect 17396 20560 17397 20600
rect 17355 20551 17397 20560
rect 17547 20600 17589 20609
rect 17547 20560 17548 20600
rect 17588 20560 17589 20600
rect 17547 20551 17589 20560
rect 17740 20600 17780 20609
rect 17451 20096 17493 20105
rect 17451 20056 17452 20096
rect 17492 20056 17493 20096
rect 17451 20047 17493 20056
rect 17452 19962 17492 20047
rect 17259 19928 17301 19937
rect 17259 19888 17260 19928
rect 17300 19888 17301 19928
rect 17259 19879 17301 19888
rect 17260 19794 17300 19879
rect 17259 19676 17301 19685
rect 17259 19636 17260 19676
rect 17300 19636 17301 19676
rect 17259 19627 17301 19636
rect 17260 19508 17300 19627
rect 17260 19459 17300 19468
rect 17548 19424 17588 20551
rect 17548 19375 17588 19384
rect 17740 19340 17780 20560
rect 17836 19433 17876 26776
rect 17932 25817 17972 28867
rect 17931 25808 17973 25817
rect 17931 25768 17932 25808
rect 17972 25768 17973 25808
rect 17931 25759 17973 25768
rect 17932 25397 17972 25759
rect 18028 25649 18068 29114
rect 18124 27656 18164 29455
rect 18220 29429 18260 29716
rect 18219 29420 18261 29429
rect 18219 29380 18220 29420
rect 18260 29380 18261 29420
rect 18219 29371 18261 29380
rect 18124 26657 18164 27616
rect 18220 29252 18260 29261
rect 18220 27581 18260 29212
rect 18316 28925 18356 29884
rect 18508 29513 18548 34336
rect 18604 34327 18644 34336
rect 18604 33881 18644 33966
rect 18603 33872 18645 33881
rect 18603 33832 18604 33872
rect 18644 33832 18645 33872
rect 18603 33823 18645 33832
rect 19180 33452 19220 34336
rect 19276 34208 19316 34217
rect 19276 33965 19316 34168
rect 19275 33956 19317 33965
rect 19275 33916 19276 33956
rect 19316 33916 19317 33956
rect 19275 33907 19317 33916
rect 19372 33788 19412 34336
rect 19659 34292 19701 34301
rect 19659 34252 19660 34292
rect 19700 34252 19701 34292
rect 19659 34243 19701 34252
rect 19563 33956 19605 33965
rect 19563 33916 19564 33956
rect 19604 33916 19605 33956
rect 19563 33907 19605 33916
rect 19564 33872 19604 33907
rect 19564 33821 19604 33832
rect 19276 33748 19412 33788
rect 19276 33536 19316 33748
rect 19383 33633 19423 33642
rect 19467 33620 19509 33629
rect 19423 33593 19468 33620
rect 19383 33580 19468 33593
rect 19508 33580 19509 33620
rect 19467 33571 19509 33580
rect 19276 33496 19412 33536
rect 19180 33412 19316 33452
rect 18699 33368 18741 33377
rect 18699 33328 18700 33368
rect 18740 33328 18741 33368
rect 18699 33319 18741 33328
rect 18700 33116 18740 33319
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 18796 33116 18836 33125
rect 18700 33076 18796 33116
rect 18796 33067 18836 33076
rect 19179 33116 19221 33125
rect 19179 33076 19180 33116
rect 19220 33076 19221 33116
rect 19179 33067 19221 33076
rect 19180 32982 19220 33067
rect 18603 32948 18645 32957
rect 18603 32908 18604 32948
rect 18644 32908 18645 32948
rect 18603 32899 18645 32908
rect 18988 32948 19028 32957
rect 18604 32814 18644 32899
rect 18795 32864 18837 32873
rect 18795 32824 18796 32864
rect 18836 32824 18837 32864
rect 18795 32815 18837 32824
rect 18603 32192 18645 32201
rect 18603 32152 18604 32192
rect 18644 32152 18645 32192
rect 18603 32143 18645 32152
rect 18796 32192 18836 32815
rect 18988 32537 19028 32908
rect 18987 32528 19029 32537
rect 18987 32488 18988 32528
rect 19028 32488 19029 32528
rect 18987 32479 19029 32488
rect 18796 32143 18836 32152
rect 18604 32058 18644 32143
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 19083 31604 19125 31613
rect 19083 31564 19084 31604
rect 19124 31564 19125 31604
rect 19083 31555 19125 31564
rect 18796 31357 18836 31366
rect 18796 30428 18836 31317
rect 18988 31184 19028 31193
rect 18988 30437 19028 31144
rect 19084 30680 19124 31555
rect 19276 30848 19316 33412
rect 19372 33116 19412 33496
rect 19564 33116 19604 33125
rect 19660 33116 19700 34243
rect 20044 34217 20084 34302
rect 20043 34208 20085 34217
rect 20043 34168 20044 34208
rect 20084 34168 20085 34208
rect 20043 34159 20085 34168
rect 19851 34124 19893 34133
rect 19851 34084 19852 34124
rect 19892 34084 19893 34124
rect 19851 34075 19893 34084
rect 19372 33076 19508 33116
rect 19372 32948 19412 32959
rect 19372 32873 19412 32908
rect 19371 32864 19413 32873
rect 19371 32824 19372 32864
rect 19412 32824 19413 32864
rect 19371 32815 19413 32824
rect 19371 31520 19413 31529
rect 19371 31480 19372 31520
rect 19412 31480 19413 31520
rect 19371 31471 19413 31480
rect 19372 31436 19412 31471
rect 19372 31385 19412 31396
rect 19468 30932 19508 33076
rect 19604 33076 19700 33116
rect 19756 33620 19796 33629
rect 19564 33067 19604 33076
rect 19756 33041 19796 33580
rect 19852 33125 19892 34075
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 19947 33872 19989 33881
rect 19947 33832 19948 33872
rect 19988 33832 19989 33872
rect 19947 33823 19989 33832
rect 19948 33738 19988 33823
rect 20043 33788 20085 33797
rect 20043 33748 20044 33788
rect 20084 33748 20085 33788
rect 20043 33739 20085 33748
rect 19851 33116 19893 33125
rect 19851 33076 19852 33116
rect 19892 33076 19893 33116
rect 19851 33067 19893 33076
rect 19755 33032 19797 33041
rect 19755 32992 19756 33032
rect 19796 32992 19797 33032
rect 19755 32983 19797 32992
rect 19947 33032 19989 33041
rect 19947 32992 19948 33032
rect 19988 32992 19989 33032
rect 19947 32983 19989 32992
rect 19756 32898 19796 32983
rect 19851 32780 19893 32789
rect 19851 32740 19852 32780
rect 19892 32740 19893 32780
rect 19851 32731 19893 32740
rect 19659 32612 19701 32621
rect 19659 32572 19660 32612
rect 19700 32572 19701 32612
rect 19659 32563 19701 32572
rect 19563 31184 19605 31193
rect 19563 31144 19564 31184
rect 19604 31144 19605 31184
rect 19563 31135 19605 31144
rect 19564 31050 19604 31135
rect 19468 30892 19604 30932
rect 19276 30799 19316 30808
rect 19084 30631 19124 30640
rect 19372 30605 19412 30690
rect 19371 30596 19413 30605
rect 19468 30596 19508 30605
rect 19371 30556 19372 30596
rect 19412 30556 19468 30596
rect 19371 30547 19413 30556
rect 19468 30547 19508 30556
rect 18604 30388 18836 30428
rect 18987 30428 19029 30437
rect 19372 30428 19412 30547
rect 18987 30388 18988 30428
rect 19028 30388 19029 30428
rect 18507 29504 18549 29513
rect 18507 29464 18508 29504
rect 18548 29464 18549 29504
rect 18507 29455 18549 29464
rect 18411 29336 18453 29345
rect 18411 29296 18412 29336
rect 18452 29296 18453 29336
rect 18411 29287 18453 29296
rect 18412 29168 18452 29287
rect 18412 29119 18452 29128
rect 18507 29168 18549 29177
rect 18507 29128 18508 29168
rect 18548 29128 18549 29168
rect 18507 29119 18549 29128
rect 18315 28916 18357 28925
rect 18315 28876 18316 28916
rect 18356 28876 18357 28916
rect 18315 28867 18357 28876
rect 18315 28664 18357 28673
rect 18315 28624 18316 28664
rect 18356 28624 18357 28664
rect 18315 28615 18357 28624
rect 18219 27572 18261 27581
rect 18219 27532 18220 27572
rect 18260 27532 18261 27572
rect 18219 27523 18261 27532
rect 18316 26816 18356 28615
rect 18508 28328 18548 29119
rect 18604 28589 18644 30388
rect 18987 30379 19029 30388
rect 19362 30388 19412 30428
rect 19467 30428 19509 30437
rect 19467 30388 19468 30428
rect 19508 30388 19509 30428
rect 19362 30344 19402 30388
rect 19467 30379 19509 30388
rect 19362 30304 19412 30344
rect 18699 30260 18741 30269
rect 18699 30220 18700 30260
rect 18740 30220 18741 30260
rect 18699 30211 18741 30220
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 18700 29840 18740 30211
rect 19228 29849 19268 29858
rect 19372 29849 19412 30304
rect 19371 29840 19413 29849
rect 19268 29809 19316 29840
rect 19228 29800 19316 29809
rect 18700 28673 18740 29800
rect 19276 29345 19316 29800
rect 19371 29800 19372 29840
rect 19412 29800 19413 29840
rect 19371 29791 19413 29800
rect 19372 29672 19412 29681
rect 19275 29336 19317 29345
rect 19275 29296 19276 29336
rect 19316 29296 19317 29336
rect 19275 29287 19317 29296
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 18699 28664 18741 28673
rect 18699 28624 18700 28664
rect 18740 28624 18741 28664
rect 18699 28615 18741 28624
rect 18603 28580 18645 28589
rect 18603 28540 18604 28580
rect 18644 28540 18645 28580
rect 18603 28531 18645 28540
rect 18987 28580 19029 28589
rect 18987 28540 18988 28580
rect 19028 28540 19029 28580
rect 18987 28531 19029 28540
rect 18988 28446 19028 28531
rect 19180 28412 19220 28421
rect 19372 28412 19412 29632
rect 19220 28372 19412 28412
rect 19180 28363 19220 28372
rect 18796 28328 18836 28337
rect 18508 28288 18796 28328
rect 18604 27656 18644 27665
rect 18604 27572 18644 27616
rect 18699 27656 18741 27665
rect 18699 27616 18700 27656
rect 18740 27616 18741 27656
rect 18699 27607 18741 27616
rect 18412 27532 18644 27572
rect 18412 27245 18452 27532
rect 18700 27522 18740 27607
rect 18796 27404 18836 28288
rect 19372 28160 19412 28169
rect 19083 28076 19125 28085
rect 19083 28036 19084 28076
rect 19124 28036 19125 28076
rect 19083 28027 19125 28036
rect 19084 27656 19124 28027
rect 19084 27581 19124 27616
rect 19180 27656 19220 27665
rect 19220 27616 19316 27656
rect 19180 27607 19220 27616
rect 19083 27572 19125 27581
rect 19083 27532 19084 27572
rect 19124 27532 19125 27572
rect 19083 27523 19125 27532
rect 18700 27364 18836 27404
rect 18411 27236 18453 27245
rect 18700 27236 18740 27364
rect 18411 27196 18412 27236
rect 18452 27196 18453 27236
rect 18411 27187 18453 27196
rect 18508 27196 18740 27236
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18220 26776 18316 26816
rect 18123 26648 18165 26657
rect 18123 26608 18124 26648
rect 18164 26608 18165 26648
rect 18123 26599 18165 26608
rect 18123 26144 18165 26153
rect 18123 26104 18124 26144
rect 18164 26104 18165 26144
rect 18123 26095 18165 26104
rect 18027 25640 18069 25649
rect 18027 25600 18028 25640
rect 18068 25600 18069 25640
rect 18027 25591 18069 25600
rect 18027 25472 18069 25481
rect 18027 25432 18028 25472
rect 18068 25432 18069 25472
rect 18027 25423 18069 25432
rect 17931 25388 17973 25397
rect 17931 25348 17932 25388
rect 17972 25348 17973 25388
rect 17931 25339 17973 25348
rect 17932 24632 17972 24643
rect 17932 24557 17972 24592
rect 17931 24548 17973 24557
rect 17931 24508 17932 24548
rect 17972 24508 17973 24548
rect 17931 24499 17973 24508
rect 17931 24380 17973 24389
rect 17931 24340 17932 24380
rect 17972 24340 17973 24380
rect 17931 24331 17973 24340
rect 17932 24246 17972 24331
rect 18028 23960 18068 25423
rect 18124 25229 18164 26095
rect 18123 25220 18165 25229
rect 18123 25180 18124 25220
rect 18164 25180 18165 25220
rect 18123 25171 18165 25180
rect 18124 24632 18164 25171
rect 18220 24809 18260 26776
rect 18316 26767 18356 26776
rect 18412 26405 18452 27187
rect 18411 26396 18453 26405
rect 18411 26356 18412 26396
rect 18452 26356 18453 26396
rect 18411 26347 18453 26356
rect 18508 26144 18548 27196
rect 18808 27187 19176 27196
rect 18796 26821 18836 26830
rect 19276 26816 19316 27616
rect 19372 27068 19412 28120
rect 19468 27572 19508 30379
rect 19564 29009 19604 30892
rect 19660 30848 19700 32563
rect 19756 31436 19796 31445
rect 19756 30941 19796 31396
rect 19755 30932 19797 30941
rect 19755 30892 19756 30932
rect 19796 30892 19797 30932
rect 19755 30883 19797 30892
rect 19660 30799 19700 30808
rect 19852 30596 19892 32731
rect 19948 31520 19988 32983
rect 20044 32948 20084 33739
rect 20044 32899 20084 32908
rect 20236 32696 20276 32705
rect 20427 32696 20469 32705
rect 20276 32656 20428 32696
rect 20468 32656 20469 32696
rect 20236 32647 20276 32656
rect 20427 32647 20469 32656
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 20236 32360 20276 32369
rect 20524 32360 20564 35335
rect 21003 32696 21045 32705
rect 21003 32656 21004 32696
rect 21044 32656 21045 32696
rect 21003 32647 21045 32656
rect 20276 32320 20564 32360
rect 20236 32311 20276 32320
rect 20043 32276 20085 32285
rect 20043 32236 20044 32276
rect 20084 32236 20085 32276
rect 20043 32227 20085 32236
rect 20044 32192 20084 32227
rect 20044 32141 20084 32152
rect 20523 31688 20565 31697
rect 20523 31648 20524 31688
rect 20564 31648 20565 31688
rect 20523 31639 20565 31648
rect 19948 31471 19988 31480
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 20524 30680 20564 31639
rect 19852 30547 19892 30556
rect 20236 30640 20564 30680
rect 20619 30680 20661 30689
rect 20619 30640 20620 30680
rect 20660 30640 20661 30680
rect 20044 30428 20084 30437
rect 19948 30388 20044 30428
rect 19755 30176 19797 30185
rect 19755 30136 19756 30176
rect 19796 30136 19797 30176
rect 19755 30127 19797 30136
rect 19660 29924 19700 29933
rect 19660 29765 19700 29884
rect 19659 29756 19701 29765
rect 19659 29716 19660 29756
rect 19700 29716 19701 29756
rect 19659 29707 19701 29716
rect 19756 29177 19796 30127
rect 19851 30092 19893 30101
rect 19851 30052 19852 30092
rect 19892 30052 19893 30092
rect 19851 30043 19893 30052
rect 19852 29958 19892 30043
rect 19851 29840 19893 29849
rect 19851 29800 19852 29840
rect 19892 29800 19893 29840
rect 19851 29791 19893 29800
rect 19852 29504 19892 29791
rect 19948 29681 19988 30388
rect 20044 30379 20084 30388
rect 20236 30092 20276 30640
rect 20619 30631 20661 30640
rect 20236 30043 20276 30052
rect 20043 29924 20085 29933
rect 20043 29884 20044 29924
rect 20084 29884 20085 29924
rect 20043 29875 20085 29884
rect 20044 29790 20084 29875
rect 19947 29672 19989 29681
rect 19947 29632 19948 29672
rect 19988 29632 19989 29672
rect 19947 29623 19989 29632
rect 20048 29504 20416 29513
rect 19852 29464 19988 29504
rect 19851 29336 19893 29345
rect 19851 29296 19852 29336
rect 19892 29296 19893 29336
rect 19851 29287 19893 29296
rect 19852 29202 19892 29287
rect 19755 29168 19797 29177
rect 19660 29126 19700 29135
rect 19659 29086 19660 29093
rect 19755 29128 19756 29168
rect 19796 29128 19797 29168
rect 19755 29119 19797 29128
rect 19700 29086 19701 29093
rect 19659 29084 19701 29086
rect 19659 29044 19660 29084
rect 19700 29044 19701 29084
rect 19659 29035 19701 29044
rect 19563 29000 19605 29009
rect 19563 28960 19564 29000
rect 19604 28960 19605 29000
rect 19660 28991 19700 29035
rect 19563 28951 19605 28960
rect 19659 28916 19701 28925
rect 19659 28876 19660 28916
rect 19700 28876 19701 28916
rect 19659 28867 19701 28876
rect 19563 28832 19605 28841
rect 19563 28792 19564 28832
rect 19604 28792 19605 28832
rect 19563 28783 19605 28792
rect 19564 28412 19604 28783
rect 19564 28363 19604 28372
rect 19660 28337 19700 28867
rect 19755 28580 19797 28589
rect 19755 28540 19756 28580
rect 19796 28540 19797 28580
rect 19948 28580 19988 29464
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 20620 29336 20660 30631
rect 20715 30008 20757 30017
rect 20715 29968 20716 30008
rect 20756 29968 20757 30008
rect 20715 29959 20757 29968
rect 20140 29296 20660 29336
rect 20043 29168 20085 29177
rect 20043 29128 20044 29168
rect 20084 29128 20085 29168
rect 20043 29119 20085 29128
rect 20044 29084 20084 29119
rect 20044 29033 20084 29044
rect 20140 28580 20180 29296
rect 20236 28916 20276 28925
rect 20276 28876 20564 28916
rect 20236 28867 20276 28876
rect 19948 28540 20084 28580
rect 19755 28531 19797 28540
rect 19756 28446 19796 28531
rect 19851 28496 19893 28505
rect 19851 28456 19852 28496
rect 19892 28456 19893 28496
rect 19851 28447 19893 28456
rect 19659 28328 19701 28337
rect 19659 28288 19660 28328
rect 19700 28288 19701 28328
rect 19659 28279 19701 28288
rect 19659 27908 19701 27917
rect 19659 27868 19660 27908
rect 19700 27868 19701 27908
rect 19659 27859 19701 27868
rect 19468 27523 19508 27532
rect 19660 27488 19700 27859
rect 19852 27572 19892 28447
rect 19947 28412 19989 28421
rect 19947 28372 19948 28412
rect 19988 28372 19989 28412
rect 19947 28363 19989 28372
rect 19948 28278 19988 28363
rect 20044 28160 20084 28540
rect 20140 28531 20180 28540
rect 19852 27523 19892 27532
rect 19948 28120 20084 28160
rect 19660 27439 19700 27448
rect 19755 27404 19797 27413
rect 19755 27364 19756 27404
rect 19796 27364 19797 27404
rect 19755 27355 19797 27364
rect 19372 27028 19508 27068
rect 19371 26900 19413 26909
rect 19371 26860 19372 26900
rect 19412 26860 19413 26900
rect 19371 26851 19413 26860
rect 18699 26312 18741 26321
rect 18699 26272 18700 26312
rect 18740 26272 18741 26312
rect 18699 26263 18741 26272
rect 18700 26178 18740 26263
rect 18316 26104 18508 26144
rect 18316 25565 18356 26104
rect 18508 26095 18548 26104
rect 18796 25892 18836 26781
rect 18892 26776 19316 26816
rect 18892 26321 18932 26776
rect 19372 26766 19412 26851
rect 19468 26741 19508 27028
rect 19756 26900 19796 27355
rect 19756 26851 19796 26860
rect 19948 26816 19988 28120
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 20043 27824 20085 27833
rect 20043 27784 20044 27824
rect 20084 27784 20085 27824
rect 20043 27775 20085 27784
rect 20044 27690 20084 27775
rect 20524 26993 20564 28876
rect 20716 27749 20756 29959
rect 20715 27740 20757 27749
rect 20715 27700 20716 27740
rect 20756 27700 20757 27740
rect 20715 27691 20757 27700
rect 20523 26984 20565 26993
rect 20523 26944 20524 26984
rect 20564 26944 20565 26984
rect 20523 26935 20565 26944
rect 19852 26776 19988 26816
rect 19467 26732 19509 26741
rect 19467 26692 19468 26732
rect 19508 26692 19509 26732
rect 19467 26683 19509 26692
rect 18988 26648 19028 26657
rect 19563 26648 19605 26657
rect 19028 26608 19412 26648
rect 18988 26599 19028 26608
rect 18987 26480 19029 26489
rect 18987 26440 18988 26480
rect 19028 26440 19029 26480
rect 18987 26431 19029 26440
rect 18891 26312 18933 26321
rect 18891 26272 18892 26312
rect 18932 26272 18933 26312
rect 18891 26263 18933 26272
rect 18891 26144 18933 26153
rect 18891 26104 18892 26144
rect 18932 26104 18933 26144
rect 18891 26095 18933 26104
rect 18988 26144 19028 26431
rect 19275 26396 19317 26405
rect 19275 26356 19276 26396
rect 19316 26356 19317 26396
rect 19275 26347 19317 26356
rect 18988 26095 19028 26104
rect 19180 26312 19220 26321
rect 18892 26010 18932 26095
rect 19180 25901 19220 26272
rect 18700 25852 18836 25892
rect 19179 25892 19221 25901
rect 19179 25852 19180 25892
rect 19220 25852 19221 25892
rect 19276 25892 19316 26347
rect 19372 26060 19412 26608
rect 19563 26608 19564 26648
rect 19604 26608 19605 26648
rect 19563 26599 19605 26608
rect 19564 26514 19604 26599
rect 19852 26396 19892 26776
rect 19947 26648 19989 26657
rect 19947 26608 19948 26648
rect 19988 26608 19989 26648
rect 19947 26599 19989 26608
rect 20811 26648 20853 26657
rect 20811 26608 20812 26648
rect 20852 26608 20853 26648
rect 20811 26599 20853 26608
rect 19948 26514 19988 26599
rect 20523 26564 20565 26573
rect 20523 26524 20524 26564
rect 20564 26524 20565 26564
rect 20523 26515 20565 26524
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 19372 26011 19412 26020
rect 19468 26356 19892 26396
rect 19276 25852 19412 25892
rect 18315 25556 18357 25565
rect 18315 25516 18316 25556
rect 18356 25516 18357 25556
rect 18315 25507 18357 25516
rect 18219 24800 18261 24809
rect 18219 24760 18220 24800
rect 18260 24760 18261 24800
rect 18219 24751 18261 24760
rect 18124 24583 18164 24592
rect 18220 24632 18260 24641
rect 18124 23960 18164 23969
rect 18028 23920 18124 23960
rect 18124 23911 18164 23920
rect 18123 23120 18165 23129
rect 18123 23080 18124 23120
rect 18164 23080 18165 23120
rect 18123 23071 18165 23080
rect 18124 22532 18164 23071
rect 18220 22961 18260 24592
rect 18316 23792 18356 25507
rect 18411 25220 18453 25229
rect 18411 25180 18412 25220
rect 18452 25180 18453 25220
rect 18411 25171 18453 25180
rect 18219 22952 18261 22961
rect 18219 22912 18220 22952
rect 18260 22912 18261 22952
rect 18219 22903 18261 22912
rect 18124 22483 18164 22492
rect 17931 22448 17973 22457
rect 17931 22408 17932 22448
rect 17972 22408 17973 22448
rect 17931 22399 17973 22408
rect 17932 22280 17972 22399
rect 17932 22231 17972 22240
rect 18023 20777 18063 20862
rect 18022 20768 18064 20777
rect 18022 20728 18023 20768
rect 18063 20728 18064 20768
rect 18022 20719 18064 20728
rect 18124 20768 18164 20777
rect 18028 20600 18068 20609
rect 17931 19592 17973 19601
rect 17931 19552 17932 19592
rect 17972 19552 17973 19592
rect 17931 19543 17973 19552
rect 17835 19424 17877 19433
rect 17835 19384 17836 19424
rect 17876 19384 17877 19424
rect 17835 19375 17877 19384
rect 17737 19300 17780 19340
rect 17547 19256 17589 19265
rect 17547 19216 17548 19256
rect 17588 19216 17589 19256
rect 17547 19207 17589 19216
rect 16972 18703 17012 18712
rect 17068 18712 17204 18752
rect 17260 19088 17300 19097
rect 16971 18500 17013 18509
rect 16971 18460 16972 18500
rect 17012 18460 17013 18500
rect 16971 18451 17013 18460
rect 16972 17828 17012 18451
rect 16972 17779 17012 17788
rect 16971 17492 17013 17501
rect 16971 17452 16972 17492
rect 17012 17452 17013 17492
rect 16971 17443 17013 17452
rect 16972 16988 17012 17443
rect 16972 16939 17012 16948
rect 16492 16360 16724 16400
rect 16780 16360 16916 16400
rect 16299 14132 16341 14141
rect 16299 14092 16300 14132
rect 16340 14092 16341 14132
rect 16299 14083 16341 14092
rect 15820 14048 15860 14057
rect 15724 14008 15820 14048
rect 15723 13880 15765 13889
rect 15723 13840 15724 13880
rect 15764 13840 15765 13880
rect 15723 13831 15765 13840
rect 15531 13124 15573 13133
rect 15531 13084 15532 13124
rect 15572 13084 15573 13124
rect 15531 13075 15573 13084
rect 15532 13044 15572 13075
rect 15147 12704 15189 12713
rect 15147 12664 15148 12704
rect 15188 12664 15189 12704
rect 15147 12655 15189 12664
rect 15340 12620 15380 12629
rect 15380 12580 15476 12620
rect 15340 12571 15380 12580
rect 14860 12536 14900 12545
rect 14860 11957 14900 12496
rect 14955 12536 14997 12545
rect 14955 12496 14956 12536
rect 14996 12496 14997 12536
rect 14955 12487 14997 12496
rect 15148 12536 15188 12545
rect 15188 12496 15284 12536
rect 15148 12487 15188 12496
rect 14956 12402 14996 12487
rect 15147 12368 15189 12377
rect 15147 12328 15148 12368
rect 15188 12328 15189 12368
rect 15147 12319 15189 12328
rect 15148 12234 15188 12319
rect 14859 11948 14901 11957
rect 14859 11908 14860 11948
rect 14900 11908 14901 11948
rect 14859 11899 14901 11908
rect 15147 11864 15189 11873
rect 15052 11824 15148 11864
rect 15188 11824 15189 11864
rect 15052 11444 15092 11824
rect 15147 11815 15189 11824
rect 15147 11696 15189 11705
rect 15147 11656 15148 11696
rect 15188 11656 15189 11696
rect 15147 11647 15189 11656
rect 15148 11562 15188 11647
rect 15052 11404 15188 11444
rect 14764 11320 14996 11360
rect 14860 11010 14900 11019
rect 14667 10940 14709 10949
rect 14667 10900 14668 10940
rect 14708 10900 14709 10940
rect 14667 10891 14709 10900
rect 14572 10135 14612 10144
rect 14668 9689 14708 10891
rect 14764 10436 14804 10445
rect 14860 10436 14900 10970
rect 14956 10940 14996 11320
rect 15052 11117 15092 11202
rect 15051 11108 15093 11117
rect 15051 11068 15052 11108
rect 15092 11068 15093 11108
rect 15051 11059 15093 11068
rect 14956 10900 15092 10940
rect 14804 10396 14900 10436
rect 14764 10387 14804 10396
rect 14956 10184 14996 10193
rect 14860 10144 14956 10184
rect 14860 9773 14900 10144
rect 14956 10135 14996 10144
rect 15052 10184 15092 10900
rect 15052 10135 15092 10144
rect 14955 9848 14997 9857
rect 14955 9808 14956 9848
rect 14996 9808 14997 9848
rect 14955 9799 14997 9808
rect 14859 9764 14901 9773
rect 14859 9724 14860 9764
rect 14900 9724 14901 9764
rect 14859 9715 14901 9724
rect 14476 9631 14516 9640
rect 14667 9680 14709 9689
rect 14667 9640 14668 9680
rect 14708 9640 14709 9680
rect 14667 9631 14709 9640
rect 14860 9521 14900 9715
rect 14572 9512 14612 9521
rect 14380 9463 14420 9472
rect 14476 9472 14572 9512
rect 14476 8177 14516 9472
rect 14572 9463 14612 9472
rect 14668 9512 14708 9521
rect 14571 9344 14613 9353
rect 14571 9304 14572 9344
rect 14612 9304 14613 9344
rect 14571 9295 14613 9304
rect 14572 8672 14612 9295
rect 14668 8849 14708 9472
rect 14823 9512 14900 9521
rect 14863 9472 14900 9512
rect 14823 9463 14900 9472
rect 14764 8924 14804 8933
rect 14860 8924 14900 9463
rect 14804 8884 14900 8924
rect 14764 8875 14804 8884
rect 14667 8840 14709 8849
rect 14667 8800 14668 8840
rect 14708 8800 14709 8840
rect 14667 8791 14709 8800
rect 14612 8632 14708 8672
rect 14572 8623 14612 8632
rect 14475 8168 14517 8177
rect 14475 8128 14476 8168
rect 14516 8128 14517 8168
rect 14475 8119 14517 8128
rect 14668 8000 14708 8632
rect 14859 8168 14901 8177
rect 14859 8128 14860 8168
rect 14900 8128 14901 8168
rect 14859 8119 14901 8128
rect 14860 8034 14900 8119
rect 14708 7960 14804 8000
rect 14668 7951 14708 7960
rect 14188 7288 14324 7328
rect 14188 7165 14228 7174
rect 14091 6908 14133 6917
rect 14091 6868 14092 6908
rect 14132 6868 14133 6908
rect 14091 6859 14133 6868
rect 14188 6656 14228 7125
rect 14188 6607 14228 6616
rect 13419 6572 13461 6581
rect 13419 6532 13420 6572
rect 13460 6532 13461 6572
rect 13419 6523 13461 6532
rect 13420 5648 13460 6523
rect 13995 6488 14037 6497
rect 13995 6448 13996 6488
rect 14036 6448 14037 6488
rect 13995 6439 14037 6448
rect 13996 6329 14036 6439
rect 13995 6320 14037 6329
rect 13995 6280 13996 6320
rect 14036 6280 14037 6320
rect 13995 6271 14037 6280
rect 13420 5599 13460 5608
rect 13803 2708 13845 2717
rect 13803 2668 13804 2708
rect 13844 2668 13845 2708
rect 13803 2659 13845 2668
rect 13804 2574 13844 2659
rect 14284 2465 14324 7288
rect 14379 6992 14421 7001
rect 14379 6952 14380 6992
rect 14420 6952 14421 6992
rect 14379 6943 14421 6952
rect 14380 6858 14420 6943
rect 14667 6236 14709 6245
rect 14667 6196 14668 6236
rect 14708 6196 14709 6236
rect 14667 6187 14709 6196
rect 14668 5648 14708 6187
rect 14668 5599 14708 5608
rect 14764 5069 14804 7960
rect 14859 7160 14901 7169
rect 14859 7120 14860 7160
rect 14900 7120 14901 7160
rect 14859 7111 14901 7120
rect 14860 5900 14900 7111
rect 14956 6665 14996 9799
rect 15052 9344 15092 9353
rect 15052 8504 15092 9304
rect 15148 9092 15188 11404
rect 15244 10856 15284 12496
rect 15339 11612 15381 11621
rect 15339 11572 15340 11612
rect 15380 11572 15381 11612
rect 15339 11563 15381 11572
rect 15340 11478 15380 11563
rect 15436 11024 15476 12580
rect 15532 12522 15572 12531
rect 15532 11696 15572 12482
rect 15628 12293 15668 13168
rect 15724 13049 15764 13831
rect 15820 13217 15860 14008
rect 15916 14048 15956 14057
rect 15956 14008 16052 14048
rect 15916 13999 15956 14008
rect 15915 13880 15957 13889
rect 15915 13840 15916 13880
rect 15956 13840 15957 13880
rect 15915 13831 15957 13840
rect 15916 13460 15956 13831
rect 16012 13805 16052 14008
rect 16300 13964 16340 13973
rect 16204 13924 16300 13964
rect 16011 13796 16053 13805
rect 16011 13756 16012 13796
rect 16052 13756 16053 13796
rect 16011 13747 16053 13756
rect 15916 13411 15956 13420
rect 16204 13376 16244 13924
rect 16300 13915 16340 13924
rect 16396 13964 16436 13973
rect 16299 13796 16341 13805
rect 16299 13756 16300 13796
rect 16340 13756 16341 13796
rect 16299 13747 16341 13756
rect 16012 13336 16244 13376
rect 15819 13208 15861 13217
rect 15819 13168 15820 13208
rect 15860 13168 15861 13208
rect 15819 13159 15861 13168
rect 15723 13040 15765 13049
rect 15723 13000 15724 13040
rect 15764 13000 15765 13040
rect 15723 12991 15765 13000
rect 15819 12704 15861 12713
rect 16012 12704 16052 13336
rect 16203 13208 16245 13217
rect 16203 13168 16204 13208
rect 16244 13168 16245 13208
rect 16203 13159 16245 13168
rect 16107 13124 16149 13133
rect 16107 13084 16108 13124
rect 16148 13084 16149 13124
rect 16107 13075 16149 13084
rect 15819 12664 15820 12704
rect 15860 12664 15861 12704
rect 15819 12655 15861 12664
rect 15916 12664 16052 12704
rect 15627 12284 15669 12293
rect 15627 12244 15628 12284
rect 15668 12244 15669 12284
rect 15627 12235 15669 12244
rect 15724 11705 15764 11790
rect 15723 11696 15765 11705
rect 15532 11656 15668 11696
rect 15531 11528 15573 11537
rect 15531 11488 15532 11528
rect 15572 11488 15573 11528
rect 15628 11528 15668 11656
rect 15723 11656 15724 11696
rect 15764 11656 15765 11696
rect 15723 11647 15765 11656
rect 15628 11488 15764 11528
rect 15531 11479 15573 11488
rect 15532 11360 15572 11479
rect 15532 11320 15668 11360
rect 15436 10975 15476 10984
rect 15628 11024 15668 11320
rect 15724 11033 15764 11488
rect 15628 10975 15668 10984
rect 15723 11024 15765 11033
rect 15723 10984 15724 11024
rect 15764 10984 15765 11024
rect 15723 10975 15765 10984
rect 15436 10856 15476 10865
rect 15244 10816 15436 10856
rect 15436 10807 15476 10816
rect 15723 10184 15765 10193
rect 15723 10144 15724 10184
rect 15764 10144 15765 10184
rect 15723 10135 15765 10144
rect 15724 10050 15764 10135
rect 15243 10016 15285 10025
rect 15243 9976 15244 10016
rect 15284 9976 15285 10016
rect 15243 9967 15285 9976
rect 15244 9882 15284 9967
rect 15340 9512 15380 9521
rect 15380 9472 15572 9512
rect 15340 9463 15380 9472
rect 15148 9052 15476 9092
rect 15339 8840 15381 8849
rect 15339 8800 15340 8840
rect 15380 8800 15381 8840
rect 15339 8791 15381 8800
rect 15340 8706 15380 8791
rect 15436 8681 15476 9052
rect 15435 8672 15477 8681
rect 15435 8632 15436 8672
rect 15476 8632 15477 8672
rect 15435 8623 15477 8632
rect 15436 8538 15476 8623
rect 15532 8513 15572 9472
rect 15052 7832 15092 8464
rect 15531 8504 15573 8513
rect 15531 8464 15532 8504
rect 15572 8464 15573 8504
rect 15531 8455 15573 8464
rect 15052 7589 15092 7792
rect 15051 7580 15093 7589
rect 15051 7540 15052 7580
rect 15092 7540 15093 7580
rect 15051 7531 15093 7540
rect 15052 7328 15092 7531
rect 14955 6656 14997 6665
rect 14955 6616 14956 6656
rect 14996 6616 14997 6656
rect 14955 6607 14997 6616
rect 14860 5851 14900 5860
rect 15052 6488 15092 7288
rect 15435 7160 15477 7169
rect 15435 7120 15436 7160
rect 15476 7120 15477 7160
rect 15435 7111 15477 7120
rect 15532 7160 15572 7171
rect 15436 7026 15476 7111
rect 15532 7085 15572 7120
rect 15531 7076 15573 7085
rect 15531 7036 15532 7076
rect 15572 7036 15573 7076
rect 15531 7027 15573 7036
rect 15532 6749 15572 7027
rect 15820 6908 15860 12655
rect 15916 11201 15956 12664
rect 16012 12536 16052 12547
rect 16012 12461 16052 12496
rect 16011 12452 16053 12461
rect 16011 12412 16012 12452
rect 16052 12412 16053 12452
rect 16011 12403 16053 12412
rect 16011 12284 16053 12293
rect 16011 12244 16012 12284
rect 16052 12244 16053 12284
rect 16011 12235 16053 12244
rect 15915 11192 15957 11201
rect 15915 11152 15916 11192
rect 15956 11152 15957 11192
rect 15915 11143 15957 11152
rect 15915 11024 15957 11033
rect 15915 10984 15916 11024
rect 15956 10984 15957 11024
rect 15915 10975 15957 10984
rect 15916 10890 15956 10975
rect 16012 10949 16052 12235
rect 16108 11360 16148 13075
rect 16204 13074 16244 13159
rect 16300 12713 16340 13747
rect 16396 13301 16436 13924
rect 16395 13292 16437 13301
rect 16395 13252 16396 13292
rect 16436 13252 16437 13292
rect 16395 13243 16437 13252
rect 16492 13217 16532 16360
rect 16587 16232 16629 16241
rect 16587 16192 16588 16232
rect 16628 16192 16629 16232
rect 16587 16183 16629 16192
rect 16588 15569 16628 16183
rect 16683 15896 16725 15905
rect 16683 15856 16684 15896
rect 16724 15856 16725 15896
rect 16683 15847 16725 15856
rect 16587 15560 16629 15569
rect 16587 15520 16588 15560
rect 16628 15520 16629 15560
rect 16587 15511 16629 15520
rect 16587 14300 16629 14309
rect 16587 14260 16588 14300
rect 16628 14260 16629 14300
rect 16587 14251 16629 14260
rect 16491 13208 16533 13217
rect 16491 13168 16492 13208
rect 16532 13168 16533 13208
rect 16491 13159 16533 13168
rect 16588 13208 16628 14251
rect 16588 13159 16628 13168
rect 16492 13074 16532 13159
rect 16299 12704 16341 12713
rect 16299 12664 16300 12704
rect 16340 12664 16341 12704
rect 16299 12655 16341 12664
rect 16587 12620 16629 12629
rect 16492 12580 16588 12620
rect 16628 12580 16629 12620
rect 16492 12536 16532 12580
rect 16587 12571 16629 12580
rect 16492 12487 16532 12496
rect 16395 12452 16437 12461
rect 16395 12412 16396 12452
rect 16436 12412 16437 12452
rect 16395 12403 16437 12412
rect 16588 12452 16628 12461
rect 16108 11320 16244 11360
rect 16204 11024 16244 11320
rect 16011 10940 16053 10949
rect 16011 10900 16012 10940
rect 16052 10900 16053 10940
rect 16011 10891 16053 10900
rect 16107 10268 16149 10277
rect 16107 10228 16108 10268
rect 16148 10228 16149 10268
rect 16107 10219 16149 10228
rect 16011 8672 16053 8681
rect 16011 8632 16012 8672
rect 16052 8632 16053 8672
rect 16011 8623 16053 8632
rect 15916 7253 15956 7284
rect 15915 7244 15957 7253
rect 15915 7204 15916 7244
rect 15956 7204 15957 7244
rect 15915 7195 15957 7204
rect 16012 7244 16052 8623
rect 16012 7195 16052 7204
rect 15724 6868 15860 6908
rect 15916 7160 15956 7195
rect 15531 6740 15573 6749
rect 15531 6700 15532 6740
rect 15572 6700 15573 6740
rect 15531 6691 15573 6700
rect 15052 5816 15092 6448
rect 15052 5144 15092 5776
rect 14763 5060 14805 5069
rect 14763 5020 14764 5060
rect 14804 5020 14805 5060
rect 14763 5011 14805 5020
rect 15052 4304 15092 5104
rect 15531 5060 15573 5069
rect 15531 5020 15532 5060
rect 15572 5020 15573 5060
rect 15531 5011 15573 5020
rect 15052 3632 15092 4264
rect 15148 3641 15188 3660
rect 15147 3632 15189 3641
rect 15092 3592 15148 3632
rect 15188 3592 15189 3632
rect 15052 2792 15092 3592
rect 15147 3583 15189 3592
rect 15052 2743 15092 2752
rect 14379 2708 14421 2717
rect 14379 2668 14380 2708
rect 14420 2668 14421 2708
rect 14379 2659 14421 2668
rect 14380 2574 14420 2659
rect 13996 2456 14036 2465
rect 13899 2120 13941 2129
rect 13899 2080 13900 2120
rect 13940 2080 13941 2120
rect 13899 2071 13941 2080
rect 13900 1986 13940 2071
rect 13324 1819 13364 1828
rect 12747 1700 12789 1709
rect 12747 1660 12748 1700
rect 12788 1660 12789 1700
rect 12747 1651 12789 1660
rect 12940 1700 12980 1709
rect 12651 776 12693 785
rect 12651 736 12652 776
rect 12692 736 12693 776
rect 12651 727 12693 736
rect 12748 80 12788 1651
rect 12940 869 12980 1660
rect 13132 1700 13172 1709
rect 13132 1457 13172 1660
rect 13899 1532 13941 1541
rect 13899 1492 13900 1532
rect 13940 1492 13941 1532
rect 13899 1483 13941 1492
rect 13131 1448 13173 1457
rect 13131 1408 13132 1448
rect 13172 1408 13173 1448
rect 13131 1399 13173 1408
rect 13707 1280 13749 1289
rect 13707 1240 13708 1280
rect 13748 1240 13749 1280
rect 13707 1231 13749 1240
rect 13035 1196 13077 1205
rect 13035 1156 13036 1196
rect 13076 1156 13077 1196
rect 13035 1147 13077 1156
rect 13419 1196 13461 1205
rect 13419 1156 13420 1196
rect 13460 1156 13461 1196
rect 13419 1147 13461 1156
rect 13036 1062 13076 1147
rect 13420 1062 13460 1147
rect 13228 944 13268 953
rect 13611 944 13653 953
rect 13268 904 13556 944
rect 13228 895 13268 904
rect 12939 860 12981 869
rect 12939 820 12940 860
rect 12980 820 12981 860
rect 12939 811 12981 820
rect 12939 524 12981 533
rect 12939 484 12940 524
rect 12980 484 12981 524
rect 12939 475 12981 484
rect 12940 80 12980 475
rect 13323 440 13365 449
rect 13323 400 13324 440
rect 13364 400 13365 440
rect 13323 391 13365 400
rect 13131 356 13173 365
rect 13131 316 13132 356
rect 13172 316 13173 356
rect 13131 307 13173 316
rect 13132 80 13172 307
rect 13324 80 13364 391
rect 13516 80 13556 904
rect 13611 904 13612 944
rect 13652 904 13653 944
rect 13611 895 13653 904
rect 13612 810 13652 895
rect 13708 80 13748 1231
rect 13803 1196 13845 1205
rect 13803 1156 13804 1196
rect 13844 1156 13845 1196
rect 13803 1147 13845 1156
rect 13804 1062 13844 1147
rect 13900 80 13940 1483
rect 13996 776 14036 2416
rect 14283 2456 14325 2465
rect 14283 2416 14284 2456
rect 14324 2416 14325 2456
rect 14283 2407 14325 2416
rect 14571 2456 14613 2465
rect 14571 2416 14572 2456
rect 14612 2416 14613 2456
rect 14571 2407 14613 2416
rect 15147 2456 15189 2465
rect 15147 2416 15148 2456
rect 15188 2416 15189 2456
rect 15147 2407 15189 2416
rect 14572 2322 14612 2407
rect 14571 2120 14613 2129
rect 14571 2080 14572 2120
rect 14612 2080 14613 2120
rect 14571 2071 14613 2080
rect 14283 1868 14325 1877
rect 14283 1828 14284 1868
rect 14324 1828 14325 1868
rect 14283 1819 14325 1828
rect 14092 1700 14132 1709
rect 14092 1037 14132 1660
rect 14188 1280 14228 1289
rect 14284 1280 14324 1819
rect 14475 1700 14517 1709
rect 14475 1660 14476 1700
rect 14516 1660 14517 1700
rect 14475 1651 14517 1660
rect 14476 1566 14516 1651
rect 14475 1364 14517 1373
rect 14475 1324 14476 1364
rect 14516 1324 14517 1364
rect 14475 1315 14517 1324
rect 14228 1240 14324 1280
rect 14188 1231 14228 1240
rect 14091 1028 14133 1037
rect 14091 988 14092 1028
rect 14132 988 14133 1028
rect 14091 979 14133 988
rect 14283 944 14325 953
rect 14283 904 14284 944
rect 14324 904 14325 944
rect 14283 895 14325 904
rect 14380 944 14420 953
rect 13996 736 14132 776
rect 14092 80 14132 736
rect 14284 80 14324 895
rect 14380 365 14420 904
rect 14379 356 14421 365
rect 14379 316 14380 356
rect 14420 316 14421 356
rect 14379 307 14421 316
rect 14476 80 14516 1315
rect 14572 1196 14612 2071
rect 14667 1868 14709 1877
rect 14667 1828 14668 1868
rect 14708 1828 14709 1868
rect 15148 1868 15188 2407
rect 15243 2120 15285 2129
rect 15243 2080 15244 2120
rect 15284 2080 15380 2120
rect 15243 2071 15285 2080
rect 15244 1986 15284 2071
rect 15148 1828 15284 1868
rect 14667 1819 14709 1828
rect 14668 1734 14708 1819
rect 14859 1700 14901 1709
rect 14859 1660 14860 1700
rect 14900 1660 14901 1700
rect 14859 1651 14901 1660
rect 14572 1147 14612 1156
rect 14667 944 14709 953
rect 14667 904 14668 944
rect 14708 904 14709 944
rect 14667 895 14709 904
rect 14764 944 14804 953
rect 14668 80 14708 895
rect 14764 533 14804 904
rect 14763 524 14805 533
rect 14763 484 14764 524
rect 14804 484 14805 524
rect 14763 475 14805 484
rect 14860 80 14900 1651
rect 14955 1196 14997 1205
rect 14955 1156 14956 1196
rect 14996 1156 14997 1196
rect 14955 1147 14997 1156
rect 14956 1062 14996 1147
rect 15148 944 15188 953
rect 15051 860 15093 869
rect 15051 820 15052 860
rect 15092 820 15093 860
rect 15051 811 15093 820
rect 15052 80 15092 811
rect 15148 449 15188 904
rect 15147 440 15189 449
rect 15147 400 15148 440
rect 15188 400 15189 440
rect 15147 391 15189 400
rect 15244 80 15284 1828
rect 15340 1196 15380 2080
rect 15435 1784 15477 1793
rect 15435 1744 15436 1784
rect 15476 1744 15477 1784
rect 15435 1735 15477 1744
rect 15436 1650 15476 1735
rect 15435 1448 15477 1457
rect 15435 1408 15436 1448
rect 15476 1408 15477 1448
rect 15435 1399 15477 1408
rect 15340 1147 15380 1156
rect 15436 80 15476 1399
rect 15532 1373 15572 5011
rect 15627 1868 15669 1877
rect 15627 1828 15628 1868
rect 15668 1828 15669 1868
rect 15627 1819 15669 1828
rect 15628 1734 15668 1819
rect 15531 1364 15573 1373
rect 15531 1324 15532 1364
rect 15572 1324 15573 1364
rect 15531 1315 15573 1324
rect 15627 1280 15669 1289
rect 15627 1240 15628 1280
rect 15668 1240 15669 1280
rect 15627 1231 15669 1240
rect 15532 944 15572 953
rect 15532 701 15572 904
rect 15531 692 15573 701
rect 15531 652 15532 692
rect 15572 652 15573 692
rect 15531 643 15573 652
rect 15628 80 15668 1231
rect 15724 1196 15764 6868
rect 15819 6740 15861 6749
rect 15819 6700 15820 6740
rect 15860 6700 15861 6740
rect 15819 6691 15861 6700
rect 15820 1877 15860 6691
rect 15916 4145 15956 7120
rect 15915 4136 15957 4145
rect 15915 4096 15916 4136
rect 15956 4096 15957 4136
rect 15915 4087 15957 4096
rect 15915 3212 15957 3221
rect 15915 3172 15916 3212
rect 15956 3172 15957 3212
rect 15915 3163 15957 3172
rect 15819 1868 15861 1877
rect 15819 1828 15820 1868
rect 15860 1828 15861 1868
rect 15819 1819 15861 1828
rect 15820 1700 15860 1709
rect 15820 1541 15860 1660
rect 15819 1532 15861 1541
rect 15819 1492 15820 1532
rect 15860 1492 15861 1532
rect 15819 1483 15861 1492
rect 15819 1364 15861 1373
rect 15819 1324 15820 1364
rect 15860 1324 15861 1364
rect 15819 1315 15861 1324
rect 15724 1147 15764 1156
rect 15820 80 15860 1315
rect 15916 1280 15956 3163
rect 16011 1868 16053 1877
rect 16011 1828 16012 1868
rect 16052 1828 16053 1868
rect 16011 1819 16053 1828
rect 16012 1734 16052 1819
rect 16108 1364 16148 10219
rect 16204 10193 16244 10984
rect 16300 11024 16340 11035
rect 16300 10949 16340 10984
rect 16299 10940 16341 10949
rect 16299 10900 16300 10940
rect 16340 10900 16341 10940
rect 16299 10891 16341 10900
rect 16203 10184 16245 10193
rect 16203 10144 16204 10184
rect 16244 10144 16245 10184
rect 16203 10135 16245 10144
rect 16396 9605 16436 12403
rect 16588 12377 16628 12412
rect 16587 12368 16629 12377
rect 16587 12328 16588 12368
rect 16628 12328 16629 12368
rect 16587 12319 16629 12328
rect 16491 12284 16533 12293
rect 16491 12244 16492 12284
rect 16532 12244 16533 12284
rect 16491 12235 16533 12244
rect 16395 9596 16437 9605
rect 16395 9556 16396 9596
rect 16436 9556 16437 9596
rect 16395 9547 16437 9556
rect 16492 7337 16532 12235
rect 16588 11453 16628 12319
rect 16587 11444 16629 11453
rect 16587 11404 16588 11444
rect 16628 11404 16629 11444
rect 16587 11395 16629 11404
rect 16587 11276 16629 11285
rect 16587 11236 16588 11276
rect 16628 11236 16629 11276
rect 16587 11227 16629 11236
rect 16588 10856 16628 11227
rect 16588 10807 16628 10816
rect 16684 9857 16724 15847
rect 16780 15728 16820 16360
rect 16875 16232 16917 16241
rect 17068 16232 17108 18712
rect 17164 18584 17204 18593
rect 17164 18425 17204 18544
rect 17260 18584 17300 19048
rect 17260 18535 17300 18544
rect 17452 18542 17492 18551
rect 17452 18500 17492 18502
rect 17452 18460 17499 18500
rect 17163 18416 17205 18425
rect 17459 18416 17499 18460
rect 17163 18376 17164 18416
rect 17204 18376 17205 18416
rect 17163 18367 17205 18376
rect 17260 18376 17499 18416
rect 17260 18173 17300 18376
rect 17259 18164 17301 18173
rect 17259 18124 17260 18164
rect 17300 18124 17301 18164
rect 17259 18115 17301 18124
rect 17163 17996 17205 18005
rect 17163 17956 17164 17996
rect 17204 17956 17205 17996
rect 17163 17947 17205 17956
rect 17164 17862 17204 17947
rect 17259 17912 17301 17921
rect 17259 17872 17260 17912
rect 17300 17872 17301 17912
rect 17259 17863 17301 17872
rect 17451 17912 17493 17921
rect 17451 17872 17452 17912
rect 17492 17872 17493 17912
rect 17451 17863 17493 17872
rect 17163 17324 17205 17333
rect 17163 17284 17164 17324
rect 17204 17284 17205 17324
rect 17163 17275 17205 17284
rect 17164 17240 17204 17275
rect 17164 17189 17204 17200
rect 17260 16484 17300 17863
rect 17355 17828 17397 17837
rect 17355 17788 17356 17828
rect 17396 17788 17397 17828
rect 17355 17779 17397 17788
rect 17356 17744 17396 17779
rect 17356 17693 17396 17704
rect 17260 16444 17396 16484
rect 17259 16316 17301 16325
rect 17259 16276 17260 16316
rect 17300 16276 17301 16316
rect 17259 16267 17301 16276
rect 16875 16192 16876 16232
rect 16916 16192 16917 16232
rect 16875 16183 16917 16192
rect 16972 16192 17108 16232
rect 16876 16098 16916 16183
rect 16972 15905 17012 16192
rect 17260 16182 17300 16267
rect 17068 16064 17108 16073
rect 16971 15896 17013 15905
rect 16971 15856 16972 15896
rect 17012 15856 17013 15896
rect 16971 15847 17013 15856
rect 16971 15728 17013 15737
rect 16780 15688 16916 15728
rect 16779 15560 16821 15569
rect 16779 15520 16780 15560
rect 16820 15520 16821 15560
rect 16779 15511 16821 15520
rect 16780 15426 16820 15511
rect 16779 14888 16821 14897
rect 16779 14848 16780 14888
rect 16820 14848 16821 14888
rect 16779 14839 16821 14848
rect 16780 14729 16820 14839
rect 16779 14720 16821 14729
rect 16779 14680 16780 14720
rect 16820 14680 16821 14720
rect 16779 14671 16821 14680
rect 16780 14586 16820 14671
rect 16876 14048 16916 15688
rect 16971 15688 16972 15728
rect 17012 15688 17013 15728
rect 16971 15679 17013 15688
rect 16972 15594 17012 15679
rect 16780 14008 16876 14048
rect 16780 12461 16820 14008
rect 16876 13999 16916 14008
rect 16972 14720 17012 14729
rect 16876 13460 16916 13469
rect 16972 13460 17012 14680
rect 17068 14720 17108 16024
rect 17164 15560 17204 15569
rect 17164 14972 17204 15520
rect 17260 15560 17300 15569
rect 17260 15149 17300 15520
rect 17259 15140 17301 15149
rect 17259 15100 17260 15140
rect 17300 15100 17301 15140
rect 17259 15091 17301 15100
rect 17260 14972 17300 14981
rect 17164 14932 17260 14972
rect 17260 14923 17300 14932
rect 17356 14897 17396 16444
rect 17452 16400 17492 17863
rect 17548 17333 17588 19207
rect 17737 19172 17777 19300
rect 17836 19256 17876 19265
rect 17737 19132 17780 19172
rect 17643 19088 17685 19097
rect 17643 19048 17644 19088
rect 17684 19048 17685 19088
rect 17643 19039 17685 19048
rect 17644 18954 17684 19039
rect 17547 17324 17589 17333
rect 17547 17284 17548 17324
rect 17588 17284 17589 17324
rect 17547 17275 17589 17284
rect 17643 17072 17685 17081
rect 17643 17032 17644 17072
rect 17684 17032 17685 17072
rect 17643 17023 17685 17032
rect 17644 16938 17684 17023
rect 17452 16351 17492 16360
rect 17643 16316 17685 16325
rect 17643 16276 17644 16316
rect 17684 16276 17685 16316
rect 17643 16267 17685 16276
rect 17644 16182 17684 16267
rect 17643 15812 17685 15821
rect 17643 15772 17644 15812
rect 17684 15772 17685 15812
rect 17643 15763 17685 15772
rect 17547 15728 17589 15737
rect 17547 15688 17548 15728
rect 17588 15688 17589 15728
rect 17547 15679 17589 15688
rect 17452 15569 17492 15654
rect 17451 15560 17493 15569
rect 17451 15520 17452 15560
rect 17492 15520 17493 15560
rect 17451 15511 17493 15520
rect 17451 15308 17493 15317
rect 17451 15268 17452 15308
rect 17492 15268 17493 15308
rect 17451 15259 17493 15268
rect 17452 15174 17492 15259
rect 17355 14888 17397 14897
rect 17355 14848 17356 14888
rect 17396 14848 17397 14888
rect 17355 14839 17397 14848
rect 17260 14720 17300 14729
rect 17452 14720 17492 14729
rect 17108 14680 17204 14720
rect 17068 14671 17108 14680
rect 17067 14552 17109 14561
rect 17067 14512 17068 14552
rect 17108 14512 17109 14552
rect 17164 14552 17204 14680
rect 17300 14680 17452 14720
rect 17260 14671 17300 14680
rect 17452 14671 17492 14680
rect 17548 14720 17588 15679
rect 17644 15560 17684 15763
rect 17740 15560 17780 19132
rect 17836 19097 17876 19216
rect 17835 19088 17877 19097
rect 17835 19048 17836 19088
rect 17876 19048 17877 19088
rect 17835 19039 17877 19048
rect 17835 17576 17877 17585
rect 17835 17536 17836 17576
rect 17876 17536 17877 17576
rect 17835 17527 17877 17536
rect 17836 16400 17876 17527
rect 17836 16351 17876 16360
rect 17932 15905 17972 19543
rect 18028 17669 18068 20560
rect 18124 19769 18164 20728
rect 18220 20768 18260 20777
rect 18220 20021 18260 20728
rect 18219 20012 18261 20021
rect 18219 19972 18220 20012
rect 18260 19972 18261 20012
rect 18219 19963 18261 19972
rect 18123 19760 18165 19769
rect 18123 19720 18124 19760
rect 18164 19720 18165 19760
rect 18123 19711 18165 19720
rect 18123 19508 18165 19517
rect 18123 19468 18124 19508
rect 18164 19468 18165 19508
rect 18123 19459 18165 19468
rect 18027 17660 18069 17669
rect 18027 17620 18028 17660
rect 18068 17620 18069 17660
rect 18027 17611 18069 17620
rect 18124 16745 18164 19459
rect 18219 18080 18261 18089
rect 18219 18040 18220 18080
rect 18260 18040 18261 18080
rect 18219 18031 18261 18040
rect 18123 16736 18165 16745
rect 18123 16696 18124 16736
rect 18164 16696 18165 16736
rect 18123 16687 18165 16696
rect 18220 16661 18260 18031
rect 18219 16652 18261 16661
rect 18219 16612 18220 16652
rect 18260 16612 18261 16652
rect 18219 16603 18261 16612
rect 18028 16232 18068 16241
rect 17931 15896 17973 15905
rect 17931 15856 17932 15896
rect 17972 15856 17973 15896
rect 17931 15847 17973 15856
rect 17740 15520 17876 15560
rect 17644 15511 17684 15520
rect 17739 15392 17781 15401
rect 17739 15352 17740 15392
rect 17780 15352 17781 15392
rect 17739 15343 17781 15352
rect 17643 15308 17685 15317
rect 17643 15268 17644 15308
rect 17684 15268 17685 15308
rect 17643 15259 17685 15268
rect 17548 14671 17588 14680
rect 17547 14552 17589 14561
rect 17644 14552 17684 15259
rect 17740 15233 17780 15343
rect 17739 15224 17781 15233
rect 17739 15184 17740 15224
rect 17780 15184 17781 15224
rect 17739 15175 17781 15184
rect 17740 14720 17780 15175
rect 17836 15065 17876 15520
rect 17931 15140 17973 15149
rect 17931 15100 17932 15140
rect 17972 15100 17973 15140
rect 17931 15091 17973 15100
rect 17835 15056 17877 15065
rect 17835 15016 17836 15056
rect 17876 15016 17877 15056
rect 17835 15007 17877 15016
rect 17740 14671 17780 14680
rect 17164 14512 17396 14552
rect 17067 14503 17109 14512
rect 16916 13420 17012 13460
rect 16876 13411 16916 13420
rect 17068 13292 17108 14503
rect 17163 14384 17205 14393
rect 17163 14344 17164 14384
rect 17204 14344 17205 14384
rect 17163 14335 17205 14344
rect 16876 13252 17108 13292
rect 16779 12452 16821 12461
rect 16779 12412 16780 12452
rect 16820 12412 16821 12452
rect 16779 12403 16821 12412
rect 16779 12032 16821 12041
rect 16876 12032 16916 13252
rect 16971 12704 17013 12713
rect 16971 12664 16972 12704
rect 17012 12664 17013 12704
rect 16971 12655 17013 12664
rect 16972 12536 17012 12655
rect 16972 12487 17012 12496
rect 17068 12536 17108 12545
rect 17068 12461 17108 12496
rect 17067 12452 17109 12461
rect 17067 12412 17068 12452
rect 17108 12412 17109 12452
rect 17067 12403 17109 12412
rect 16779 11992 16780 12032
rect 16820 11992 16916 12032
rect 16779 11983 16821 11992
rect 16780 11024 16820 11983
rect 16971 11696 17013 11705
rect 16971 11656 16972 11696
rect 17012 11656 17013 11696
rect 16971 11647 17013 11656
rect 16972 11562 17012 11647
rect 17068 11621 17108 12403
rect 17164 12293 17204 14335
rect 17356 14057 17396 14512
rect 17547 14512 17548 14552
rect 17588 14512 17684 14552
rect 17547 14503 17589 14512
rect 17547 14384 17589 14393
rect 17547 14344 17548 14384
rect 17588 14344 17589 14384
rect 17547 14335 17589 14344
rect 17451 14300 17493 14309
rect 17451 14260 17452 14300
rect 17492 14260 17493 14300
rect 17451 14251 17493 14260
rect 17355 14048 17397 14057
rect 17355 14003 17356 14048
rect 17396 14003 17397 14048
rect 17355 13999 17397 14003
rect 17356 13914 17396 13999
rect 17259 13208 17301 13217
rect 17259 13168 17260 13208
rect 17300 13168 17301 13208
rect 17259 13159 17301 13168
rect 17356 13208 17396 13217
rect 17452 13208 17492 14251
rect 17548 14216 17588 14335
rect 17836 14309 17876 15007
rect 17835 14300 17877 14309
rect 17835 14260 17836 14300
rect 17876 14260 17877 14300
rect 17835 14251 17877 14260
rect 17932 14216 17972 15091
rect 18028 14393 18068 16192
rect 18220 16232 18260 16241
rect 18124 16064 18164 16073
rect 18124 15569 18164 16024
rect 18220 15737 18260 16192
rect 18219 15728 18261 15737
rect 18219 15688 18220 15728
rect 18260 15688 18261 15728
rect 18219 15679 18261 15688
rect 18123 15560 18165 15569
rect 18123 15520 18124 15560
rect 18164 15520 18165 15560
rect 18123 15511 18165 15520
rect 18316 15392 18356 23752
rect 18412 22709 18452 25171
rect 18603 24884 18645 24893
rect 18603 24844 18604 24884
rect 18644 24844 18645 24884
rect 18603 24835 18645 24844
rect 18604 24632 18644 24835
rect 18508 24613 18548 24622
rect 18604 24583 18644 24592
rect 18508 23129 18548 24573
rect 18603 23960 18645 23969
rect 18603 23920 18604 23960
rect 18644 23920 18645 23960
rect 18603 23911 18645 23920
rect 18507 23120 18549 23129
rect 18507 23080 18508 23120
rect 18548 23080 18549 23120
rect 18604 23120 18644 23911
rect 18700 23372 18740 25852
rect 19179 25843 19221 25852
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 19083 25556 19125 25565
rect 19083 25516 19084 25556
rect 19124 25516 19125 25556
rect 19083 25507 19125 25516
rect 19084 25422 19124 25507
rect 19179 25472 19221 25481
rect 19179 25432 19180 25472
rect 19220 25432 19221 25472
rect 19179 25423 19221 25432
rect 18892 25304 18932 25315
rect 18892 25229 18932 25264
rect 18891 25220 18933 25229
rect 18891 25180 18892 25220
rect 18932 25180 18933 25220
rect 18891 25171 18933 25180
rect 19180 24716 19220 25423
rect 19372 25304 19412 25852
rect 19468 25481 19508 26356
rect 19660 26272 19988 26312
rect 19563 25892 19605 25901
rect 19563 25852 19564 25892
rect 19604 25852 19605 25892
rect 19563 25843 19605 25852
rect 19564 25758 19604 25843
rect 19660 25640 19700 26272
rect 19755 26144 19797 26153
rect 19755 26104 19756 26144
rect 19796 26104 19797 26144
rect 19755 26095 19797 26104
rect 19852 26144 19892 26153
rect 19756 26010 19796 26095
rect 19564 25600 19700 25640
rect 19467 25472 19509 25481
rect 19467 25432 19468 25472
rect 19508 25432 19509 25472
rect 19467 25423 19509 25432
rect 19276 25283 19316 25292
rect 19564 25304 19604 25600
rect 19852 25481 19892 26104
rect 19948 26144 19988 26272
rect 19948 26095 19988 26104
rect 20044 26144 20084 26153
rect 19659 25472 19701 25481
rect 19659 25432 19660 25472
rect 19700 25432 19701 25472
rect 19659 25423 19701 25432
rect 19851 25472 19893 25481
rect 19851 25432 19852 25472
rect 19892 25432 19893 25472
rect 19851 25423 19893 25432
rect 19372 25255 19412 25264
rect 19468 25283 19508 25292
rect 19276 24893 19316 25243
rect 19564 25255 19604 25264
rect 19468 25145 19508 25243
rect 19467 25136 19509 25145
rect 19467 25096 19468 25136
rect 19508 25096 19509 25136
rect 19660 25136 19700 25423
rect 19755 25388 19797 25397
rect 20044 25388 20084 26104
rect 19755 25348 19756 25388
rect 19796 25348 19797 25388
rect 19755 25339 19797 25348
rect 19948 25348 20084 25388
rect 19756 25304 19796 25339
rect 19756 25253 19796 25264
rect 19852 25304 19892 25313
rect 19660 25096 19796 25136
rect 19467 25087 19509 25096
rect 19275 24884 19317 24893
rect 19275 24844 19276 24884
rect 19316 24844 19317 24884
rect 19275 24835 19317 24844
rect 19371 24800 19413 24809
rect 19371 24760 19372 24800
rect 19412 24760 19413 24800
rect 19371 24751 19413 24760
rect 19659 24800 19701 24809
rect 19659 24760 19660 24800
rect 19700 24760 19701 24800
rect 19659 24751 19701 24760
rect 19180 24676 19316 24716
rect 18987 24632 19029 24641
rect 18987 24592 18988 24632
rect 19028 24592 19029 24632
rect 18987 24583 19029 24592
rect 18988 24389 19028 24583
rect 19083 24548 19125 24557
rect 19083 24508 19084 24548
rect 19124 24508 19125 24548
rect 19083 24499 19125 24508
rect 19084 24414 19124 24499
rect 18987 24380 19029 24389
rect 18987 24340 18988 24380
rect 19028 24340 19029 24380
rect 18987 24331 19029 24340
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 19276 23801 19316 24676
rect 19275 23792 19317 23801
rect 19275 23752 19276 23792
rect 19316 23752 19317 23792
rect 19275 23743 19317 23752
rect 18700 23332 18836 23372
rect 18796 23288 18836 23332
rect 18892 23288 18932 23297
rect 18796 23248 18892 23288
rect 18892 23239 18932 23248
rect 19120 23288 19162 23297
rect 19120 23248 19121 23288
rect 19161 23248 19162 23288
rect 19372 23288 19412 24751
rect 19564 24632 19604 24641
rect 19564 24305 19604 24592
rect 19563 24296 19605 24305
rect 19563 24256 19564 24296
rect 19604 24256 19605 24296
rect 19563 24247 19605 24256
rect 19660 23969 19700 24751
rect 19659 23960 19701 23969
rect 19659 23920 19660 23960
rect 19700 23920 19701 23960
rect 19659 23911 19701 23920
rect 19563 23792 19605 23801
rect 19563 23752 19564 23792
rect 19604 23752 19605 23792
rect 19563 23743 19605 23752
rect 19564 23658 19604 23743
rect 19756 23624 19796 25096
rect 19852 24893 19892 25264
rect 19851 24884 19893 24893
rect 19851 24844 19852 24884
rect 19892 24844 19893 24884
rect 19851 24835 19893 24844
rect 19948 24716 19988 25348
rect 20044 25145 20084 25230
rect 20043 25136 20085 25145
rect 20043 25096 20044 25136
rect 20084 25096 20085 25136
rect 20043 25087 20085 25096
rect 20524 24977 20564 26515
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 20523 24968 20565 24977
rect 20523 24928 20524 24968
rect 20564 24928 20565 24968
rect 20523 24919 20565 24928
rect 20043 24800 20085 24809
rect 20043 24760 20044 24800
rect 20084 24760 20085 24800
rect 20043 24751 20085 24760
rect 19756 23575 19796 23584
rect 19852 24676 19988 24716
rect 19852 23297 19892 24676
rect 20044 24618 20084 24751
rect 20044 24473 20084 24578
rect 20236 24716 20276 24725
rect 20043 24464 20085 24473
rect 20043 24424 20044 24464
rect 20084 24424 20085 24464
rect 20043 24415 20085 24424
rect 20236 23960 20276 24676
rect 20523 24464 20565 24473
rect 20523 24424 20524 24464
rect 20564 24424 20565 24464
rect 20523 24415 20565 24424
rect 19948 23920 20276 23960
rect 19948 23792 19988 23920
rect 19948 23743 19988 23752
rect 20044 23792 20084 23801
rect 20044 23624 20084 23752
rect 19948 23584 20084 23624
rect 19851 23288 19893 23297
rect 19372 23248 19508 23288
rect 19120 23239 19162 23248
rect 18700 23120 18740 23129
rect 18604 23080 18700 23120
rect 18507 23071 18549 23080
rect 18411 22700 18453 22709
rect 18411 22660 18412 22700
rect 18452 22660 18453 22700
rect 18411 22651 18453 22660
rect 18700 22532 18740 23080
rect 19121 23120 19161 23239
rect 19121 23071 19161 23080
rect 19276 23120 19316 23129
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 18700 22492 18932 22532
rect 18604 22280 18644 22289
rect 18412 22112 18452 22121
rect 18604 22112 18644 22240
rect 18452 22072 18644 22112
rect 18412 22063 18452 22072
rect 18412 20768 18452 20777
rect 18412 19937 18452 20728
rect 18508 20768 18548 20777
rect 18508 20189 18548 20728
rect 18604 20609 18644 22072
rect 18699 21692 18741 21701
rect 18699 21652 18700 21692
rect 18740 21652 18741 21692
rect 18699 21643 18741 21652
rect 18603 20600 18645 20609
rect 18603 20560 18604 20600
rect 18644 20560 18645 20600
rect 18603 20551 18645 20560
rect 18700 20264 18740 21643
rect 18892 21608 18932 22492
rect 19276 21944 19316 23080
rect 19084 21904 19316 21944
rect 19372 23120 19412 23129
rect 19084 21776 19124 21904
rect 19084 21727 19124 21736
rect 19180 21617 19220 21904
rect 19276 21776 19316 21785
rect 19372 21776 19412 23080
rect 19316 21736 19412 21776
rect 19276 21727 19316 21736
rect 18892 21440 18932 21568
rect 19179 21608 19221 21617
rect 19179 21568 19180 21608
rect 19220 21568 19221 21608
rect 19179 21559 19221 21568
rect 19468 21608 19508 23248
rect 19851 23248 19852 23288
rect 19892 23248 19893 23288
rect 19851 23239 19893 23248
rect 19564 23120 19604 23129
rect 19564 21785 19604 23080
rect 19660 23120 19700 23129
rect 19851 23120 19893 23129
rect 19700 23080 19796 23120
rect 19660 23071 19700 23080
rect 19659 22868 19701 22877
rect 19659 22828 19660 22868
rect 19700 22828 19701 22868
rect 19659 22819 19701 22828
rect 19660 22734 19700 22819
rect 19563 21776 19605 21785
rect 19563 21736 19564 21776
rect 19604 21736 19605 21776
rect 19563 21727 19605 21736
rect 18892 21400 19316 21440
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 19276 21020 19316 21400
rect 19084 20980 19316 21020
rect 18796 20768 18836 20777
rect 18796 20441 18836 20728
rect 18795 20432 18837 20441
rect 18795 20392 18796 20432
rect 18836 20392 18837 20432
rect 18795 20383 18837 20392
rect 18892 20264 18932 20273
rect 18700 20224 18892 20264
rect 18892 20215 18932 20224
rect 18507 20180 18549 20189
rect 18507 20140 18508 20180
rect 18548 20140 18549 20180
rect 18507 20131 18549 20140
rect 18700 20096 18740 20105
rect 19084 20096 19124 20980
rect 19468 20945 19508 21568
rect 19563 21608 19605 21617
rect 19563 21568 19564 21608
rect 19604 21568 19605 21608
rect 19563 21559 19605 21568
rect 19564 21474 19604 21559
rect 19756 21440 19796 23080
rect 19851 23080 19852 23120
rect 19892 23080 19893 23120
rect 19851 23071 19893 23080
rect 19948 23120 19988 23584
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 20139 23288 20181 23297
rect 20139 23248 20140 23288
rect 20180 23248 20181 23288
rect 20139 23239 20181 23248
rect 20140 23154 20180 23239
rect 19988 23080 20084 23120
rect 19948 23071 19988 23080
rect 19852 22986 19892 23071
rect 20044 22532 20084 23080
rect 20044 22483 20084 22492
rect 19851 22448 19893 22457
rect 19851 22408 19852 22448
rect 19892 22408 19893 22448
rect 19851 22399 19893 22408
rect 19852 22280 19892 22399
rect 19892 22240 19988 22280
rect 19852 22231 19892 22240
rect 19948 21776 19988 22240
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 20524 21776 20564 24415
rect 20812 24305 20852 26599
rect 20811 24296 20853 24305
rect 20811 24256 20812 24296
rect 20852 24256 20853 24296
rect 20811 24247 20853 24256
rect 21004 23960 21044 32647
rect 21388 29345 21428 38704
rect 21387 29336 21429 29345
rect 21387 29296 21388 29336
rect 21428 29296 21429 29336
rect 21387 29287 21429 29296
rect 21004 23920 21428 23960
rect 21388 22961 21428 23920
rect 21387 22952 21429 22961
rect 21387 22912 21388 22952
rect 21428 22912 21429 22952
rect 21387 22903 21429 22912
rect 20811 22616 20853 22625
rect 20811 22576 20812 22616
rect 20852 22576 20853 22616
rect 20811 22567 20853 22576
rect 20619 21944 20661 21953
rect 20619 21904 20620 21944
rect 20660 21904 20661 21944
rect 20619 21895 20661 21904
rect 19948 21736 20084 21776
rect 19851 21692 19893 21701
rect 19851 21652 19852 21692
rect 19892 21652 19893 21692
rect 19851 21643 19893 21652
rect 19852 21608 19892 21643
rect 19852 21557 19892 21568
rect 19947 21608 19989 21617
rect 19947 21568 19948 21608
rect 19988 21568 19989 21608
rect 19947 21559 19989 21568
rect 19948 21474 19988 21559
rect 19852 21440 19892 21449
rect 19756 21400 19852 21440
rect 19852 21391 19892 21400
rect 19467 20936 19509 20945
rect 19467 20896 19468 20936
rect 19508 20896 19509 20936
rect 19467 20887 19509 20896
rect 19179 20768 19221 20777
rect 20044 20768 20084 21736
rect 20236 21736 20564 21776
rect 20139 21608 20181 21617
rect 20139 21568 20140 21608
rect 20180 21568 20181 21608
rect 20139 21559 20181 21568
rect 20140 21474 20180 21559
rect 20236 21020 20276 21736
rect 20236 20971 20276 20980
rect 19179 20728 19180 20768
rect 19220 20728 19221 20768
rect 19179 20719 19221 20728
rect 19948 20728 20044 20768
rect 19180 20264 19220 20719
rect 19948 20357 19988 20728
rect 20044 20719 20084 20728
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 19947 20348 19989 20357
rect 19947 20308 19948 20348
rect 19988 20308 19989 20348
rect 19947 20299 19989 20308
rect 19180 20224 19508 20264
rect 19180 20180 19220 20224
rect 18604 20056 18700 20096
rect 18740 20056 19124 20096
rect 19175 20140 19220 20180
rect 19175 20096 19215 20140
rect 18411 19928 18453 19937
rect 18411 19888 18412 19928
rect 18452 19888 18453 19928
rect 18411 19879 18453 19888
rect 18604 19181 18644 20056
rect 18700 20047 18740 20056
rect 19175 20047 19215 20056
rect 19276 20096 19316 20105
rect 18808 19676 19176 19685
rect 19276 19676 19316 20056
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 19228 19636 19316 19676
rect 19372 20096 19412 20105
rect 19228 19592 19268 19636
rect 19200 19552 19268 19592
rect 19200 19508 19240 19552
rect 19180 19468 19240 19508
rect 19084 19256 19124 19265
rect 18988 19216 19084 19256
rect 18603 19172 18645 19181
rect 18603 19132 18604 19172
rect 18644 19132 18645 19172
rect 18603 19123 18645 19132
rect 18604 17744 18644 19123
rect 18988 18920 19028 19216
rect 19084 19207 19124 19216
rect 19180 19088 19220 19468
rect 19275 19172 19317 19181
rect 19275 19132 19276 19172
rect 19316 19132 19317 19172
rect 19275 19123 19317 19132
rect 18411 17408 18453 17417
rect 18411 17368 18412 17408
rect 18452 17368 18453 17408
rect 18411 17359 18453 17368
rect 18124 15352 18356 15392
rect 18027 14384 18069 14393
rect 18027 14344 18028 14384
rect 18068 14344 18069 14384
rect 18027 14335 18069 14344
rect 18028 14216 18068 14225
rect 17932 14176 18028 14216
rect 17548 14167 17588 14176
rect 18028 14167 18068 14176
rect 17739 14048 17781 14057
rect 17739 14008 17740 14048
rect 17780 14008 17781 14048
rect 17739 13999 17781 14008
rect 17836 14048 17876 14057
rect 17740 13914 17780 13999
rect 17836 13889 17876 14008
rect 17835 13880 17877 13889
rect 17835 13840 17836 13880
rect 17876 13840 17877 13880
rect 17835 13831 17877 13840
rect 18124 13712 18164 15352
rect 18219 15224 18261 15233
rect 18219 15184 18220 15224
rect 18260 15184 18261 15224
rect 18219 15175 18261 15184
rect 17396 13168 17492 13208
rect 17836 13672 18164 13712
rect 17163 12284 17205 12293
rect 17163 12244 17164 12284
rect 17204 12244 17205 12284
rect 17163 12235 17205 12244
rect 17260 11705 17300 13159
rect 17356 12704 17396 13168
rect 17356 12655 17396 12664
rect 17547 12704 17589 12713
rect 17547 12664 17548 12704
rect 17588 12664 17589 12704
rect 17547 12655 17589 12664
rect 17164 11696 17204 11705
rect 17067 11612 17109 11621
rect 17067 11572 17068 11612
rect 17108 11572 17109 11612
rect 17067 11563 17109 11572
rect 17164 11360 17204 11656
rect 17259 11696 17301 11705
rect 17259 11656 17260 11696
rect 17300 11656 17301 11696
rect 17259 11647 17301 11656
rect 17356 11696 17396 11707
rect 17260 11562 17300 11647
rect 17356 11621 17396 11656
rect 17355 11612 17397 11621
rect 17355 11572 17356 11612
rect 17396 11572 17397 11612
rect 17355 11563 17397 11572
rect 16876 11320 17204 11360
rect 17452 11528 17492 11537
rect 16876 11033 16916 11320
rect 17452 11276 17492 11488
rect 17548 11360 17588 12655
rect 17644 12536 17684 12547
rect 17644 12461 17684 12496
rect 17740 12536 17780 12545
rect 17643 12452 17685 12461
rect 17643 12412 17644 12452
rect 17684 12412 17685 12452
rect 17643 12403 17685 12412
rect 17740 11369 17780 12496
rect 17739 11360 17781 11369
rect 17548 11320 17684 11360
rect 17068 11236 17492 11276
rect 16971 11192 17013 11201
rect 16971 11152 16972 11192
rect 17012 11152 17013 11192
rect 16971 11143 17013 11152
rect 16972 11058 17012 11143
rect 16780 10975 16820 10984
rect 16875 11024 16917 11033
rect 16875 10984 16876 11024
rect 16916 10984 16917 11024
rect 16875 10975 16917 10984
rect 17068 11024 17108 11236
rect 17644 11033 17684 11320
rect 17739 11320 17740 11360
rect 17780 11320 17781 11360
rect 17739 11311 17781 11320
rect 17740 11192 17780 11201
rect 17068 10975 17108 10984
rect 17260 11024 17300 11033
rect 16683 9848 16725 9857
rect 16683 9808 16684 9848
rect 16724 9808 16725 9848
rect 16683 9799 16725 9808
rect 16780 9680 16820 9689
rect 16876 9680 16916 10975
rect 17067 10856 17109 10865
rect 17067 10816 17068 10856
rect 17108 10816 17109 10856
rect 17067 10807 17109 10816
rect 16971 10268 17013 10277
rect 16971 10228 16972 10268
rect 17012 10228 17013 10268
rect 16971 10219 17013 10228
rect 16972 10184 17012 10219
rect 16972 10133 17012 10144
rect 16971 10016 17013 10025
rect 16971 9976 16972 10016
rect 17012 9976 17013 10016
rect 16971 9967 17013 9976
rect 16820 9640 16916 9680
rect 16780 9631 16820 9640
rect 16587 9512 16629 9521
rect 16587 9472 16588 9512
rect 16628 9472 16629 9512
rect 16587 9463 16629 9472
rect 16491 7328 16533 7337
rect 16491 7288 16492 7328
rect 16532 7288 16533 7328
rect 16491 7279 16533 7288
rect 16492 7160 16532 7279
rect 16492 7111 16532 7120
rect 16588 6992 16628 9463
rect 16876 8672 16916 8681
rect 16876 8504 16916 8632
rect 16972 8672 17012 9967
rect 16972 8623 17012 8632
rect 17068 8504 17108 10807
rect 17163 10688 17205 10697
rect 17163 10648 17164 10688
rect 17204 10648 17205 10688
rect 17163 10639 17205 10648
rect 17164 10436 17204 10639
rect 17260 10529 17300 10984
rect 17356 11024 17396 11033
rect 17259 10520 17301 10529
rect 17259 10480 17260 10520
rect 17300 10480 17301 10520
rect 17259 10471 17301 10480
rect 17164 10387 17204 10396
rect 17356 10184 17396 10984
rect 17452 11024 17492 11033
rect 17452 10529 17492 10984
rect 17548 11024 17588 11033
rect 17548 10865 17588 10984
rect 17643 11024 17685 11033
rect 17643 10984 17644 11024
rect 17684 10984 17685 11024
rect 17643 10975 17685 10984
rect 17547 10856 17589 10865
rect 17547 10816 17548 10856
rect 17588 10816 17589 10856
rect 17547 10807 17589 10816
rect 17451 10520 17493 10529
rect 17451 10480 17452 10520
rect 17492 10480 17493 10520
rect 17451 10471 17493 10480
rect 17260 10144 17396 10184
rect 17163 8840 17205 8849
rect 17163 8800 17164 8840
rect 17204 8800 17205 8840
rect 17163 8791 17205 8800
rect 16876 8464 17108 8504
rect 17164 8504 17204 8791
rect 17164 8455 17204 8464
rect 17260 8177 17300 10144
rect 17356 10016 17396 10025
rect 17644 10016 17684 10975
rect 17740 10865 17780 11152
rect 17739 10856 17781 10865
rect 17739 10816 17740 10856
rect 17780 10816 17781 10856
rect 17739 10807 17781 10816
rect 17739 10520 17781 10529
rect 17739 10480 17740 10520
rect 17780 10480 17781 10520
rect 17739 10471 17781 10480
rect 17740 10184 17780 10471
rect 17836 10361 17876 13672
rect 18220 13628 18260 15175
rect 18412 14048 18452 17359
rect 18604 16829 18644 17704
rect 18700 18880 19028 18920
rect 19084 19048 19220 19088
rect 18700 18584 18740 18880
rect 19084 18677 19124 19048
rect 19276 19038 19316 19123
rect 19372 18794 19412 20056
rect 19372 18745 19412 18754
rect 18892 18668 18932 18677
rect 19083 18668 19125 18677
rect 19468 18668 19508 20224
rect 20620 20180 20660 21895
rect 20812 20180 20852 22567
rect 21195 21272 21237 21281
rect 21195 21232 21196 21272
rect 21236 21232 21237 21272
rect 21195 21223 21237 21232
rect 21099 20936 21141 20945
rect 21099 20896 21100 20936
rect 21140 20896 21141 20936
rect 21099 20887 21141 20896
rect 21100 20189 21140 20887
rect 20524 20140 20660 20180
rect 20716 20140 20852 20180
rect 21099 20180 21141 20189
rect 21099 20140 21100 20180
rect 21140 20140 21141 20180
rect 19564 20096 19604 20105
rect 19564 19508 19604 20056
rect 19660 20096 19700 20105
rect 19852 20096 19892 20105
rect 19700 20056 19796 20096
rect 19660 20047 19700 20056
rect 19659 19844 19701 19853
rect 19659 19804 19660 19844
rect 19700 19804 19701 19844
rect 19659 19795 19701 19804
rect 19660 19710 19700 19795
rect 19564 19468 19632 19508
rect 19592 19424 19632 19468
rect 19756 19424 19796 20056
rect 19852 19937 19892 20056
rect 19948 20096 19988 20105
rect 19851 19928 19893 19937
rect 19851 19888 19852 19928
rect 19892 19888 19893 19928
rect 19851 19879 19893 19888
rect 19948 19769 19988 20056
rect 20043 20096 20085 20105
rect 20043 20056 20044 20096
rect 20084 20056 20085 20096
rect 20043 20047 20085 20056
rect 20140 20091 20180 20100
rect 20044 19962 20084 20047
rect 19947 19760 19989 19769
rect 20140 19760 20180 20051
rect 19947 19720 19948 19760
rect 19988 19720 19989 19760
rect 19947 19711 19989 19720
rect 20044 19720 20180 19760
rect 19592 19384 19700 19424
rect 19660 19256 19700 19384
rect 19756 19375 19796 19384
rect 19947 19340 19989 19349
rect 20044 19340 20084 19720
rect 19947 19300 19948 19340
rect 19988 19300 20084 19340
rect 19947 19291 19989 19300
rect 19660 19181 19700 19216
rect 19756 19256 19796 19265
rect 19659 19172 19701 19181
rect 19659 19132 19660 19172
rect 19700 19132 19701 19172
rect 19659 19123 19701 19132
rect 19660 19092 19700 19123
rect 19756 18677 19796 19216
rect 19948 19256 19988 19291
rect 19948 19205 19988 19216
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 20043 18752 20085 18761
rect 20043 18712 20044 18752
rect 20084 18712 20085 18752
rect 20043 18703 20085 18712
rect 20235 18752 20277 18761
rect 20235 18712 20236 18752
rect 20276 18712 20277 18752
rect 20235 18703 20277 18712
rect 18932 18628 19084 18668
rect 19124 18628 19125 18668
rect 18892 18619 18932 18628
rect 19083 18619 19125 18628
rect 19372 18628 19508 18668
rect 19755 18668 19797 18677
rect 19755 18628 19756 18668
rect 19796 18628 19797 18668
rect 18700 16997 18740 18544
rect 19084 18584 19124 18619
rect 19084 18534 19124 18544
rect 19180 18584 19220 18593
rect 19180 18425 19220 18544
rect 19179 18416 19221 18425
rect 19179 18376 19180 18416
rect 19220 18376 19221 18416
rect 19179 18367 19221 18376
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 18795 17996 18837 18005
rect 18795 17956 18796 17996
rect 18836 17956 18837 17996
rect 18795 17947 18837 17956
rect 18796 17862 18836 17947
rect 19372 17912 19412 18628
rect 19755 18619 19797 18628
rect 19564 18584 19604 18593
rect 19468 18544 19564 18584
rect 19468 18005 19508 18544
rect 19564 18535 19604 18544
rect 19660 18584 19700 18593
rect 19564 18416 19604 18425
rect 19467 17996 19509 18005
rect 19467 17956 19468 17996
rect 19508 17956 19509 17996
rect 19467 17947 19509 17956
rect 19079 17872 19412 17912
rect 18891 17744 18933 17753
rect 18891 17704 18892 17744
rect 18932 17704 18933 17744
rect 18891 17695 18933 17704
rect 19079 17744 19119 17872
rect 19079 17695 19119 17704
rect 19180 17744 19220 17753
rect 18892 17576 18932 17695
rect 19084 17576 19124 17585
rect 18892 17536 19084 17576
rect 19084 17527 19124 17536
rect 19180 17501 19220 17704
rect 19275 17744 19317 17753
rect 19275 17704 19276 17744
rect 19316 17704 19317 17744
rect 19275 17695 19317 17704
rect 19276 17610 19316 17695
rect 19372 17576 19412 17872
rect 19468 17744 19508 17947
rect 19468 17695 19508 17704
rect 19564 17744 19604 18376
rect 19564 17695 19604 17704
rect 19660 17744 19700 18544
rect 19852 18584 19892 18593
rect 19892 18544 19988 18584
rect 19852 18535 19892 18544
rect 19851 18416 19893 18425
rect 19851 18376 19852 18416
rect 19892 18376 19893 18416
rect 19851 18367 19893 18376
rect 19756 17744 19796 17753
rect 19660 17704 19756 17744
rect 19372 17536 19604 17576
rect 19179 17492 19221 17501
rect 19179 17452 19180 17492
rect 19220 17452 19221 17492
rect 19179 17443 19221 17452
rect 19084 17240 19124 17249
rect 19180 17240 19220 17443
rect 19124 17200 19220 17240
rect 19084 17191 19124 17200
rect 19275 17156 19317 17165
rect 19275 17116 19276 17156
rect 19316 17116 19317 17156
rect 19275 17107 19317 17116
rect 18892 17072 18932 17081
rect 18699 16988 18741 16997
rect 18699 16948 18700 16988
rect 18740 16948 18741 16988
rect 18699 16939 18741 16948
rect 18603 16820 18645 16829
rect 18603 16780 18604 16820
rect 18644 16780 18645 16820
rect 18603 16771 18645 16780
rect 18603 16652 18645 16661
rect 18603 16612 18604 16652
rect 18644 16612 18645 16652
rect 18603 16603 18645 16612
rect 18515 16237 18555 16246
rect 18604 16232 18644 16603
rect 18700 16484 18740 16939
rect 18892 16829 18932 17032
rect 19276 16988 19316 17107
rect 19276 16939 19316 16948
rect 18891 16820 18933 16829
rect 18891 16780 18892 16820
rect 18932 16780 18933 16820
rect 18891 16771 18933 16780
rect 19468 16820 19508 16829
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 18700 16444 18932 16484
rect 18555 16197 18644 16232
rect 18515 16192 18644 16197
rect 18700 16232 18740 16243
rect 18515 16188 18555 16192
rect 18700 16157 18740 16192
rect 18795 16232 18837 16241
rect 18795 16192 18796 16232
rect 18836 16192 18837 16232
rect 18795 16183 18837 16192
rect 18699 16148 18741 16157
rect 18699 16108 18700 16148
rect 18740 16108 18741 16148
rect 18699 16099 18741 16108
rect 18796 16098 18836 16183
rect 18604 16064 18644 16073
rect 18604 15980 18644 16024
rect 18699 15980 18741 15989
rect 18604 15940 18700 15980
rect 18740 15940 18741 15980
rect 18699 15931 18741 15940
rect 18892 15560 18932 16444
rect 19468 16409 19508 16780
rect 19467 16400 19509 16409
rect 19467 16360 19468 16400
rect 19508 16360 19509 16400
rect 19467 16351 19509 16360
rect 19179 16316 19221 16325
rect 19179 16276 19180 16316
rect 19220 16276 19221 16316
rect 19179 16267 19221 16276
rect 18988 16232 19028 16241
rect 18988 15989 19028 16192
rect 19083 16232 19125 16241
rect 19083 16192 19084 16232
rect 19124 16192 19125 16232
rect 19083 16183 19125 16192
rect 18987 15980 19029 15989
rect 18987 15940 18988 15980
rect 19028 15940 19029 15980
rect 18987 15931 19029 15940
rect 19084 15728 19124 16183
rect 19180 16064 19220 16267
rect 19372 16241 19412 16326
rect 19564 16241 19604 17536
rect 19660 17501 19700 17704
rect 19756 17695 19796 17704
rect 19852 17744 19892 18367
rect 19948 18089 19988 18544
rect 20044 18500 20084 18703
rect 20236 18618 20276 18703
rect 20044 18451 20084 18460
rect 19947 18080 19989 18089
rect 19947 18040 19948 18080
rect 19988 18040 19989 18080
rect 19947 18031 19989 18040
rect 19659 17492 19701 17501
rect 19852 17492 19892 17704
rect 20043 17744 20085 17753
rect 20043 17704 20044 17744
rect 20084 17704 20085 17744
rect 20043 17695 20085 17704
rect 19947 17660 19989 17669
rect 19947 17620 19948 17660
rect 19988 17620 19989 17660
rect 19947 17611 19989 17620
rect 19659 17452 19660 17492
rect 19700 17452 19701 17492
rect 19659 17443 19701 17452
rect 19756 17452 19892 17492
rect 19756 17072 19796 17452
rect 19851 17324 19893 17333
rect 19851 17284 19852 17324
rect 19892 17284 19893 17324
rect 19851 17275 19893 17284
rect 19852 17240 19892 17275
rect 19852 17189 19892 17200
rect 19756 17032 19892 17072
rect 19659 16988 19701 16997
rect 19659 16948 19660 16988
rect 19700 16948 19701 16988
rect 19659 16939 19701 16948
rect 19660 16854 19700 16939
rect 19756 16241 19796 16326
rect 19276 16232 19316 16241
rect 19276 16073 19316 16192
rect 19371 16232 19413 16241
rect 19371 16192 19372 16232
rect 19412 16192 19413 16232
rect 19371 16183 19413 16192
rect 19527 16232 19604 16241
rect 19567 16192 19604 16232
rect 19527 16183 19604 16192
rect 19755 16232 19797 16241
rect 19755 16192 19756 16232
rect 19796 16192 19797 16232
rect 19755 16183 19797 16192
rect 19852 16232 19892 17032
rect 19852 16183 19892 16192
rect 19180 16015 19220 16024
rect 19275 16064 19317 16073
rect 19275 16024 19276 16064
rect 19316 16024 19317 16064
rect 19275 16015 19317 16024
rect 19275 15896 19317 15905
rect 19275 15856 19276 15896
rect 19316 15856 19317 15896
rect 19275 15847 19317 15856
rect 19084 15679 19124 15688
rect 18892 15308 18932 15520
rect 19276 15476 19316 15847
rect 19276 15427 19316 15436
rect 18700 15268 18932 15308
rect 18700 14972 18740 15268
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 19180 14972 19220 14981
rect 19372 14972 19412 16183
rect 19467 15896 19509 15905
rect 19467 15856 19468 15896
rect 19508 15856 19509 15896
rect 19467 15847 19509 15856
rect 19468 15728 19508 15847
rect 19468 15679 19508 15688
rect 19564 15317 19604 16183
rect 19851 15812 19893 15821
rect 19851 15772 19852 15812
rect 19892 15772 19893 15812
rect 19851 15763 19893 15772
rect 19852 15728 19892 15763
rect 19852 15677 19892 15688
rect 19659 15476 19701 15485
rect 19659 15436 19660 15476
rect 19700 15436 19701 15476
rect 19948 15476 19988 17611
rect 20044 17576 20084 17695
rect 20044 17527 20084 17536
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 20236 17240 20276 17249
rect 20524 17240 20564 20140
rect 20276 17200 20564 17240
rect 20236 17191 20276 17200
rect 20044 16988 20084 16997
rect 20044 16493 20084 16948
rect 20043 16484 20085 16493
rect 20043 16444 20044 16484
rect 20084 16444 20085 16484
rect 20043 16435 20085 16444
rect 20044 16073 20084 16158
rect 20043 16064 20085 16073
rect 20043 16024 20044 16064
rect 20084 16024 20085 16064
rect 20043 16015 20085 16024
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 20716 15812 20756 20140
rect 21099 20131 21141 20140
rect 20907 19928 20949 19937
rect 20907 19888 20908 19928
rect 20948 19888 20949 19928
rect 20907 19879 20949 19888
rect 20811 19592 20853 19601
rect 20811 19552 20812 19592
rect 20852 19552 20853 19592
rect 20811 19543 20853 19552
rect 20524 15772 20756 15812
rect 20236 15728 20276 15737
rect 20524 15728 20564 15772
rect 20276 15688 20564 15728
rect 20236 15679 20276 15688
rect 20044 15476 20084 15485
rect 19948 15436 20044 15476
rect 19659 15427 19701 15436
rect 20044 15427 20084 15436
rect 19660 15342 19700 15427
rect 19563 15308 19605 15317
rect 19563 15268 19564 15308
rect 19604 15268 19605 15308
rect 19563 15259 19605 15268
rect 20043 15308 20085 15317
rect 20812 15308 20852 19543
rect 20043 15268 20044 15308
rect 20084 15268 20085 15308
rect 20043 15259 20085 15268
rect 20524 15268 20852 15308
rect 18700 14932 19028 14972
rect 18988 14720 19028 14932
rect 19220 14932 19412 14972
rect 20044 14972 20084 15259
rect 19180 14923 19220 14932
rect 20044 14923 20084 14932
rect 19468 14848 19796 14888
rect 19372 14729 19412 14814
rect 18699 14636 18741 14645
rect 18699 14596 18700 14636
rect 18740 14596 18741 14636
rect 18699 14587 18741 14596
rect 18603 14468 18645 14477
rect 18603 14428 18604 14468
rect 18644 14428 18645 14468
rect 18603 14419 18645 14428
rect 18412 13999 18452 14008
rect 18124 13588 18260 13628
rect 17932 12704 17972 12713
rect 17932 12545 17972 12664
rect 17931 12536 17973 12545
rect 17931 12496 17932 12536
rect 17972 12496 17973 12536
rect 17931 12487 17973 12496
rect 17932 11957 17972 12042
rect 17931 11948 17973 11957
rect 17931 11908 17932 11948
rect 17972 11908 17973 11948
rect 17931 11899 17973 11908
rect 17932 11696 17972 11705
rect 17932 11201 17972 11656
rect 18027 11276 18069 11285
rect 18027 11236 18028 11276
rect 18068 11236 18069 11276
rect 18027 11227 18069 11236
rect 17931 11192 17973 11201
rect 17931 11152 17932 11192
rect 17972 11152 17973 11192
rect 17931 11143 17973 11152
rect 17932 11024 17972 11033
rect 17835 10352 17877 10361
rect 17835 10312 17836 10352
rect 17876 10312 17877 10352
rect 17932 10352 17972 10984
rect 18028 11024 18068 11227
rect 18028 10697 18068 10984
rect 18027 10688 18069 10697
rect 18027 10648 18028 10688
rect 18068 10648 18069 10688
rect 18027 10639 18069 10648
rect 18124 10529 18164 13588
rect 18604 13208 18644 14419
rect 18604 13159 18644 13168
rect 18603 12620 18645 12629
rect 18603 12580 18604 12620
rect 18644 12580 18645 12620
rect 18603 12571 18645 12580
rect 18507 12536 18549 12545
rect 18507 12496 18508 12536
rect 18548 12496 18549 12536
rect 18507 12487 18549 12496
rect 18604 12536 18644 12571
rect 18220 11696 18260 11705
rect 18220 11537 18260 11656
rect 18219 11528 18261 11537
rect 18219 11488 18220 11528
rect 18260 11488 18261 11528
rect 18219 11479 18261 11488
rect 18508 11360 18548 12487
rect 18604 11528 18644 12496
rect 18700 11696 18740 14587
rect 18988 13805 19028 14680
rect 19371 14720 19413 14729
rect 19371 14680 19372 14720
rect 19412 14680 19413 14720
rect 19371 14671 19413 14680
rect 19468 14720 19508 14848
rect 19468 14671 19508 14680
rect 19659 14720 19701 14729
rect 19659 14680 19660 14720
rect 19700 14680 19701 14720
rect 19659 14671 19701 14680
rect 19660 14586 19700 14671
rect 19564 14552 19604 14561
rect 19372 14512 19564 14552
rect 18987 13796 19029 13805
rect 18987 13756 18988 13796
rect 19028 13756 19029 13796
rect 18987 13747 19029 13756
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 19275 13544 19317 13553
rect 19275 13504 19276 13544
rect 19316 13504 19317 13544
rect 19275 13495 19317 13504
rect 19083 13376 19125 13385
rect 19083 13336 19084 13376
rect 19124 13336 19125 13376
rect 19083 13327 19125 13336
rect 19084 13242 19124 13327
rect 19276 13301 19316 13495
rect 19275 13292 19317 13301
rect 19275 13252 19276 13292
rect 19316 13252 19317 13292
rect 19275 13243 19317 13252
rect 18796 13040 18836 13049
rect 18796 12545 18836 13000
rect 18795 12536 18837 12545
rect 18795 12496 18796 12536
rect 18836 12496 18837 12536
rect 19276 12536 19316 13243
rect 19372 13208 19412 14512
rect 19564 14503 19604 14512
rect 19659 14468 19701 14477
rect 19659 14428 19660 14468
rect 19700 14428 19701 14468
rect 19659 14419 19701 14428
rect 19660 14048 19700 14419
rect 19564 14008 19660 14048
rect 19372 13159 19412 13168
rect 19468 13208 19508 13217
rect 19468 12797 19508 13168
rect 19467 12788 19509 12797
rect 19467 12748 19468 12788
rect 19508 12748 19509 12788
rect 19467 12739 19509 12748
rect 19564 12713 19604 14008
rect 19660 13999 19700 14008
rect 19756 13376 19796 14848
rect 19851 14804 19893 14813
rect 19851 14764 19852 14804
rect 19892 14764 19893 14804
rect 19851 14755 19893 14764
rect 19852 14670 19892 14755
rect 19947 14720 19989 14729
rect 19947 14680 19948 14720
rect 19988 14680 19989 14720
rect 19947 14671 19989 14680
rect 19660 13336 19796 13376
rect 19852 13796 19892 13805
rect 19563 12704 19605 12713
rect 19563 12664 19564 12704
rect 19604 12664 19605 12704
rect 19563 12655 19605 12664
rect 19563 12536 19605 12545
rect 19276 12496 19508 12536
rect 18795 12487 18837 12496
rect 18988 12452 19028 12461
rect 18988 12284 19028 12412
rect 19084 12452 19124 12461
rect 19124 12412 19412 12452
rect 19084 12403 19124 12412
rect 18988 12244 19316 12284
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 18700 11647 18740 11656
rect 18604 11488 18740 11528
rect 18508 11320 18644 11360
rect 18219 11276 18261 11285
rect 18219 11236 18220 11276
rect 18260 11236 18261 11276
rect 18219 11227 18261 11236
rect 18220 11044 18260 11227
rect 18220 11024 18273 11044
rect 18508 11033 18548 11118
rect 18412 11024 18452 11033
rect 18220 11014 18281 11024
rect 18220 11004 18412 11014
rect 18233 10984 18412 11004
rect 18241 10974 18452 10984
rect 18507 11024 18549 11033
rect 18507 10984 18508 11024
rect 18548 10984 18549 11024
rect 18507 10975 18549 10984
rect 18219 10856 18261 10865
rect 18219 10816 18220 10856
rect 18260 10816 18261 10856
rect 18219 10807 18261 10816
rect 18123 10520 18165 10529
rect 18123 10480 18124 10520
rect 18164 10480 18165 10520
rect 18123 10471 18165 10480
rect 17932 10312 18164 10352
rect 17835 10303 17877 10312
rect 17740 10135 17780 10144
rect 17836 10184 17876 10193
rect 17644 9976 17780 10016
rect 17356 9857 17396 9976
rect 17355 9848 17397 9857
rect 17355 9808 17356 9848
rect 17396 9808 17397 9848
rect 17355 9799 17397 9808
rect 17356 9344 17396 9799
rect 17643 9512 17685 9521
rect 17643 9472 17644 9512
rect 17684 9472 17685 9512
rect 17643 9463 17685 9472
rect 17644 9378 17684 9463
rect 17356 8504 17396 9304
rect 17644 8681 17684 8766
rect 17643 8672 17685 8681
rect 17643 8632 17644 8672
rect 17684 8632 17685 8672
rect 17643 8623 17685 8632
rect 17259 8168 17301 8177
rect 17259 8128 17260 8168
rect 17300 8128 17301 8168
rect 17259 8119 17301 8128
rect 17356 7832 17396 8464
rect 17643 8504 17685 8513
rect 17643 8464 17644 8504
rect 17684 8464 17685 8504
rect 17643 8455 17685 8464
rect 17644 8000 17684 8455
rect 17644 7951 17684 7960
rect 16396 6952 16628 6992
rect 16972 7165 17012 7174
rect 16300 6488 16340 6497
rect 16396 6488 16436 6952
rect 16972 6740 17012 7125
rect 17356 7160 17396 7792
rect 17163 7076 17205 7085
rect 17163 7036 17164 7076
rect 17204 7036 17205 7076
rect 17163 7027 17205 7036
rect 17164 6942 17204 7027
rect 16492 6700 17012 6740
rect 16492 6656 16532 6700
rect 16492 6607 16532 6616
rect 16683 6572 16725 6581
rect 16683 6532 16684 6572
rect 16724 6532 16725 6572
rect 16683 6523 16725 6532
rect 16340 6448 16436 6488
rect 16300 6439 16340 6448
rect 16396 6245 16436 6448
rect 16491 6488 16533 6497
rect 16491 6448 16492 6488
rect 16532 6448 16533 6488
rect 16491 6439 16533 6448
rect 16395 6236 16437 6245
rect 16395 6196 16396 6236
rect 16436 6196 16437 6236
rect 16395 6187 16437 6196
rect 16395 1868 16437 1877
rect 16395 1828 16396 1868
rect 16436 1828 16437 1868
rect 16395 1819 16437 1828
rect 16396 1734 16436 1819
rect 16203 1700 16245 1709
rect 16203 1660 16204 1700
rect 16244 1660 16245 1700
rect 16203 1651 16245 1660
rect 16204 1566 16244 1651
rect 16108 1324 16244 1364
rect 15916 1240 16052 1280
rect 15915 944 15957 953
rect 15915 904 15916 944
rect 15956 904 15957 944
rect 15915 895 15957 904
rect 15916 810 15956 895
rect 16012 80 16052 1240
rect 16107 1196 16149 1205
rect 16107 1156 16108 1196
rect 16148 1156 16149 1196
rect 16107 1147 16149 1156
rect 16108 1062 16148 1147
rect 16204 80 16244 1324
rect 16492 1112 16532 6439
rect 16588 1700 16628 1709
rect 16588 1457 16628 1660
rect 16587 1448 16629 1457
rect 16587 1408 16588 1448
rect 16628 1408 16629 1448
rect 16587 1399 16629 1408
rect 16684 1280 16724 6523
rect 16875 6404 16917 6413
rect 16875 6364 16876 6404
rect 16916 6364 16917 6404
rect 16875 6355 16917 6364
rect 16779 1868 16821 1877
rect 16779 1828 16780 1868
rect 16820 1828 16821 1868
rect 16779 1819 16821 1828
rect 16780 1734 16820 1819
rect 16396 1072 16532 1112
rect 16588 1240 16724 1280
rect 16396 80 16436 1072
rect 16588 80 16628 1240
rect 16876 1112 16916 6355
rect 16971 6320 17013 6329
rect 16971 6280 16972 6320
rect 17012 6280 17013 6320
rect 16971 6271 17013 6280
rect 17356 6320 17396 7120
rect 16780 1072 16916 1112
rect 16780 80 16820 1072
rect 16972 80 17012 6271
rect 17163 6236 17205 6245
rect 17163 6196 17164 6236
rect 17204 6196 17205 6236
rect 17163 6187 17205 6196
rect 17164 80 17204 6187
rect 17356 5480 17396 6280
rect 17356 4808 17396 5440
rect 17356 3968 17396 4768
rect 17356 3641 17396 3928
rect 17355 3632 17397 3641
rect 17355 3592 17356 3632
rect 17396 3592 17397 3632
rect 17355 3583 17397 3592
rect 17356 3498 17396 3583
rect 17259 2120 17301 2129
rect 17259 2080 17260 2120
rect 17300 2080 17301 2120
rect 17259 2071 17301 2080
rect 17643 2120 17685 2129
rect 17643 2080 17644 2120
rect 17684 2080 17685 2120
rect 17643 2071 17685 2080
rect 17260 1986 17300 2071
rect 17644 1986 17684 2071
rect 17452 1868 17492 1877
rect 17356 1828 17452 1868
rect 17356 80 17396 1828
rect 17452 1819 17492 1828
rect 17547 1868 17589 1877
rect 17547 1828 17548 1868
rect 17588 1828 17589 1868
rect 17547 1819 17589 1828
rect 17548 80 17588 1819
rect 17740 1784 17780 9976
rect 17836 8849 17876 10144
rect 17931 10184 17973 10193
rect 17931 10144 17932 10184
rect 17972 10144 17973 10184
rect 17931 10135 17973 10144
rect 18028 10184 18068 10193
rect 17932 10050 17972 10135
rect 18028 10025 18068 10144
rect 18027 10016 18069 10025
rect 18027 9976 18028 10016
rect 18068 9976 18069 10016
rect 18027 9967 18069 9976
rect 17931 9848 17973 9857
rect 17931 9808 17932 9848
rect 17972 9808 17973 9848
rect 17931 9799 17973 9808
rect 17835 8840 17877 8849
rect 17835 8800 17836 8840
rect 17876 8800 17877 8840
rect 17835 8791 17877 8800
rect 17932 6497 17972 9799
rect 18027 9764 18069 9773
rect 18027 9724 18028 9764
rect 18068 9724 18069 9764
rect 18027 9715 18069 9724
rect 18028 6581 18068 9715
rect 18124 9689 18164 10312
rect 18220 10184 18260 10807
rect 18604 10604 18644 11320
rect 18412 10564 18644 10604
rect 18315 10520 18357 10529
rect 18315 10480 18316 10520
rect 18356 10480 18357 10520
rect 18315 10471 18357 10480
rect 18316 10268 18356 10471
rect 18316 10219 18356 10228
rect 18220 10135 18260 10144
rect 18412 10100 18452 10564
rect 18603 10436 18645 10445
rect 18603 10396 18604 10436
rect 18644 10396 18645 10436
rect 18603 10387 18645 10396
rect 18604 10268 18644 10387
rect 18700 10352 18740 11488
rect 19276 11360 19316 12244
rect 19372 12125 19412 12412
rect 19371 12116 19413 12125
rect 19371 12076 19372 12116
rect 19412 12076 19413 12116
rect 19371 12067 19413 12076
rect 19372 11873 19412 12067
rect 19371 11864 19413 11873
rect 19371 11824 19372 11864
rect 19412 11824 19413 11864
rect 19371 11815 19413 11824
rect 19276 11320 19412 11360
rect 18891 11276 18933 11285
rect 18891 11236 18892 11276
rect 18932 11236 18933 11276
rect 18891 11227 18933 11236
rect 18892 11024 18932 11227
rect 18892 10865 18932 10984
rect 18988 10940 19028 10949
rect 19028 10900 19316 10940
rect 18988 10891 19028 10900
rect 18891 10856 18933 10865
rect 18891 10816 18892 10856
rect 18932 10816 18933 10856
rect 18891 10807 18933 10816
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 18700 10312 18836 10352
rect 18604 10228 18740 10268
rect 18700 10184 18740 10228
rect 18509 10169 18549 10178
rect 18700 10135 18740 10144
rect 18509 10100 18549 10129
rect 18412 10060 18549 10100
rect 18509 10016 18549 10060
rect 18508 9976 18549 10016
rect 18603 10016 18645 10025
rect 18796 10016 18836 10312
rect 18891 10268 18933 10277
rect 18891 10228 18892 10268
rect 18932 10228 18933 10268
rect 18891 10219 18933 10228
rect 18603 9976 18604 10016
rect 18644 9976 18645 10016
rect 18123 9680 18165 9689
rect 18123 9640 18124 9680
rect 18164 9640 18165 9680
rect 18123 9631 18165 9640
rect 18508 9353 18548 9976
rect 18603 9967 18645 9976
rect 18700 9976 18836 10016
rect 18507 9344 18549 9353
rect 18507 9304 18508 9344
rect 18548 9304 18549 9344
rect 18507 9295 18549 9304
rect 18604 7328 18644 9967
rect 18508 7288 18644 7328
rect 18027 6572 18069 6581
rect 18027 6532 18028 6572
rect 18068 6532 18069 6572
rect 18027 6523 18069 6532
rect 17931 6488 17973 6497
rect 17931 6448 17932 6488
rect 17972 6448 17973 6488
rect 17931 6439 17973 6448
rect 18508 2540 18548 7288
rect 18700 7169 18740 9976
rect 18892 9512 18932 10219
rect 19276 9773 19316 10900
rect 19275 9764 19317 9773
rect 19275 9724 19276 9764
rect 19316 9724 19317 9764
rect 19275 9715 19317 9724
rect 19372 9689 19412 11320
rect 19468 11024 19508 12496
rect 19563 12496 19564 12536
rect 19604 12496 19605 12536
rect 19563 12487 19605 12496
rect 19564 12377 19604 12487
rect 19563 12368 19605 12377
rect 19563 12328 19564 12368
rect 19604 12328 19605 12368
rect 19563 12319 19605 12328
rect 19468 10975 19508 10984
rect 19467 9848 19509 9857
rect 19467 9808 19468 9848
rect 19508 9808 19509 9848
rect 19467 9799 19509 9808
rect 19083 9680 19125 9689
rect 19083 9640 19084 9680
rect 19124 9640 19125 9680
rect 19083 9631 19125 9640
rect 19371 9680 19413 9689
rect 19371 9640 19372 9680
rect 19412 9640 19413 9680
rect 19371 9631 19413 9640
rect 19084 9546 19124 9631
rect 18892 9463 18932 9472
rect 19366 9512 19408 9521
rect 19366 9472 19367 9512
rect 19407 9472 19408 9512
rect 19366 9463 19408 9472
rect 19468 9512 19508 9799
rect 19468 9463 19508 9472
rect 19563 9512 19605 9521
rect 19563 9472 19564 9512
rect 19604 9472 19605 9512
rect 19563 9463 19605 9472
rect 19084 9269 19124 9354
rect 19083 9260 19125 9269
rect 19083 9220 19084 9260
rect 19124 9220 19125 9260
rect 19083 9211 19125 9220
rect 19367 9176 19407 9463
rect 19564 9378 19604 9463
rect 19660 9437 19700 13336
rect 19756 13208 19796 13217
rect 19852 13208 19892 13756
rect 19796 13168 19892 13208
rect 19756 13159 19796 13168
rect 19851 12704 19893 12713
rect 19851 12664 19852 12704
rect 19892 12664 19893 12704
rect 19948 12704 19988 14671
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 20236 14216 20276 14225
rect 20524 14216 20564 15268
rect 20908 15056 20948 19879
rect 21099 16316 21141 16325
rect 21099 16276 21100 16316
rect 21140 16276 21141 16316
rect 21099 16267 21141 16276
rect 21003 16232 21045 16241
rect 21003 16192 21004 16232
rect 21044 16192 21045 16232
rect 21003 16183 21045 16192
rect 20276 14176 20564 14216
rect 20620 15016 20948 15056
rect 20236 14167 20276 14176
rect 20620 14048 20660 15016
rect 20811 14888 20853 14897
rect 20811 14848 20812 14888
rect 20852 14848 20853 14888
rect 20811 14839 20853 14848
rect 20236 14008 20660 14048
rect 20043 13964 20085 13973
rect 20043 13924 20044 13964
rect 20084 13924 20085 13964
rect 20043 13915 20085 13924
rect 20044 13830 20084 13915
rect 20236 13460 20276 14008
rect 20715 13712 20757 13721
rect 20715 13672 20716 13712
rect 20756 13672 20757 13712
rect 20715 13663 20757 13672
rect 20236 13411 20276 13420
rect 20043 13292 20085 13301
rect 20043 13252 20044 13292
rect 20084 13252 20085 13292
rect 20043 13243 20085 13252
rect 20044 13158 20084 13243
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 19948 12664 20084 12704
rect 19851 12655 19893 12664
rect 19852 11696 19892 12655
rect 20044 12531 20084 12664
rect 20235 12620 20277 12629
rect 20235 12580 20236 12620
rect 20276 12580 20277 12620
rect 20235 12571 20277 12580
rect 20044 11948 20084 12491
rect 20236 12486 20276 12571
rect 20140 11948 20180 11957
rect 20044 11908 20140 11948
rect 20140 11880 20180 11908
rect 19948 11696 19988 11705
rect 19852 11656 19948 11696
rect 19852 10268 19892 11656
rect 19948 11647 19988 11656
rect 20048 11360 20416 11369
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 20140 11108 20180 11117
rect 20180 11068 20660 11108
rect 20140 11059 20180 11068
rect 19996 10982 20036 10991
rect 19996 10940 20036 10942
rect 19996 10900 20180 10940
rect 19947 10268 19989 10277
rect 19852 10228 19948 10268
rect 19988 10228 19989 10268
rect 19947 10219 19989 10228
rect 19948 10184 19988 10219
rect 20140 10193 20180 10900
rect 19948 10133 19988 10144
rect 20139 10184 20181 10193
rect 20139 10144 20140 10184
rect 20180 10144 20181 10184
rect 20139 10135 20181 10144
rect 20140 10100 20180 10135
rect 20140 10049 20180 10060
rect 20620 10016 20660 11068
rect 20716 10193 20756 13663
rect 20812 12545 20852 14839
rect 20811 12536 20853 12545
rect 20811 12496 20812 12536
rect 20852 12496 20853 12536
rect 20811 12487 20853 12496
rect 20715 10184 20757 10193
rect 20715 10144 20716 10184
rect 20756 10144 20757 10184
rect 20715 10135 20757 10144
rect 20620 9976 20756 10016
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 20044 9521 20084 9606
rect 19756 9512 19796 9521
rect 19659 9428 19701 9437
rect 19659 9388 19660 9428
rect 19700 9388 19701 9428
rect 19659 9379 19701 9388
rect 19467 9260 19509 9269
rect 19467 9220 19468 9260
rect 19508 9220 19509 9260
rect 19467 9211 19509 9220
rect 19367 9136 19412 9176
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 19372 9017 19412 9136
rect 19371 9008 19413 9017
rect 19371 8968 19372 9008
rect 19412 8968 19413 9008
rect 19371 8959 19413 8968
rect 19083 8924 19125 8933
rect 19083 8884 19084 8924
rect 19124 8884 19125 8924
rect 19083 8875 19125 8884
rect 19084 8790 19124 8875
rect 18892 8672 18932 8681
rect 18892 8009 18932 8632
rect 19276 8672 19316 8681
rect 19084 8504 19124 8513
rect 19124 8464 19220 8504
rect 19084 8455 19124 8464
rect 18891 8000 18933 8009
rect 18891 7960 18892 8000
rect 18932 7960 18933 8000
rect 18891 7951 18933 7960
rect 18892 7866 18932 7951
rect 19180 7925 19220 8464
rect 19179 7916 19221 7925
rect 19179 7876 19180 7916
rect 19220 7876 19221 7916
rect 19179 7867 19221 7876
rect 19084 7757 19124 7842
rect 19083 7748 19125 7757
rect 19083 7708 19084 7748
rect 19124 7708 19125 7748
rect 19083 7699 19125 7708
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 18987 7412 19029 7421
rect 18987 7372 18988 7412
rect 19028 7372 19029 7412
rect 18987 7363 19029 7372
rect 18795 7328 18837 7337
rect 18795 7288 18796 7328
rect 18836 7288 18837 7328
rect 18795 7279 18837 7288
rect 18796 7194 18836 7279
rect 18604 7160 18644 7169
rect 18604 7001 18644 7120
rect 18699 7160 18741 7169
rect 18699 7120 18700 7160
rect 18740 7120 18741 7160
rect 18699 7111 18741 7120
rect 18988 7160 19028 7363
rect 19276 7328 19316 8632
rect 19372 8672 19412 8681
rect 19372 7337 19412 8632
rect 19468 8000 19508 9211
rect 19756 8933 19796 9472
rect 19852 9512 19892 9521
rect 20043 9512 20085 9521
rect 19892 9472 19988 9512
rect 19852 9463 19892 9472
rect 19948 9344 19988 9472
rect 20043 9472 20044 9512
rect 20084 9472 20085 9512
rect 20043 9463 20085 9472
rect 20236 9512 20276 9521
rect 20139 9428 20181 9437
rect 20139 9388 20140 9428
rect 20180 9388 20181 9428
rect 20139 9379 20181 9388
rect 19948 9304 20084 9344
rect 19852 9260 19892 9269
rect 19892 9220 19988 9260
rect 19852 9211 19892 9220
rect 19851 9008 19893 9017
rect 19851 8968 19852 9008
rect 19892 8968 19893 9008
rect 19851 8959 19893 8968
rect 19755 8924 19797 8933
rect 19755 8884 19756 8924
rect 19796 8884 19797 8924
rect 19755 8875 19797 8884
rect 19852 8756 19892 8959
rect 19817 8716 19892 8756
rect 19948 8756 19988 9220
rect 20044 8924 20084 9304
rect 20140 9294 20180 9379
rect 20236 9353 20276 9472
rect 20235 9344 20277 9353
rect 20235 9304 20236 9344
rect 20276 9304 20277 9344
rect 20235 9295 20277 9304
rect 20523 9176 20565 9185
rect 20523 9136 20524 9176
rect 20564 9136 20565 9176
rect 20523 9127 20565 9136
rect 20235 8924 20277 8933
rect 20044 8884 20180 8924
rect 20044 8756 20084 8765
rect 19948 8716 20044 8756
rect 19817 8687 19857 8716
rect 20044 8707 20084 8716
rect 19563 8672 19605 8681
rect 19563 8632 19564 8672
rect 19604 8632 19605 8672
rect 19563 8623 19605 8632
rect 19660 8672 19700 8681
rect 19817 8638 19857 8647
rect 19564 8538 19604 8623
rect 19468 7951 19508 7960
rect 19563 8000 19605 8009
rect 19563 7960 19564 8000
rect 19604 7960 19605 8000
rect 19563 7951 19605 7960
rect 19564 7866 19604 7951
rect 19276 7279 19316 7288
rect 19371 7328 19413 7337
rect 19371 7288 19372 7328
rect 19412 7288 19413 7328
rect 19371 7279 19413 7288
rect 18988 7111 19028 7120
rect 19180 7160 19220 7169
rect 18603 6992 18645 7001
rect 18603 6952 18604 6992
rect 18644 6952 18645 6992
rect 18603 6943 18645 6952
rect 18604 6413 18644 6943
rect 19180 6908 19220 7120
rect 19276 7160 19316 7169
rect 19316 7120 19321 7160
rect 19276 7111 19321 7120
rect 19281 7076 19321 7111
rect 19372 7076 19412 7279
rect 19660 7160 19700 8632
rect 20140 8588 20180 8884
rect 20235 8884 20236 8924
rect 20276 8884 20277 8924
rect 20235 8875 20277 8884
rect 20236 8840 20276 8875
rect 20236 8789 20276 8800
rect 19948 8548 20180 8588
rect 19756 8504 19796 8513
rect 19796 8464 19892 8504
rect 19756 8455 19796 8464
rect 19755 8168 19797 8177
rect 19755 8128 19756 8168
rect 19796 8128 19797 8168
rect 19755 8119 19797 8128
rect 19756 8034 19796 8119
rect 19755 7832 19797 7841
rect 19755 7792 19756 7832
rect 19796 7792 19797 7832
rect 19755 7783 19797 7792
rect 19756 7664 19796 7783
rect 19852 7748 19892 8464
rect 19948 8177 19988 8548
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19947 8168 19989 8177
rect 19947 8128 19948 8168
rect 19988 8128 19989 8168
rect 19947 8119 19989 8128
rect 20139 8168 20181 8177
rect 20524 8168 20564 9127
rect 20716 8177 20756 9976
rect 20139 8128 20140 8168
rect 20180 8128 20181 8168
rect 20139 8119 20181 8128
rect 20236 8128 20564 8168
rect 20715 8168 20757 8177
rect 20715 8128 20716 8168
rect 20756 8128 20757 8168
rect 20140 8034 20180 8119
rect 19947 8000 19989 8009
rect 19947 7960 19948 8000
rect 19988 7960 19989 8000
rect 19947 7951 19989 7960
rect 20044 8000 20084 8011
rect 19948 7866 19988 7951
rect 20044 7925 20084 7960
rect 20236 8000 20276 8128
rect 20715 8119 20757 8128
rect 21004 8000 21044 16183
rect 21100 9932 21140 16267
rect 21196 15821 21236 21223
rect 21291 20600 21333 20609
rect 21291 20560 21292 20600
rect 21332 20560 21333 20600
rect 21291 20551 21333 20560
rect 21292 15989 21332 20551
rect 21387 20096 21429 20105
rect 21387 20056 21388 20096
rect 21428 20056 21429 20096
rect 21387 20047 21429 20056
rect 21291 15980 21333 15989
rect 21291 15940 21292 15980
rect 21332 15940 21333 15980
rect 21291 15931 21333 15940
rect 21195 15812 21237 15821
rect 21195 15772 21196 15812
rect 21236 15772 21237 15812
rect 21195 15763 21237 15772
rect 21388 15401 21428 20047
rect 21387 15392 21429 15401
rect 21387 15352 21388 15392
rect 21428 15352 21429 15392
rect 21387 15343 21429 15352
rect 21195 13460 21237 13469
rect 21195 13420 21196 13460
rect 21236 13420 21237 13460
rect 21195 13411 21237 13420
rect 21196 10529 21236 13411
rect 21195 10520 21237 10529
rect 21195 10480 21196 10520
rect 21236 10480 21237 10520
rect 21195 10471 21237 10480
rect 21100 9892 21236 9932
rect 21099 9764 21141 9773
rect 21099 9724 21100 9764
rect 21140 9724 21141 9764
rect 21099 9715 21141 9724
rect 21100 8177 21140 9715
rect 21196 8933 21236 9892
rect 21195 8924 21237 8933
rect 21195 8884 21196 8924
rect 21236 8884 21237 8924
rect 21195 8875 21237 8884
rect 21099 8168 21141 8177
rect 21099 8128 21100 8168
rect 21140 8128 21141 8168
rect 21099 8119 21141 8128
rect 20236 7951 20276 7960
rect 20332 7960 21044 8000
rect 20043 7916 20085 7925
rect 20043 7876 20044 7916
rect 20084 7876 20085 7916
rect 20043 7867 20085 7876
rect 19852 7708 20084 7748
rect 19756 7624 19892 7664
rect 19281 7036 19412 7076
rect 19468 7120 19700 7160
rect 19468 6908 19508 7120
rect 19563 6992 19605 7001
rect 19563 6952 19564 6992
rect 19604 6952 19605 6992
rect 19563 6943 19605 6952
rect 19180 6868 19508 6908
rect 19564 6858 19604 6943
rect 18699 6740 18741 6749
rect 18699 6700 18700 6740
rect 18740 6700 18741 6740
rect 18699 6691 18741 6700
rect 19563 6740 19605 6749
rect 19563 6700 19564 6740
rect 19604 6700 19605 6740
rect 19563 6691 19605 6700
rect 18700 6488 18740 6691
rect 18700 6439 18740 6448
rect 18603 6404 18645 6413
rect 18603 6364 18604 6404
rect 18644 6364 18645 6404
rect 18603 6355 18645 6364
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19564 5648 19604 6691
rect 19660 6656 19700 7120
rect 19756 7160 19796 7169
rect 19756 6833 19796 7120
rect 19852 7160 19892 7624
rect 20044 7244 20084 7708
rect 20236 7412 20276 7421
rect 20332 7412 20372 7960
rect 20276 7372 20372 7412
rect 20236 7363 20276 7372
rect 20044 7195 20084 7204
rect 19852 7111 19892 7120
rect 19755 6824 19797 6833
rect 19755 6784 19756 6824
rect 19796 6784 19797 6824
rect 19755 6775 19797 6784
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20140 6656 20180 6665
rect 19660 6616 20140 6656
rect 19660 5648 19700 5657
rect 19564 5608 19660 5648
rect 19660 5599 19700 5608
rect 19756 5648 19796 6616
rect 20140 6607 20180 6616
rect 19948 6488 19988 6499
rect 19948 6413 19988 6448
rect 19947 6404 19989 6413
rect 19947 6364 19948 6404
rect 19988 6364 19989 6404
rect 19947 6355 19989 6364
rect 19756 5599 19796 5608
rect 19467 5480 19509 5489
rect 19467 5440 19468 5480
rect 19508 5440 19509 5480
rect 19467 5431 19509 5440
rect 19468 5346 19508 5431
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 19947 5060 19989 5069
rect 19947 5020 19948 5060
rect 19988 5020 19989 5060
rect 19947 5011 19989 5020
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 18508 2500 18740 2540
rect 18027 2120 18069 2129
rect 18027 2080 18028 2120
rect 18068 2080 18069 2120
rect 18027 2071 18069 2080
rect 18411 2120 18453 2129
rect 18411 2080 18412 2120
rect 18452 2080 18453 2120
rect 18411 2071 18453 2080
rect 18028 1986 18068 2071
rect 18412 1986 18452 2071
rect 17835 1868 17877 1877
rect 18220 1868 18260 1877
rect 18604 1868 18644 1877
rect 17835 1828 17836 1868
rect 17876 1828 17877 1868
rect 17835 1819 17877 1828
rect 17932 1828 18220 1868
rect 17644 1744 17780 1784
rect 17644 197 17684 1744
rect 17836 1734 17876 1819
rect 17932 524 17972 1828
rect 18220 1819 18260 1828
rect 18316 1828 18604 1868
rect 18027 1280 18069 1289
rect 18027 1240 18028 1280
rect 18068 1240 18069 1280
rect 18027 1231 18069 1240
rect 18028 1146 18068 1231
rect 18220 1196 18260 1205
rect 18124 1156 18220 1196
rect 17740 484 17972 524
rect 17643 188 17685 197
rect 17643 148 17644 188
rect 17684 148 17685 188
rect 17643 139 17685 148
rect 17740 80 17780 484
rect 17931 356 17973 365
rect 17931 316 17932 356
rect 17972 316 17973 356
rect 17931 307 17973 316
rect 17932 80 17972 307
rect 18124 80 18164 1156
rect 18220 1147 18260 1156
rect 18316 365 18356 1828
rect 18604 1819 18644 1828
rect 18507 1700 18549 1709
rect 18507 1660 18508 1700
rect 18548 1660 18549 1700
rect 18507 1651 18549 1660
rect 18508 1373 18548 1651
rect 18507 1364 18549 1373
rect 18507 1324 18508 1364
rect 18548 1324 18549 1364
rect 18507 1315 18549 1324
rect 18411 1280 18453 1289
rect 18411 1240 18412 1280
rect 18452 1240 18453 1280
rect 18700 1280 18740 2500
rect 18795 2288 18837 2297
rect 18795 2248 18796 2288
rect 18836 2248 18837 2288
rect 18795 2239 18837 2248
rect 18796 2120 18836 2239
rect 18796 2071 18836 2080
rect 19179 2120 19221 2129
rect 19179 2080 19180 2120
rect 19220 2080 19221 2120
rect 19179 2071 19221 2080
rect 19563 2120 19605 2129
rect 19563 2080 19564 2120
rect 19604 2080 19605 2120
rect 19563 2071 19605 2080
rect 19948 2120 19988 5011
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19948 2071 19988 2080
rect 19180 1986 19220 2071
rect 19564 1986 19604 2071
rect 18988 1868 19028 1877
rect 18988 1709 19028 1828
rect 19372 1868 19412 1877
rect 19756 1868 19796 1877
rect 18987 1700 19029 1709
rect 18987 1660 18988 1700
rect 19028 1660 19029 1700
rect 18987 1651 19029 1660
rect 19372 1541 19412 1828
rect 19468 1828 19756 1868
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 19371 1532 19413 1541
rect 19371 1492 19372 1532
rect 19412 1492 19413 1532
rect 19371 1483 19413 1492
rect 19468 1364 19508 1828
rect 19756 1819 19796 1828
rect 20121 1865 20161 1874
rect 20121 1532 20161 1825
rect 21291 1784 21333 1793
rect 21291 1744 21292 1784
rect 21332 1744 21333 1784
rect 21291 1735 21333 1744
rect 19084 1324 19508 1364
rect 19948 1492 20161 1532
rect 18796 1280 18836 1289
rect 18700 1240 18796 1280
rect 18411 1231 18453 1240
rect 18796 1231 18836 1240
rect 18412 1146 18452 1231
rect 18604 1196 18644 1205
rect 18988 1196 19028 1205
rect 18508 1156 18604 1196
rect 18411 1028 18453 1037
rect 18411 988 18412 1028
rect 18452 988 18453 1028
rect 18411 979 18453 988
rect 18315 356 18357 365
rect 18315 316 18316 356
rect 18356 316 18357 356
rect 18315 307 18357 316
rect 18412 188 18452 979
rect 18316 148 18452 188
rect 18316 80 18356 148
rect 18508 80 18548 1156
rect 18604 1147 18644 1156
rect 18892 1156 18988 1196
rect 18699 1112 18741 1121
rect 18699 1072 18700 1112
rect 18740 1072 18741 1112
rect 18699 1063 18741 1072
rect 18700 80 18740 1063
rect 18892 80 18932 1156
rect 18988 1147 19028 1156
rect 19084 80 19124 1324
rect 19372 1196 19412 1205
rect 19276 1156 19372 1196
rect 19179 944 19221 953
rect 19179 904 19180 944
rect 19220 904 19221 944
rect 19179 895 19221 904
rect 19180 810 19220 895
rect 19276 80 19316 1156
rect 19372 1147 19412 1156
rect 19468 80 19700 104
rect 7028 64 7048 80
rect 6968 0 7048 64
rect 7160 0 7240 80
rect 7352 0 7432 80
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 0 8008 80
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 64 19700 80
rect 19448 0 19528 64
rect 19660 60 19700 64
rect 19948 60 19988 1492
rect 21292 1448 21332 1735
rect 21387 1448 21429 1457
rect 21292 1408 21388 1448
rect 21428 1408 21429 1448
rect 21387 1399 21429 1408
rect 20523 1364 20565 1373
rect 20523 1324 20524 1364
rect 20564 1324 20565 1364
rect 20523 1315 20565 1324
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 20524 449 20564 1315
rect 20523 440 20565 449
rect 20523 400 20524 440
rect 20564 400 20565 440
rect 20523 391 20565 400
rect 19660 20 19988 60
<< via2 >>
rect 1036 85072 1076 85112
rect 172 78520 212 78560
rect 76 66424 116 66464
rect 268 73816 308 73856
rect 844 70456 884 70496
rect 844 65500 884 65540
rect 748 65080 788 65120
rect 268 60964 308 61004
rect 172 59788 212 59828
rect 364 59704 404 59744
rect 172 59032 212 59072
rect 172 46600 212 46640
rect 940 60376 980 60416
rect 2188 83560 2228 83600
rect 1516 83476 1556 83516
rect 2092 83476 2132 83516
rect 2668 83560 2708 83600
rect 3436 84820 3476 84860
rect 3436 84400 3476 84440
rect 3340 83812 3380 83852
rect 3724 84820 3764 84860
rect 4108 84988 4148 85028
rect 3688 84652 3728 84692
rect 3770 84652 3810 84692
rect 3852 84652 3892 84692
rect 3934 84652 3974 84692
rect 4016 84652 4056 84692
rect 4396 84988 4436 85028
rect 4108 83812 4148 83852
rect 2860 83476 2900 83516
rect 2860 82804 2900 82844
rect 3244 82804 3284 82844
rect 2380 81124 2420 81164
rect 1516 72724 1556 72764
rect 1324 72304 1364 72344
rect 1324 70372 1364 70412
rect 1516 69952 1556 69992
rect 1324 67348 1364 67388
rect 1228 66928 1268 66968
rect 1420 66088 1460 66128
rect 1132 64408 1172 64448
rect 1036 54160 1076 54200
rect 364 44416 404 44456
rect 748 41728 788 41768
rect 172 38452 212 38492
rect 76 36604 116 36644
rect 76 35512 116 35552
rect 652 37276 692 37316
rect 940 41392 980 41432
rect 844 40384 884 40424
rect 844 39880 884 39920
rect 748 33748 788 33788
rect 652 31480 692 31520
rect 268 29212 308 29252
rect 268 20056 308 20096
rect 460 19552 500 19592
rect 172 17368 212 17408
rect 364 16528 404 16568
rect 76 10312 116 10352
rect 1324 62308 1364 62348
rect 1996 74488 2036 74528
rect 1900 73144 1940 73184
rect 1804 65500 1844 65540
rect 1708 64072 1748 64112
rect 1708 62812 1748 62852
rect 1708 62308 1748 62348
rect 1612 61888 1652 61928
rect 1516 61468 1556 61508
rect 1420 60544 1460 60584
rect 1324 59368 1364 59408
rect 1612 60796 1652 60836
rect 1516 57604 1556 57644
rect 1324 56596 1364 56636
rect 1420 56008 1460 56048
rect 1324 55672 1364 55712
rect 1420 54916 1460 54956
rect 1420 54328 1460 54368
rect 1708 57604 1748 57644
rect 1612 56512 1652 56552
rect 1612 55000 1652 55040
rect 1228 53656 1268 53696
rect 1324 53320 1364 53360
rect 1516 52816 1556 52856
rect 1420 52564 1460 52604
rect 1420 51808 1460 51848
rect 1324 50884 1364 50924
rect 1420 50212 1460 50252
rect 1420 49624 1460 49664
rect 1324 48952 1364 48992
rect 1708 50296 1748 50336
rect 1612 50128 1652 50168
rect 1516 48952 1556 48992
rect 1324 48196 1364 48236
rect 1708 47944 1748 47984
rect 1612 46936 1652 46976
rect 1420 46768 1460 46808
rect 1324 46600 1364 46640
rect 1228 45592 1268 45632
rect 1708 46600 1748 46640
rect 1324 41476 1364 41516
rect 1228 37864 1268 37904
rect 1324 37192 1364 37232
rect 1228 36688 1268 36728
rect 1228 35428 1268 35468
rect 1228 34336 1268 34376
rect 1036 33748 1076 33788
rect 940 15436 980 15476
rect 844 15016 884 15056
rect 2284 70792 2324 70832
rect 2092 67768 2132 67808
rect 1996 62644 2036 62684
rect 1900 61132 1940 61172
rect 1996 60544 2036 60584
rect 1900 57016 1940 57056
rect 2476 72388 2516 72428
rect 2284 66928 2324 66968
rect 2476 70036 2516 70076
rect 2476 67600 2516 67640
rect 2572 67432 2612 67472
rect 2956 70708 2996 70748
rect 2956 69112 2996 69152
rect 4012 83476 4052 83516
rect 3628 83308 3668 83348
rect 3688 83140 3728 83180
rect 3770 83140 3810 83180
rect 3852 83140 3892 83180
rect 3934 83140 3974 83180
rect 4016 83140 4056 83180
rect 4300 84400 4340 84440
rect 4492 84316 4532 84356
rect 5068 84652 5108 84692
rect 5644 85156 5684 85196
rect 5260 84568 5300 84608
rect 4876 84064 4916 84104
rect 5356 84064 5396 84104
rect 4928 83896 4968 83936
rect 5010 83896 5050 83936
rect 5092 83896 5132 83936
rect 5174 83896 5214 83936
rect 5256 83896 5296 83936
rect 6028 85072 6068 85112
rect 6412 85576 6452 85616
rect 6604 84484 6644 84524
rect 5836 84400 5876 84440
rect 6220 84400 6260 84440
rect 6796 84400 6836 84440
rect 6604 83812 6644 83852
rect 4396 83308 4436 83348
rect 5548 83644 5588 83684
rect 6124 83476 6164 83516
rect 5164 83224 5204 83264
rect 4780 83140 4820 83180
rect 5548 83140 5588 83180
rect 6508 83140 6548 83180
rect 3628 82804 3668 82844
rect 4108 82804 4148 82844
rect 4780 82804 4820 82844
rect 4928 82384 4968 82424
rect 5010 82384 5050 82424
rect 5092 82384 5132 82424
rect 5174 82384 5214 82424
rect 5256 82384 5296 82424
rect 3688 81628 3728 81668
rect 3770 81628 3810 81668
rect 3852 81628 3892 81668
rect 3934 81628 3974 81668
rect 4016 81628 4056 81668
rect 5452 81208 5492 81248
rect 4928 80872 4968 80912
rect 5010 80872 5050 80912
rect 5092 80872 5132 80912
rect 5174 80872 5214 80912
rect 5256 80872 5296 80912
rect 3688 80116 3728 80156
rect 3770 80116 3810 80156
rect 3852 80116 3892 80156
rect 3934 80116 3974 80156
rect 4016 80116 4056 80156
rect 3532 79444 3572 79484
rect 4928 79360 4968 79400
rect 5010 79360 5050 79400
rect 5092 79360 5132 79400
rect 5174 79360 5214 79400
rect 5256 79360 5296 79400
rect 5356 78772 5396 78812
rect 3688 78604 3728 78644
rect 3770 78604 3810 78644
rect 3852 78604 3892 78644
rect 3934 78604 3974 78644
rect 4016 78604 4056 78644
rect 4928 77848 4968 77888
rect 5010 77848 5050 77888
rect 5092 77848 5132 77888
rect 5174 77848 5214 77888
rect 5256 77848 5296 77888
rect 3688 77092 3728 77132
rect 3770 77092 3810 77132
rect 3852 77092 3892 77132
rect 3934 77092 3974 77132
rect 4016 77092 4056 77132
rect 4300 76756 4340 76796
rect 3688 75580 3728 75620
rect 3770 75580 3810 75620
rect 3852 75580 3892 75620
rect 3934 75580 3974 75620
rect 4016 75580 4056 75620
rect 3688 74068 3728 74108
rect 3770 74068 3810 74108
rect 3852 74068 3892 74108
rect 3934 74068 3974 74108
rect 4016 74068 4056 74108
rect 3436 72388 3476 72428
rect 3916 72724 3956 72764
rect 4108 72724 4148 72764
rect 3688 72556 3728 72596
rect 3770 72556 3810 72596
rect 3852 72556 3892 72596
rect 3934 72556 3974 72596
rect 4016 72556 4056 72596
rect 3688 71044 3728 71084
rect 3770 71044 3810 71084
rect 3852 71044 3892 71084
rect 3934 71044 3974 71084
rect 4016 71044 4056 71084
rect 4012 70708 4052 70748
rect 3532 70624 3572 70664
rect 3820 70456 3860 70496
rect 3628 70288 3668 70328
rect 3688 69532 3728 69572
rect 3770 69532 3810 69572
rect 3852 69532 3892 69572
rect 3934 69532 3974 69572
rect 4016 69532 4056 69572
rect 3532 69112 3572 69152
rect 3436 69028 3476 69068
rect 3340 68692 3380 68732
rect 3916 69112 3956 69152
rect 4012 69028 4052 69068
rect 3916 68692 3956 68732
rect 4928 76336 4968 76376
rect 5010 76336 5050 76376
rect 5092 76336 5132 76376
rect 5174 76336 5214 76376
rect 5256 76336 5296 76376
rect 4928 74824 4968 74864
rect 5010 74824 5050 74864
rect 5092 74824 5132 74864
rect 5174 74824 5214 74864
rect 5256 74824 5296 74864
rect 5356 74656 5396 74696
rect 4972 74488 5012 74528
rect 5452 73816 5492 73856
rect 6316 81964 6356 82004
rect 6124 79108 6164 79148
rect 5644 74656 5684 74696
rect 5164 73564 5204 73604
rect 5452 73564 5492 73604
rect 4928 73312 4968 73352
rect 5010 73312 5050 73352
rect 5092 73312 5132 73352
rect 5174 73312 5214 73352
rect 5256 73312 5296 73352
rect 4300 70456 4340 70496
rect 4204 70288 4244 70328
rect 4396 70372 4436 70412
rect 5164 71968 5204 72008
rect 4928 71800 4968 71840
rect 5010 71800 5050 71840
rect 5092 71800 5132 71840
rect 5174 71800 5214 71840
rect 5256 71800 5296 71840
rect 5068 71548 5108 71588
rect 4588 71464 4628 71504
rect 4588 70372 4628 70412
rect 4492 70204 4532 70244
rect 4396 70120 4436 70160
rect 4492 69952 4532 69992
rect 4492 69112 4532 69152
rect 5356 71464 5396 71504
rect 5260 71380 5300 71420
rect 5164 71212 5204 71252
rect 5548 72136 5588 72176
rect 5932 73816 5972 73856
rect 6028 73648 6068 73688
rect 6700 83728 6740 83768
rect 7180 85828 7220 85868
rect 7756 84820 7796 84860
rect 7756 84484 7796 84524
rect 7564 83980 7604 84020
rect 7468 83728 7508 83768
rect 7852 83896 7892 83936
rect 6988 83476 7028 83516
rect 6412 74488 6452 74528
rect 6700 76336 6740 76376
rect 6796 75412 6836 75452
rect 6700 74656 6740 74696
rect 6604 74236 6644 74276
rect 5260 70540 5300 70580
rect 5068 70456 5108 70496
rect 4928 70288 4968 70328
rect 5010 70288 5050 70328
rect 5092 70288 5132 70328
rect 5174 70288 5214 70328
rect 5256 70288 5296 70328
rect 4972 70120 5012 70160
rect 4684 69280 4724 69320
rect 3916 68356 3956 68396
rect 3628 68188 3668 68228
rect 3688 68020 3728 68060
rect 3770 68020 3810 68060
rect 3852 68020 3892 68060
rect 3934 68020 3974 68060
rect 4016 68020 4056 68060
rect 2956 67768 2996 67808
rect 2764 67600 2804 67640
rect 2956 67516 2996 67556
rect 2188 66088 2228 66128
rect 2668 66676 2708 66716
rect 2092 58612 2132 58652
rect 3052 67432 3092 67472
rect 2956 66676 2996 66716
rect 2860 66088 2900 66128
rect 2860 65584 2900 65624
rect 2860 65416 2900 65456
rect 2668 64744 2708 64784
rect 2572 64576 2612 64616
rect 2764 64072 2804 64112
rect 2572 62728 2612 62768
rect 2476 62224 2516 62264
rect 2284 60796 2324 60836
rect 2956 63904 2996 63944
rect 2956 63064 2996 63104
rect 3532 67768 3572 67808
rect 3436 66340 3476 66380
rect 3244 66256 3284 66296
rect 4204 67600 4244 67640
rect 3688 66508 3728 66548
rect 3770 66508 3810 66548
rect 3852 66508 3892 66548
rect 3934 66508 3974 66548
rect 4016 66508 4056 66548
rect 3724 66340 3764 66380
rect 4588 68944 4628 68984
rect 4780 69112 4820 69152
rect 4972 69112 5012 69152
rect 4928 68776 4968 68816
rect 5010 68776 5050 68816
rect 5092 68776 5132 68816
rect 5174 68776 5214 68816
rect 5256 68776 5296 68816
rect 5452 70960 5492 71000
rect 5452 70708 5492 70748
rect 5356 68692 5396 68732
rect 4300 67012 4340 67052
rect 3244 66004 3284 66044
rect 3148 65500 3188 65540
rect 3628 65584 3668 65624
rect 4108 66004 4148 66044
rect 3916 65668 3956 65708
rect 3820 65500 3860 65540
rect 3724 65416 3764 65456
rect 3148 65080 3188 65120
rect 3148 64744 3188 64784
rect 3244 64240 3284 64280
rect 3148 63904 3188 63944
rect 3148 63652 3188 63692
rect 3148 63400 3188 63440
rect 3148 63064 3188 63104
rect 3052 62728 3092 62768
rect 2956 62392 2996 62432
rect 2764 61720 2804 61760
rect 2668 61552 2708 61592
rect 2572 60880 2612 60920
rect 2668 60712 2708 60752
rect 2284 59368 2324 59408
rect 2188 56008 2228 56048
rect 2284 53908 2324 53948
rect 1996 51808 2036 51848
rect 2188 53320 2228 53360
rect 2860 61552 2900 61592
rect 3052 61384 3092 61424
rect 2860 61048 2900 61088
rect 4396 66172 4436 66212
rect 4300 66088 4340 66128
rect 4204 65584 4244 65624
rect 4588 66928 4628 66968
rect 4588 66088 4628 66128
rect 4928 67264 4968 67304
rect 5010 67264 5050 67304
rect 5092 67264 5132 67304
rect 5174 67264 5214 67304
rect 5256 67264 5296 67304
rect 4972 67012 5012 67052
rect 5356 66844 5396 66884
rect 4780 66760 4820 66800
rect 5164 66172 5204 66212
rect 4396 65416 4436 65456
rect 4300 65248 4340 65288
rect 3436 65080 3476 65120
rect 3688 64996 3728 65036
rect 3770 64996 3810 65036
rect 3852 64996 3892 65036
rect 3934 64996 3974 65036
rect 4016 64996 4056 65036
rect 3820 64744 3860 64784
rect 4492 65248 4532 65288
rect 4012 64156 4052 64196
rect 3532 64072 3572 64112
rect 3436 63736 3476 63776
rect 3340 63232 3380 63272
rect 4108 64072 4148 64112
rect 4012 63820 4052 63860
rect 3916 63736 3956 63776
rect 4204 63736 4244 63776
rect 3688 63484 3728 63524
rect 3770 63484 3810 63524
rect 3852 63484 3892 63524
rect 3934 63484 3974 63524
rect 4016 63484 4056 63524
rect 3532 63400 3572 63440
rect 3916 63316 3956 63356
rect 3532 63232 3572 63272
rect 3340 63064 3380 63104
rect 3436 61636 3476 61676
rect 3340 61552 3380 61592
rect 3436 61384 3476 61424
rect 3148 60880 3188 60920
rect 3052 60040 3092 60080
rect 3244 59536 3284 59576
rect 2764 59368 2804 59408
rect 3244 59368 3284 59408
rect 2764 59116 2804 59156
rect 2668 58780 2708 58820
rect 3148 59116 3188 59156
rect 3688 61972 3728 62012
rect 3770 61972 3810 62012
rect 3852 61972 3892 62012
rect 3934 61972 3974 62012
rect 4016 61972 4056 62012
rect 3724 61636 3764 61676
rect 4204 63064 4244 63104
rect 4204 62392 4244 62432
rect 4396 64576 4436 64616
rect 4492 64324 4532 64364
rect 4780 66004 4820 66044
rect 4684 65500 4724 65540
rect 4396 63652 4436 63692
rect 4492 63316 4532 63356
rect 4588 63232 4628 63272
rect 4684 62980 4724 63020
rect 3628 60712 3668 60752
rect 3724 60628 3764 60668
rect 4108 60628 4148 60668
rect 3688 60460 3728 60500
rect 3770 60460 3810 60500
rect 3852 60460 3892 60500
rect 3934 60460 3974 60500
rect 4016 60460 4056 60500
rect 3724 59368 3764 59408
rect 3628 59116 3668 59156
rect 3688 58948 3728 58988
rect 3770 58948 3810 58988
rect 3852 58948 3892 58988
rect 3934 58948 3974 58988
rect 4016 58948 4056 58988
rect 4396 61720 4436 61760
rect 4684 61720 4724 61760
rect 4396 61048 4436 61088
rect 4204 60040 4244 60080
rect 4204 59620 4244 59660
rect 4204 59200 4244 59240
rect 4300 58780 4340 58820
rect 4108 58696 4148 58736
rect 3532 58528 3572 58568
rect 3244 58024 3284 58064
rect 3436 58024 3476 58064
rect 2572 57016 2612 57056
rect 3340 57772 3380 57812
rect 3244 57688 3284 57728
rect 2764 57268 2804 57308
rect 2860 57016 2900 57056
rect 2668 56680 2708 56720
rect 3052 56848 3092 56888
rect 3443 57604 3483 57644
rect 3340 57268 3380 57308
rect 3724 57856 3764 57896
rect 3916 57772 3956 57812
rect 4113 57688 4153 57728
rect 3628 57604 3668 57644
rect 4012 57604 4052 57644
rect 3688 57436 3728 57476
rect 3770 57436 3810 57476
rect 3852 57436 3892 57476
rect 3934 57436 3974 57476
rect 4016 57436 4056 57476
rect 3244 56848 3284 56888
rect 3436 56344 3476 56384
rect 2764 55336 2804 55376
rect 2092 50884 2132 50924
rect 1900 46768 1940 46808
rect 1996 43996 2036 44036
rect 1804 41896 1844 41936
rect 1804 41224 1844 41264
rect 1900 40384 1940 40424
rect 1708 37528 1748 37568
rect 1516 36688 1556 36728
rect 1420 34420 1460 34460
rect 1228 32740 1268 32780
rect 2668 54664 2708 54704
rect 2860 55084 2900 55124
rect 3628 56176 3668 56216
rect 3532 55924 3572 55964
rect 3688 55924 3728 55964
rect 3770 55924 3810 55964
rect 3852 55924 3892 55964
rect 3934 55924 3974 55964
rect 4016 55924 4056 55964
rect 3244 55504 3284 55544
rect 4012 55672 4052 55712
rect 3916 55504 3956 55544
rect 3340 55084 3380 55124
rect 3148 54748 3188 54788
rect 3340 54832 3380 54872
rect 3244 53656 3284 53696
rect 2572 53152 2612 53192
rect 2956 53152 2996 53192
rect 2476 51304 2516 51344
rect 2284 50716 2324 50756
rect 2860 52312 2900 52352
rect 2860 51808 2900 51848
rect 2860 51640 2900 51680
rect 2764 51052 2804 51092
rect 2860 50968 2900 51008
rect 2668 50800 2708 50840
rect 2380 50044 2420 50084
rect 2668 49372 2708 49412
rect 2284 48280 2324 48320
rect 2860 50044 2900 50084
rect 2860 49288 2900 49328
rect 2764 48700 2804 48740
rect 2476 48028 2516 48068
rect 2380 47860 2420 47900
rect 2188 47020 2228 47060
rect 2188 46600 2228 46640
rect 2476 47776 2516 47816
rect 2764 48532 2804 48572
rect 3244 53320 3284 53360
rect 3628 55336 3668 55376
rect 3688 54412 3728 54452
rect 3770 54412 3810 54452
rect 3852 54412 3892 54452
rect 3934 54412 3974 54452
rect 4016 54412 4056 54452
rect 3724 54244 3764 54284
rect 4204 55588 4244 55628
rect 3628 53908 3668 53948
rect 4300 53824 4340 53864
rect 4108 53740 4148 53780
rect 3688 52900 3728 52940
rect 3770 52900 3810 52940
rect 3852 52900 3892 52940
rect 3934 52900 3974 52940
rect 4016 52900 4056 52940
rect 3052 51724 3092 51764
rect 3244 51843 3284 51848
rect 3244 51808 3284 51843
rect 3532 52312 3572 52352
rect 3340 51640 3380 51680
rect 3340 51052 3380 51092
rect 3244 50044 3284 50084
rect 3052 48952 3092 48992
rect 2956 48364 2996 48404
rect 2572 47692 2612 47732
rect 2188 44752 2228 44792
rect 2092 42904 2132 42944
rect 2092 37696 2132 37736
rect 1996 36856 2036 36896
rect 1996 36016 2036 36056
rect 1900 34924 1940 34964
rect 1516 32404 1556 32444
rect 1324 32320 1364 32360
rect 1132 32236 1172 32276
rect 1900 32068 1940 32108
rect 1132 30808 1172 30848
rect 1804 30724 1844 30764
rect 1420 29632 1460 29672
rect 1228 28120 1268 28160
rect 1228 27616 1268 27656
rect 1324 26944 1364 26984
rect 1228 26776 1268 26816
rect 1516 27868 1556 27908
rect 2092 32740 2132 32780
rect 3724 51808 3764 51848
rect 3916 51724 3956 51764
rect 4928 65752 4968 65792
rect 5010 65752 5050 65792
rect 5092 65752 5132 65792
rect 5174 65752 5214 65792
rect 5256 65752 5296 65792
rect 5740 71464 5780 71504
rect 5644 70624 5684 70664
rect 5836 70540 5876 70580
rect 5548 70372 5588 70412
rect 5644 69280 5684 69320
rect 5548 68608 5588 68648
rect 5452 65584 5492 65624
rect 5356 65500 5396 65540
rect 5452 65416 5492 65456
rect 4928 64240 4968 64280
rect 5010 64240 5050 64280
rect 5092 64240 5132 64280
rect 5174 64240 5214 64280
rect 5256 64240 5296 64280
rect 4972 64072 5012 64112
rect 5164 63988 5204 64028
rect 5356 63316 5396 63356
rect 4928 62728 4968 62768
rect 5010 62728 5050 62768
rect 5092 62728 5132 62768
rect 5174 62728 5214 62768
rect 5256 62728 5296 62768
rect 5452 62896 5492 62936
rect 5356 61552 5396 61592
rect 4928 61216 4968 61256
rect 5010 61216 5050 61256
rect 5092 61216 5132 61256
rect 5174 61216 5214 61256
rect 5256 61216 5296 61256
rect 4780 60460 4820 60500
rect 4876 60124 4916 60164
rect 4928 59704 4968 59744
rect 5010 59704 5050 59744
rect 5092 59704 5132 59744
rect 5174 59704 5214 59744
rect 5256 59704 5296 59744
rect 4876 59452 4916 59492
rect 5452 61048 5492 61088
rect 5452 60796 5492 60836
rect 5452 59368 5492 59408
rect 5356 58948 5396 58988
rect 4780 58780 4820 58820
rect 4492 58696 4532 58736
rect 5356 58444 5396 58484
rect 4780 58276 4820 58316
rect 4684 57940 4724 57980
rect 4588 56680 4628 56720
rect 4928 58192 4968 58232
rect 5010 58192 5050 58232
rect 5092 58192 5132 58232
rect 5174 58192 5214 58232
rect 5256 58192 5296 58232
rect 4972 57688 5012 57728
rect 5260 57856 5300 57896
rect 5356 57772 5396 57812
rect 5356 57604 5396 57644
rect 4928 56680 4968 56720
rect 5010 56680 5050 56720
rect 5092 56680 5132 56720
rect 5174 56680 5214 56720
rect 5256 56680 5296 56720
rect 4492 56008 4532 56048
rect 4588 55672 4628 55712
rect 4588 54664 4628 54704
rect 5164 55924 5204 55964
rect 5356 55924 5396 55964
rect 4928 55168 4968 55208
rect 5010 55168 5050 55208
rect 5092 55168 5132 55208
rect 5174 55168 5214 55208
rect 5256 55168 5296 55208
rect 6316 71380 6356 71420
rect 6124 70960 6164 71000
rect 6028 69952 6068 69992
rect 6220 69952 6260 69992
rect 6028 69700 6068 69740
rect 5932 69280 5972 69320
rect 6412 68440 6452 68480
rect 6604 71464 6644 71504
rect 6604 71212 6644 71252
rect 6988 74236 7028 74276
rect 7372 83476 7412 83516
rect 7660 82804 7700 82844
rect 7756 75412 7796 75452
rect 7660 74488 7700 74528
rect 7660 74320 7700 74360
rect 6892 70960 6932 71000
rect 6892 70540 6932 70580
rect 6604 69112 6644 69152
rect 6220 67768 6260 67808
rect 5836 67600 5876 67640
rect 6028 67432 6068 67472
rect 6220 67096 6260 67136
rect 5836 66928 5876 66968
rect 5836 66760 5876 66800
rect 5740 66592 5780 66632
rect 5644 66424 5684 66464
rect 5740 66256 5780 66296
rect 6220 66592 6260 66632
rect 5932 65584 5972 65624
rect 5644 64492 5684 64532
rect 5740 63988 5780 64028
rect 5644 63064 5684 63104
rect 5644 61552 5684 61592
rect 6124 65416 6164 65456
rect 6124 65164 6164 65204
rect 6028 63736 6068 63776
rect 5932 62896 5972 62936
rect 6412 66508 6452 66548
rect 6316 66088 6356 66128
rect 6220 63820 6260 63860
rect 6220 62980 6260 63020
rect 5932 61552 5972 61592
rect 5836 60712 5876 60752
rect 6220 61972 6260 62012
rect 6220 60880 6260 60920
rect 6220 60040 6260 60080
rect 6028 59368 6068 59408
rect 5932 58948 5972 58988
rect 5740 58780 5780 58820
rect 5836 58696 5876 58736
rect 5932 56596 5972 56636
rect 5644 56344 5684 56384
rect 5836 56344 5876 56384
rect 5740 54664 5780 54704
rect 5548 54580 5588 54620
rect 5740 54328 5780 54368
rect 5452 54160 5492 54200
rect 4396 53740 4436 53780
rect 4684 53572 4724 53612
rect 4396 53152 4436 53192
rect 4204 52732 4244 52772
rect 4300 52648 4340 52688
rect 4204 52144 4244 52184
rect 4300 51808 4340 51848
rect 3688 51388 3728 51428
rect 3770 51388 3810 51428
rect 3852 51388 3892 51428
rect 3934 51388 3974 51428
rect 4016 51388 4056 51428
rect 3628 51220 3668 51260
rect 4012 51052 4052 51092
rect 3916 50968 3956 51008
rect 4108 50968 4148 51008
rect 3820 50296 3860 50336
rect 4012 50044 4052 50084
rect 3688 49876 3728 49916
rect 3770 49876 3810 49916
rect 3852 49876 3892 49916
rect 3934 49876 3974 49916
rect 4016 49876 4056 49916
rect 3820 49624 3860 49664
rect 3916 49540 3956 49580
rect 3340 48952 3380 48992
rect 3148 48532 3188 48572
rect 3148 48364 3188 48404
rect 2956 47776 2996 47816
rect 2860 46936 2900 46976
rect 2860 46516 2900 46556
rect 2668 46012 2708 46052
rect 2860 45928 2900 45968
rect 3052 45592 3092 45632
rect 2956 45424 2996 45464
rect 2572 44080 2612 44120
rect 2764 44080 2804 44120
rect 2476 42400 2516 42440
rect 2476 41896 2516 41936
rect 2668 42736 2708 42776
rect 2572 41476 2612 41516
rect 2572 40468 2612 40508
rect 2476 40300 2516 40340
rect 2764 41392 2804 41432
rect 2668 40048 2708 40088
rect 2860 41224 2900 41264
rect 3436 48616 3476 48656
rect 3628 48616 3668 48656
rect 3340 48028 3380 48068
rect 3244 47692 3284 47732
rect 4300 50884 4340 50924
rect 4396 50800 4436 50840
rect 4204 49624 4244 49664
rect 4108 48700 4148 48740
rect 3688 48364 3728 48404
rect 3770 48364 3810 48404
rect 3852 48364 3892 48404
rect 3934 48364 3974 48404
rect 4016 48364 4056 48404
rect 3820 48196 3860 48236
rect 3688 46852 3728 46892
rect 3770 46852 3810 46892
rect 3852 46852 3892 46892
rect 3934 46852 3974 46892
rect 4016 46852 4056 46892
rect 4300 49456 4340 49496
rect 4300 49204 4340 49244
rect 4588 52816 4628 52856
rect 4876 53824 4916 53864
rect 5932 55756 5972 55796
rect 5836 54244 5876 54284
rect 5068 53824 5108 53864
rect 5260 53824 5300 53864
rect 4928 53656 4968 53696
rect 5010 53656 5050 53696
rect 5092 53656 5132 53696
rect 5174 53656 5214 53696
rect 5256 53656 5296 53696
rect 5452 53656 5492 53696
rect 5548 53488 5588 53528
rect 5836 53656 5876 53696
rect 5452 52816 5492 52856
rect 6796 69700 6836 69740
rect 7180 72136 7220 72176
rect 7084 71716 7124 71756
rect 7180 71548 7220 71588
rect 7660 73060 7700 73100
rect 7660 72724 7700 72764
rect 7564 72136 7604 72176
rect 7372 71968 7412 72008
rect 7372 71716 7412 71756
rect 7276 71464 7316 71504
rect 7180 71212 7220 71252
rect 7276 70792 7316 70832
rect 7084 69196 7124 69236
rect 7276 70624 7316 70664
rect 7468 70540 7508 70580
rect 7180 69112 7220 69152
rect 6892 68524 6932 68564
rect 6796 68356 6836 68396
rect 6700 68020 6740 68060
rect 6604 63232 6644 63272
rect 6508 61972 6548 62012
rect 6796 67852 6836 67892
rect 6892 66424 6932 66464
rect 7084 65416 7124 65456
rect 6892 65248 6932 65288
rect 7084 64660 7124 64700
rect 6892 64324 6932 64364
rect 6796 64156 6836 64196
rect 6988 63820 7028 63860
rect 6796 62308 6836 62348
rect 6412 61720 6452 61760
rect 6700 61720 6740 61760
rect 6604 61552 6644 61592
rect 6796 61384 6836 61424
rect 7084 62980 7124 63020
rect 7372 69112 7412 69152
rect 7276 68356 7316 68396
rect 7660 71464 7700 71504
rect 7660 70540 7700 70580
rect 8140 83980 8180 84020
rect 7948 83728 7988 83768
rect 8524 85408 8564 85448
rect 8524 84652 8564 84692
rect 8428 84400 8468 84440
rect 8140 83476 8180 83516
rect 7948 83140 7988 83180
rect 8716 83896 8756 83936
rect 8716 83476 8756 83516
rect 8620 83308 8660 83348
rect 8524 83224 8564 83264
rect 8428 76840 8468 76880
rect 8524 76672 8564 76712
rect 8428 76168 8468 76208
rect 7948 76000 7988 76040
rect 8812 77428 8852 77468
rect 9004 80452 9044 80492
rect 8716 76588 8756 76628
rect 7948 74908 7988 74948
rect 7852 73900 7892 73940
rect 7852 73060 7892 73100
rect 7852 72892 7892 72932
rect 7756 69952 7796 69992
rect 7564 68440 7604 68480
rect 7468 68020 7508 68060
rect 7372 67936 7412 67976
rect 7468 67600 7508 67640
rect 7372 67432 7412 67472
rect 7468 67348 7508 67388
rect 7852 69280 7892 69320
rect 7852 68188 7892 68228
rect 7660 67600 7700 67640
rect 8140 74992 8180 75032
rect 8044 74320 8084 74360
rect 8620 74488 8660 74528
rect 8908 76840 8948 76880
rect 9292 83896 9332 83936
rect 9292 83476 9332 83516
rect 9196 83224 9236 83264
rect 9100 79192 9140 79232
rect 9100 78856 9140 78896
rect 9196 77512 9236 77552
rect 9004 76672 9044 76712
rect 8908 76168 8948 76208
rect 8908 75328 8948 75368
rect 8812 74908 8852 74948
rect 9196 76840 9236 76880
rect 9196 75328 9236 75368
rect 9196 74908 9236 74948
rect 9004 74488 9044 74528
rect 9100 74404 9140 74444
rect 8908 73816 8948 73856
rect 9004 73732 9044 73772
rect 8716 73648 8756 73688
rect 8236 73564 8276 73604
rect 8140 71968 8180 72008
rect 9100 73648 9140 73688
rect 8524 72976 8564 73016
rect 8332 72892 8372 72932
rect 8812 72892 8852 72932
rect 8332 72556 8372 72596
rect 8428 71716 8468 71756
rect 8236 70708 8276 70748
rect 8524 71380 8564 71420
rect 8716 71212 8756 71252
rect 8716 70876 8756 70916
rect 9100 71464 9140 71504
rect 9004 70708 9044 70748
rect 8236 70036 8276 70076
rect 8044 68524 8084 68564
rect 7948 67852 7988 67892
rect 8044 67600 8084 67640
rect 7276 64576 7316 64616
rect 7276 64408 7316 64448
rect 8428 69952 8468 69992
rect 8332 69196 8372 69236
rect 8236 68440 8276 68480
rect 8620 68356 8660 68396
rect 8524 66928 8564 66968
rect 8428 66844 8468 66884
rect 7564 64492 7604 64532
rect 7660 64240 7700 64280
rect 7276 64072 7316 64112
rect 7468 64072 7508 64112
rect 7180 61720 7220 61760
rect 7084 61468 7124 61508
rect 7180 61300 7220 61340
rect 6508 60796 6548 60836
rect 6700 60712 6740 60752
rect 6700 60124 6740 60164
rect 6604 60040 6644 60080
rect 6700 59872 6740 59912
rect 6412 59284 6452 59324
rect 6316 58528 6356 58568
rect 6220 58360 6260 58400
rect 6220 57436 6260 57476
rect 6220 55756 6260 55796
rect 7468 63904 7508 63944
rect 7372 63064 7412 63104
rect 7276 61048 7316 61088
rect 7276 60880 7316 60920
rect 6988 60796 7028 60836
rect 6892 60628 6932 60668
rect 6796 59200 6836 59240
rect 6700 58444 6740 58484
rect 6604 57940 6644 57980
rect 6796 56176 6836 56216
rect 6796 55672 6836 55712
rect 6604 55588 6644 55628
rect 6700 55504 6740 55544
rect 6508 55168 6548 55208
rect 6412 55000 6452 55040
rect 6124 54328 6164 54368
rect 6316 54328 6356 54368
rect 6316 53824 6356 53864
rect 6220 53572 6260 53612
rect 5932 52816 5972 52856
rect 6220 53404 6260 53444
rect 4928 52144 4968 52184
rect 5010 52144 5050 52184
rect 5092 52144 5132 52184
rect 5174 52144 5214 52184
rect 5256 52144 5296 52184
rect 5356 52144 5396 52184
rect 5452 51976 5492 52016
rect 5356 51892 5396 51932
rect 4876 51304 4916 51344
rect 4780 51052 4820 51092
rect 4684 50716 4724 50756
rect 4928 50632 4968 50672
rect 5010 50632 5050 50672
rect 5092 50632 5132 50672
rect 5174 50632 5214 50672
rect 5256 50632 5296 50672
rect 4588 49960 4628 50000
rect 4684 49288 4724 49328
rect 5452 49624 5492 49664
rect 4972 49372 5012 49412
rect 4780 49120 4820 49160
rect 4928 49120 4968 49160
rect 5010 49120 5050 49160
rect 5092 49120 5132 49160
rect 5174 49120 5214 49160
rect 5256 49120 5296 49160
rect 4876 48952 4916 48992
rect 4780 48868 4820 48908
rect 5452 48868 5492 48908
rect 5260 48784 5300 48824
rect 4588 48532 4628 48572
rect 5356 48532 5396 48572
rect 4204 48196 4244 48236
rect 4204 47860 4244 47900
rect 5356 48364 5396 48404
rect 4684 47944 4724 47984
rect 6796 55000 6836 55040
rect 6796 54664 6836 54704
rect 6604 53908 6644 53948
rect 6412 53740 6452 53780
rect 6508 53656 6548 53696
rect 6508 53320 6548 53360
rect 6412 52648 6452 52688
rect 5644 52144 5684 52184
rect 6796 54160 6836 54200
rect 6700 53824 6740 53864
rect 6604 52648 6644 52688
rect 6604 52396 6644 52436
rect 5932 51640 5972 51680
rect 5644 51556 5684 51596
rect 5932 51304 5972 51344
rect 6124 51808 6164 51848
rect 6412 51976 6452 52016
rect 7180 59872 7220 59912
rect 6988 59368 7028 59408
rect 7564 62980 7604 63020
rect 7660 62392 7700 62432
rect 7468 62308 7508 62348
rect 7564 62056 7604 62096
rect 7468 60040 7508 60080
rect 7660 61636 7700 61676
rect 7660 61468 7700 61508
rect 7660 60796 7700 60836
rect 7660 60628 7700 60668
rect 7756 60124 7796 60164
rect 7564 59872 7604 59912
rect 7180 59200 7220 59240
rect 7180 58444 7220 58484
rect 6988 56680 7028 56720
rect 7180 57268 7220 57308
rect 7180 57016 7220 57056
rect 7660 58696 7700 58736
rect 7372 58360 7412 58400
rect 7564 57940 7604 57980
rect 7564 57352 7604 57392
rect 7084 56596 7124 56636
rect 6988 56512 7028 56552
rect 6988 55168 7028 55208
rect 6988 55000 7028 55040
rect 7276 56596 7316 56636
rect 7372 56512 7412 56552
rect 7660 56848 7700 56888
rect 7276 56176 7316 56216
rect 7276 55504 7316 55544
rect 7180 55168 7220 55208
rect 7564 56176 7604 56216
rect 7468 55504 7508 55544
rect 7084 54664 7124 54704
rect 7180 54160 7220 54200
rect 7468 55000 7508 55040
rect 8716 67936 8756 67976
rect 8716 66760 8756 66800
rect 8140 66592 8180 66632
rect 7948 64408 7988 64448
rect 8044 64324 8084 64364
rect 8332 63988 8372 64028
rect 8140 63820 8180 63860
rect 7948 62476 7988 62516
rect 7852 60040 7892 60080
rect 7852 59872 7892 59912
rect 7852 59536 7892 59576
rect 7852 59284 7892 59324
rect 8044 62308 8084 62348
rect 8236 62392 8276 62432
rect 8044 61888 8084 61928
rect 8044 61384 8084 61424
rect 8044 58528 8084 58568
rect 8236 59116 8276 59156
rect 8140 58444 8180 58484
rect 7948 57940 7988 57980
rect 8140 56848 8180 56888
rect 7948 56764 7988 56804
rect 7852 56512 7892 56552
rect 7852 56344 7892 56384
rect 7756 55509 7796 55544
rect 7756 55504 7796 55509
rect 7756 55336 7796 55376
rect 7564 54916 7604 54956
rect 7372 54412 7412 54452
rect 6892 52480 6932 52520
rect 6220 51640 6260 51680
rect 6316 50884 6356 50924
rect 5740 50044 5780 50084
rect 5548 48028 5588 48068
rect 6028 50296 6068 50336
rect 6028 50044 6068 50084
rect 5836 49876 5876 49916
rect 6124 49876 6164 49916
rect 5836 49456 5876 49496
rect 6508 50380 6548 50420
rect 6316 49456 6356 49496
rect 6124 49372 6164 49412
rect 4928 47608 4968 47648
rect 5010 47608 5050 47648
rect 5092 47608 5132 47648
rect 5174 47608 5214 47648
rect 5256 47608 5296 47648
rect 4588 47272 4628 47312
rect 3532 46264 3572 46304
rect 4012 46264 4052 46304
rect 3340 46012 3380 46052
rect 3340 45844 3380 45884
rect 5644 47524 5684 47564
rect 5548 47188 5588 47228
rect 4972 46432 5012 46472
rect 5452 46600 5492 46640
rect 5068 46348 5108 46388
rect 4684 46264 4724 46304
rect 4684 45844 4724 45884
rect 4204 45424 4244 45464
rect 3688 45340 3728 45380
rect 3770 45340 3810 45380
rect 3852 45340 3892 45380
rect 3934 45340 3974 45380
rect 4016 45340 4056 45380
rect 4588 45676 4628 45716
rect 4492 45508 4532 45548
rect 4396 45256 4436 45296
rect 3916 45172 3956 45212
rect 4012 44920 4052 44960
rect 4300 44836 4340 44876
rect 4204 44752 4244 44792
rect 3244 44584 3284 44624
rect 3340 44416 3380 44456
rect 3148 44080 3188 44120
rect 3052 43408 3092 43448
rect 4108 44248 4148 44288
rect 3688 43828 3728 43868
rect 3770 43828 3810 43868
rect 3852 43828 3892 43868
rect 3934 43828 3974 43868
rect 4016 43828 4056 43868
rect 3052 42904 3092 42944
rect 3052 42064 3092 42104
rect 3244 42736 3284 42776
rect 3244 41896 3284 41936
rect 3148 41392 3188 41432
rect 3724 42652 3764 42692
rect 3628 42568 3668 42608
rect 3688 42316 3728 42356
rect 3770 42316 3810 42356
rect 3852 42316 3892 42356
rect 3934 42316 3974 42356
rect 4016 42316 4056 42356
rect 4928 46096 4968 46136
rect 5010 46096 5050 46136
rect 5092 46096 5132 46136
rect 5174 46096 5214 46136
rect 5256 46096 5296 46136
rect 5356 46012 5396 46052
rect 5068 45928 5108 45968
rect 4972 45592 5012 45632
rect 4972 45340 5012 45380
rect 4972 45088 5012 45128
rect 4780 44920 4820 44960
rect 4396 44584 4436 44624
rect 4928 44584 4968 44624
rect 5010 44584 5050 44624
rect 5092 44584 5132 44624
rect 5174 44584 5214 44624
rect 5256 44584 5296 44624
rect 4588 44416 4628 44456
rect 4204 42820 4244 42860
rect 4300 42736 4340 42776
rect 3916 42148 3956 42188
rect 3724 42064 3764 42104
rect 3820 41560 3860 41600
rect 3724 41224 3764 41264
rect 2284 39628 2324 39668
rect 2188 32152 2228 32192
rect 2092 31312 2132 31352
rect 1996 30052 2036 30092
rect 1996 29884 2036 29924
rect 1420 26272 1460 26312
rect 1228 26188 1268 26228
rect 1324 26104 1364 26144
rect 1516 25852 1556 25892
rect 1132 24676 1172 24716
rect 1324 25096 1364 25136
rect 1420 24928 1460 24968
rect 1612 25264 1652 25304
rect 1228 24592 1268 24632
rect 1996 27868 2036 27908
rect 1996 26776 2036 26816
rect 1996 26356 2036 26396
rect 1900 26188 1940 26228
rect 2188 29800 2228 29840
rect 2668 39712 2708 39752
rect 2572 38536 2612 38576
rect 3148 40300 3188 40340
rect 3148 40048 3188 40088
rect 2956 38872 2996 38912
rect 3052 38704 3092 38744
rect 3052 38536 3092 38576
rect 2380 37360 2420 37400
rect 2476 36940 2516 36980
rect 2668 36856 2708 36896
rect 2476 35932 2516 35972
rect 2668 35176 2708 35216
rect 3148 36184 3188 36224
rect 3052 35260 3092 35300
rect 3052 35092 3092 35132
rect 3148 35008 3188 35048
rect 3052 34336 3092 34376
rect 2764 34168 2804 34208
rect 4204 41896 4244 41936
rect 4876 44248 4916 44288
rect 4876 43408 4916 43448
rect 4928 43072 4968 43112
rect 5010 43072 5050 43112
rect 5092 43072 5132 43112
rect 5174 43072 5214 43112
rect 5256 43072 5296 43112
rect 5356 42904 5396 42944
rect 4492 42736 4532 42776
rect 4396 42652 4436 42692
rect 4492 42568 4532 42608
rect 4396 41980 4436 42020
rect 4108 41560 4148 41600
rect 4300 41560 4340 41600
rect 4012 40972 4052 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 3340 40552 3380 40592
rect 3532 40468 3572 40508
rect 3820 39712 3860 39752
rect 4204 41056 4244 41096
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 4684 42148 4724 42188
rect 4780 41980 4820 42020
rect 5260 42820 5300 42860
rect 5068 42736 5108 42776
rect 5164 42484 5204 42524
rect 5356 42652 5396 42692
rect 5356 42400 5396 42440
rect 5356 42064 5396 42104
rect 5068 41728 5108 41768
rect 4492 41056 4532 41096
rect 4300 39628 4340 39668
rect 4204 39208 4244 39248
rect 4108 39040 4148 39080
rect 3340 38872 3380 38912
rect 3532 38704 3572 38744
rect 3340 38200 3380 38240
rect 3628 38116 3668 38156
rect 4012 38032 4052 38072
rect 4108 37948 4148 37988
rect 3436 37024 3476 37064
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3724 37360 3764 37400
rect 4108 37192 4148 37232
rect 3628 37024 3668 37064
rect 3340 36604 3380 36644
rect 3340 36352 3380 36392
rect 3340 35932 3380 35972
rect 3244 34084 3284 34124
rect 3052 33916 3092 33956
rect 2956 33832 2996 33872
rect 2956 33664 2996 33704
rect 2668 33412 2708 33452
rect 2860 32824 2900 32864
rect 3244 33832 3284 33872
rect 3532 36856 3572 36896
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 3724 36100 3764 36140
rect 4012 36100 4052 36140
rect 3436 35092 3476 35132
rect 3628 35176 3668 35216
rect 3532 35008 3572 35048
rect 4492 37948 4532 37988
rect 5260 41728 5300 41768
rect 4780 41560 4820 41600
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 5548 42232 5588 42272
rect 5740 47356 5780 47396
rect 5836 46180 5876 46220
rect 6220 49036 6260 49076
rect 6316 48868 6356 48908
rect 6220 48784 6260 48824
rect 6124 47776 6164 47816
rect 6124 47272 6164 47312
rect 6508 49204 6548 49244
rect 6508 48784 6548 48824
rect 6412 47608 6452 47648
rect 6316 46852 6356 46892
rect 6220 46516 6260 46556
rect 6412 46432 6452 46472
rect 6316 46012 6356 46052
rect 6220 45844 6260 45884
rect 5836 45592 5876 45632
rect 6028 45676 6068 45716
rect 5932 45340 5972 45380
rect 5740 42820 5780 42860
rect 5836 42736 5876 42776
rect 5740 42484 5780 42524
rect 5644 41560 5684 41600
rect 5740 41392 5780 41432
rect 5164 40972 5204 41012
rect 4780 40720 4820 40760
rect 5356 40552 5396 40592
rect 5164 40384 5204 40424
rect 4972 40300 5012 40340
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 5164 39712 5204 39752
rect 4684 38956 4724 38996
rect 5164 38872 5204 38912
rect 5356 38872 5396 38912
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 5644 40384 5684 40424
rect 5452 38368 5492 38408
rect 5452 38116 5492 38156
rect 4012 35176 4052 35216
rect 3724 34924 3764 34964
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 3436 33748 3476 33788
rect 3916 33664 3956 33704
rect 4588 37360 4628 37400
rect 5356 37360 5396 37400
rect 5260 37192 5300 37232
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 4876 36520 4916 36560
rect 4300 34420 4340 34460
rect 4300 34084 4340 34124
rect 4204 33916 4244 33956
rect 4492 35008 4532 35048
rect 4588 34336 4628 34376
rect 4492 34252 4532 34292
rect 4492 34000 4532 34040
rect 4396 33832 4436 33872
rect 4204 33664 4244 33704
rect 4108 33412 4148 33452
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 4396 33580 4436 33620
rect 4492 33412 4532 33452
rect 4396 33244 4436 33284
rect 3340 32992 3380 33032
rect 2860 32152 2900 32192
rect 2476 32068 2516 32108
rect 2764 32068 2804 32108
rect 2476 31900 2516 31940
rect 2380 31312 2420 31352
rect 2476 30640 2516 30680
rect 2668 30052 2708 30092
rect 2668 29380 2708 29420
rect 2284 29296 2324 29336
rect 2188 29128 2228 29168
rect 2284 29044 2324 29084
rect 2380 28792 2420 28832
rect 2284 26440 2324 26480
rect 2188 25348 2228 25388
rect 1900 25096 1940 25136
rect 1324 23164 1364 23204
rect 1324 22240 1364 22280
rect 1516 21568 1556 21608
rect 1516 20896 1556 20936
rect 1420 20056 1460 20096
rect 1324 19048 1364 19088
rect 1132 18292 1172 18332
rect 1324 17200 1364 17240
rect 1804 23836 1844 23876
rect 1996 24424 2036 24464
rect 1996 23836 2036 23876
rect 1900 23668 1940 23708
rect 2092 23584 2132 23624
rect 1996 23500 2036 23540
rect 1708 20308 1748 20348
rect 1708 19720 1748 19760
rect 1612 18292 1652 18332
rect 1516 17956 1556 17996
rect 1804 18292 1844 18332
rect 1900 17757 1940 17786
rect 1900 17746 1940 17757
rect 1804 17368 1844 17408
rect 1708 16192 1748 16232
rect 1612 15772 1652 15812
rect 1324 14680 1364 14720
rect 1228 14512 1268 14552
rect 1036 13672 1076 13712
rect 1516 13252 1556 13292
rect 1420 12496 1460 12536
rect 460 11320 500 11360
rect 1516 11824 1556 11864
rect 1324 11488 1364 11528
rect 1516 11404 1556 11444
rect 1228 11152 1268 11192
rect 1324 10984 1364 11024
rect 2188 20728 2228 20768
rect 2092 18460 2132 18500
rect 2188 17956 2228 17996
rect 2188 17788 2228 17828
rect 2188 17368 2228 17408
rect 2092 17200 2132 17240
rect 1996 15940 2036 15980
rect 1900 15772 1940 15812
rect 1996 15688 2036 15728
rect 1900 15520 1940 15560
rect 1804 14176 1844 14216
rect 1708 13168 1748 13208
rect 1708 12916 1748 12956
rect 1804 12748 1844 12788
rect 1996 13168 2036 13208
rect 1996 12496 2036 12536
rect 2572 26692 2612 26732
rect 2380 23500 2420 23540
rect 2476 22324 2516 22364
rect 2668 25264 2708 25304
rect 3148 32656 3188 32696
rect 2860 31060 2900 31100
rect 3532 32488 3572 32528
rect 3820 32824 3860 32864
rect 4108 32824 4148 32864
rect 5740 39712 5780 39752
rect 5740 39040 5780 39080
rect 5644 38872 5684 38912
rect 6124 44248 6164 44288
rect 6412 45844 6452 45884
rect 6604 47860 6644 47900
rect 6892 50632 6932 50672
rect 6892 49372 6932 49412
rect 7276 53992 7316 54032
rect 7276 53236 7316 53276
rect 7180 52648 7220 52688
rect 7084 52564 7124 52604
rect 7084 52396 7124 52436
rect 7180 51976 7220 52016
rect 7180 51808 7220 51848
rect 7564 54160 7604 54200
rect 7564 53572 7604 53612
rect 7468 53488 7508 53528
rect 7084 51304 7124 51344
rect 7084 50548 7124 50588
rect 7084 49708 7124 49748
rect 7372 51640 7412 51680
rect 7948 56092 7988 56132
rect 8524 66340 8564 66380
rect 8524 65500 8564 65540
rect 8524 64660 8564 64700
rect 8716 64660 8756 64700
rect 8620 64492 8660 64532
rect 8524 64072 8564 64112
rect 8524 63820 8564 63860
rect 8428 63484 8468 63524
rect 8620 63064 8660 63104
rect 8428 61552 8468 61592
rect 8428 61384 8468 61424
rect 9388 83140 9428 83180
rect 9292 71464 9332 71504
rect 9580 83896 9620 83936
rect 9580 79528 9620 79568
rect 9484 76672 9524 76712
rect 9580 75580 9620 75620
rect 9484 74488 9524 74528
rect 10060 84400 10100 84440
rect 10156 82300 10196 82340
rect 9772 79192 9812 79232
rect 9676 73732 9716 73772
rect 9580 73648 9620 73688
rect 9676 71548 9716 71588
rect 9196 70624 9236 70664
rect 9004 70456 9044 70496
rect 8908 70372 8948 70412
rect 9580 70708 9620 70748
rect 9676 70624 9716 70664
rect 9196 69112 9236 69152
rect 9004 68272 9044 68312
rect 9100 67852 9140 67892
rect 9100 67684 9140 67724
rect 9100 66088 9140 66128
rect 9100 65332 9140 65372
rect 8812 63232 8852 63272
rect 9100 63652 9140 63692
rect 9100 63232 9140 63272
rect 9004 63148 9044 63188
rect 8812 62728 8852 62768
rect 8620 62392 8660 62432
rect 8908 61720 8948 61760
rect 9484 68440 9524 68480
rect 9484 67684 9524 67724
rect 9388 66088 9428 66128
rect 9292 64408 9332 64448
rect 9292 62644 9332 62684
rect 9004 60796 9044 60836
rect 9004 60628 9044 60668
rect 8524 60544 8564 60584
rect 9196 60208 9236 60248
rect 8812 59200 8852 59240
rect 8620 59116 8660 59156
rect 9100 58948 9140 58988
rect 9100 57856 9140 57896
rect 8620 57100 8660 57140
rect 8812 57016 8852 57056
rect 8428 56848 8468 56888
rect 8236 56344 8276 56384
rect 8428 56176 8468 56216
rect 8140 55756 8180 55796
rect 8332 55672 8372 55712
rect 9100 56764 9140 56804
rect 8908 56344 8948 56384
rect 8620 55756 8660 55796
rect 9100 55672 9140 55712
rect 8620 55588 8660 55628
rect 9004 54832 9044 54872
rect 8332 54748 8372 54788
rect 8140 54664 8180 54704
rect 7852 54244 7892 54284
rect 7756 53572 7796 53612
rect 7660 53404 7700 53444
rect 7756 53320 7796 53360
rect 7948 53992 7988 54032
rect 7948 53236 7988 53276
rect 7564 51220 7604 51260
rect 7756 52648 7796 52688
rect 7756 52060 7796 52100
rect 7852 51556 7892 51596
rect 9004 54412 9044 54452
rect 8620 54160 8660 54200
rect 8524 53992 8564 54032
rect 8428 53824 8468 53864
rect 8236 53320 8276 53360
rect 8140 52900 8180 52940
rect 8044 52816 8084 52856
rect 8044 52564 8084 52604
rect 7948 51304 7988 51344
rect 8332 53068 8372 53108
rect 8332 52732 8372 52772
rect 8236 52312 8276 52352
rect 8044 51220 8084 51260
rect 7660 51136 7700 51176
rect 8332 51808 8372 51848
rect 7468 50968 7508 51008
rect 7468 50548 7508 50588
rect 7756 50884 7796 50924
rect 8044 50884 8084 50924
rect 8332 50884 8372 50924
rect 8236 50800 8276 50840
rect 7660 50632 7700 50672
rect 8236 50464 8276 50504
rect 7948 50380 7988 50420
rect 7660 50251 7700 50252
rect 7660 50212 7700 50251
rect 7660 49624 7700 49664
rect 7468 49288 7508 49328
rect 6988 48868 7028 48908
rect 6796 48784 6836 48824
rect 7276 48819 7316 48824
rect 7276 48784 7316 48819
rect 7564 48700 7604 48740
rect 7468 48616 7508 48656
rect 7468 48364 7508 48404
rect 6988 48196 7028 48236
rect 6796 48028 6836 48068
rect 6892 47944 6932 47984
rect 7084 48028 7124 48068
rect 6700 47272 6740 47312
rect 7276 47944 7316 47984
rect 7660 48616 7700 48656
rect 7564 48028 7604 48068
rect 7660 47944 7700 47984
rect 8236 49792 8276 49832
rect 7852 49708 7892 49748
rect 8524 53488 8564 53528
rect 9100 54076 9140 54116
rect 8716 53992 8756 54032
rect 9004 53992 9044 54032
rect 8908 53572 8948 53612
rect 8620 53320 8660 53360
rect 8620 53068 8660 53108
rect 8524 51556 8564 51596
rect 8716 52480 8756 52520
rect 8620 51304 8660 51344
rect 8620 51136 8660 51176
rect 8620 49960 8660 50000
rect 8428 49624 8468 49664
rect 7948 48784 7988 48824
rect 8428 49456 8468 49496
rect 8236 48616 8276 48656
rect 8044 48532 8084 48572
rect 8620 48532 8660 48572
rect 8140 48028 8180 48068
rect 6988 47272 7028 47312
rect 6700 46684 6740 46724
rect 6604 46516 6644 46556
rect 7564 46684 7604 46724
rect 7084 46600 7124 46640
rect 7276 46516 7316 46556
rect 6604 46348 6644 46388
rect 7180 46432 7220 46472
rect 6796 46264 6836 46304
rect 6604 46198 6644 46220
rect 6604 46180 6644 46198
rect 6988 46096 7028 46136
rect 6316 45592 6356 45632
rect 6700 45592 6740 45632
rect 6412 45508 6452 45548
rect 6508 44920 6548 44960
rect 6508 44248 6548 44288
rect 6988 45508 7028 45548
rect 6892 45424 6932 45464
rect 6796 44920 6836 44960
rect 8716 47272 8756 47312
rect 8812 46852 8852 46892
rect 8620 46684 8660 46724
rect 8140 46600 8180 46640
rect 8236 46516 8276 46556
rect 7852 46432 7892 46472
rect 7756 46348 7796 46388
rect 7180 45508 7220 45548
rect 7372 45508 7412 45548
rect 7276 45172 7316 45212
rect 7564 45760 7604 45800
rect 7756 45760 7796 45800
rect 7948 45760 7988 45800
rect 7468 45088 7508 45128
rect 7756 44920 7796 44960
rect 8428 46264 8468 46304
rect 8524 45760 8564 45800
rect 8236 45592 8276 45632
rect 8140 45088 8180 45128
rect 8332 45088 8372 45128
rect 8236 44920 8276 44960
rect 7852 44752 7892 44792
rect 8044 44752 8084 44792
rect 7468 44668 7508 44708
rect 6892 44332 6932 44372
rect 6892 44164 6932 44204
rect 6796 44080 6836 44120
rect 6508 43492 6548 43532
rect 6220 43408 6260 43448
rect 5932 41560 5972 41600
rect 5836 38116 5876 38156
rect 5548 37612 5588 37652
rect 5740 37108 5780 37148
rect 5548 36940 5588 36980
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 5068 34924 5108 34964
rect 5260 34672 5300 34712
rect 5260 34420 5300 34460
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 5452 34840 5492 34880
rect 5548 34168 5588 34208
rect 5452 33916 5492 33956
rect 5164 33748 5204 33788
rect 4876 33496 4916 33536
rect 6028 40384 6068 40424
rect 6604 42736 6644 42776
rect 6604 42484 6644 42524
rect 6700 42316 6740 42356
rect 6316 41560 6356 41600
rect 6700 41560 6740 41600
rect 6220 41392 6260 41432
rect 6892 41560 6932 41600
rect 6796 41476 6836 41516
rect 6412 40888 6452 40928
rect 6124 40132 6164 40172
rect 6796 40636 6836 40676
rect 6700 40384 6740 40424
rect 6316 40300 6356 40340
rect 6604 40300 6644 40340
rect 6124 39460 6164 39500
rect 6028 39040 6068 39080
rect 6028 38704 6068 38744
rect 5932 37696 5972 37736
rect 5836 35344 5876 35384
rect 5932 34840 5972 34880
rect 6508 39628 6548 39668
rect 7084 44248 7124 44288
rect 6988 39796 7028 39836
rect 6316 39040 6356 39080
rect 6700 38536 6740 38576
rect 6604 38368 6644 38408
rect 6316 38200 6356 38240
rect 6508 37864 6548 37904
rect 6220 37612 6260 37652
rect 6508 36940 6548 36980
rect 6124 36604 6164 36644
rect 6892 39124 6932 39164
rect 6988 39040 7028 39080
rect 6700 38032 6740 38072
rect 6988 37360 7028 37400
rect 6796 36856 6836 36896
rect 7468 44080 7508 44120
rect 8140 44248 8180 44288
rect 8332 44500 8372 44540
rect 8332 44080 8372 44120
rect 8236 43996 8276 44036
rect 8716 45508 8756 45548
rect 8620 45088 8660 45128
rect 8620 44836 8660 44876
rect 8524 43828 8564 43868
rect 8140 43492 8180 43532
rect 8044 43324 8084 43364
rect 7372 42988 7412 43028
rect 7276 40552 7316 40592
rect 8716 43996 8756 44036
rect 8812 43744 8852 43784
rect 8140 41812 8180 41852
rect 8044 41560 8084 41600
rect 7660 41476 7700 41516
rect 7564 40972 7604 41012
rect 7564 40720 7604 40760
rect 7372 39460 7412 39500
rect 7180 39040 7220 39080
rect 7468 39208 7508 39248
rect 8236 41308 8276 41348
rect 8812 41812 8852 41852
rect 8620 41560 8660 41600
rect 8620 41224 8660 41264
rect 8044 40888 8084 40928
rect 7660 40468 7700 40508
rect 7564 39124 7604 39164
rect 7468 38956 7508 38996
rect 7276 38368 7316 38408
rect 7276 37948 7316 37988
rect 7180 37612 7220 37652
rect 6796 36688 6836 36728
rect 7084 36688 7124 36728
rect 6988 36520 7028 36560
rect 7180 36100 7220 36140
rect 6220 35260 6260 35300
rect 6124 34588 6164 34628
rect 5740 34504 5780 34544
rect 6028 34504 6068 34544
rect 6124 34420 6164 34460
rect 5740 34336 5780 34376
rect 5644 34000 5684 34040
rect 5932 33916 5972 33956
rect 5452 33412 5492 33452
rect 5356 33328 5396 33368
rect 4972 33244 5012 33284
rect 4876 33076 4916 33116
rect 4684 32908 4724 32948
rect 6124 33748 6164 33788
rect 5932 33496 5972 33536
rect 3532 32152 3572 32192
rect 3244 32068 3284 32108
rect 3436 30724 3476 30764
rect 3340 30640 3380 30680
rect 3148 29968 3188 30008
rect 3148 29800 3188 29840
rect 4492 32152 4532 32192
rect 4588 32068 4628 32108
rect 5644 32572 5684 32612
rect 6028 32572 6068 32612
rect 4780 32488 4820 32528
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 4780 31900 4820 31940
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 4684 31648 4724 31688
rect 4588 31564 4628 31604
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 4108 29968 4148 30008
rect 3052 29044 3092 29084
rect 2956 28876 2996 28916
rect 2860 27952 2900 27992
rect 3148 28456 3188 28496
rect 3340 29044 3380 29084
rect 3244 27952 3284 27992
rect 3148 27784 3188 27824
rect 2956 27616 2996 27656
rect 2956 27448 2996 27488
rect 2860 26692 2900 26732
rect 2860 26020 2900 26060
rect 2860 25348 2900 25388
rect 2860 25180 2900 25220
rect 2764 23752 2804 23792
rect 3148 27532 3188 27572
rect 3052 26608 3092 26648
rect 3340 27448 3380 27488
rect 3628 29632 3668 29672
rect 3820 29800 3860 29840
rect 3820 29464 3860 29504
rect 3724 29296 3764 29336
rect 4108 29632 4148 29672
rect 4012 29548 4052 29588
rect 3916 29128 3956 29168
rect 3724 28876 3764 28916
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 4108 28456 4148 28496
rect 3532 28372 3572 28412
rect 3628 28288 3668 28328
rect 4108 28288 4148 28328
rect 3628 27700 3668 27740
rect 3532 27616 3572 27656
rect 4108 27616 4148 27656
rect 3532 27364 3572 27404
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 3244 26692 3284 26732
rect 3148 26356 3188 26396
rect 3148 26104 3188 26144
rect 3244 26020 3284 26060
rect 3244 25852 3284 25892
rect 3148 25348 3188 25388
rect 3052 24760 3092 24800
rect 3052 24004 3092 24044
rect 3244 25180 3284 25220
rect 3628 26944 3668 26984
rect 3628 26608 3668 26648
rect 3436 26272 3476 26312
rect 3820 26356 3860 26396
rect 3532 25936 3572 25976
rect 3436 25264 3476 25304
rect 3820 25852 3860 25892
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 4012 25516 4052 25556
rect 4492 30892 4532 30932
rect 4396 30640 4436 30680
rect 4588 29800 4628 29840
rect 4396 29548 4436 29588
rect 5068 31312 5108 31352
rect 5164 31228 5204 31268
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 4780 30640 4820 30680
rect 5068 30640 5108 30680
rect 5452 31480 5492 31520
rect 5932 31480 5972 31520
rect 5644 31144 5684 31184
rect 5452 30976 5492 31016
rect 5356 30472 5396 30512
rect 5164 30388 5204 30428
rect 4780 30220 4820 30260
rect 5548 30556 5588 30596
rect 5644 30472 5684 30512
rect 5740 30388 5780 30428
rect 5452 29884 5492 29924
rect 5356 29800 5396 29840
rect 4684 29632 4724 29672
rect 4588 29464 4628 29504
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 5356 29464 5396 29504
rect 4300 28624 4340 28664
rect 4300 28456 4340 28496
rect 4204 26272 4244 26312
rect 4108 24928 4148 24968
rect 3532 24844 3572 24884
rect 3916 24627 3956 24632
rect 3916 24592 3956 24627
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 3628 24004 3668 24044
rect 3148 23752 3188 23792
rect 2668 22576 2708 22616
rect 3148 23080 3188 23120
rect 3052 22492 3092 22532
rect 2860 22408 2900 22448
rect 2668 22324 2708 22364
rect 2956 21736 2996 21776
rect 2668 21484 2708 21524
rect 2860 21484 2900 21524
rect 2572 20476 2612 20516
rect 2668 20140 2708 20180
rect 2572 19300 2612 19340
rect 2476 18628 2516 18668
rect 2476 17956 2516 17996
rect 2476 17620 2516 17660
rect 3148 21988 3188 22028
rect 2860 20560 2900 20600
rect 3052 20140 3092 20180
rect 3052 18124 3092 18164
rect 3532 23752 3572 23792
rect 4012 23752 4052 23792
rect 3916 23668 3956 23708
rect 3340 23500 3380 23540
rect 3436 23248 3476 23288
rect 4972 29296 5012 29336
rect 5164 29296 5204 29336
rect 4485 29044 4525 29084
rect 4588 28960 4628 29000
rect 5164 29128 5204 29168
rect 5548 29800 5588 29840
rect 5068 29044 5108 29084
rect 4492 28624 4532 28664
rect 4396 27028 4436 27068
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4588 27784 4628 27824
rect 5644 29044 5684 29084
rect 5836 29800 5876 29840
rect 6412 34504 6452 34544
rect 6412 34168 6452 34208
rect 6124 32152 6164 32192
rect 6412 33496 6452 33536
rect 7372 37108 7412 37148
rect 7372 36184 7412 36224
rect 7372 36016 7412 36056
rect 6700 35176 6740 35216
rect 6988 35344 7028 35384
rect 6892 34756 6932 34796
rect 6796 34588 6836 34628
rect 6700 34504 6740 34544
rect 6604 34336 6644 34376
rect 6700 34252 6740 34292
rect 6028 30220 6068 30260
rect 6220 30136 6260 30176
rect 6892 34168 6932 34208
rect 6892 33664 6932 33704
rect 7372 35596 7412 35636
rect 6796 32908 6836 32948
rect 6700 31480 6740 31520
rect 7372 35211 7412 35216
rect 7372 35176 7412 35211
rect 7372 34504 7412 34544
rect 7564 38200 7604 38240
rect 8812 40720 8852 40760
rect 8236 40636 8276 40676
rect 8044 40384 8084 40424
rect 8620 40384 8660 40424
rect 8428 40216 8468 40256
rect 8140 39796 8180 39836
rect 7948 39040 7988 39080
rect 8812 39544 8852 39584
rect 8812 39040 8852 39080
rect 8620 38956 8660 38996
rect 7660 37696 7700 37736
rect 7756 37612 7796 37652
rect 8140 38200 8180 38240
rect 8140 37948 8180 37988
rect 7948 37444 7988 37484
rect 9004 53488 9044 53528
rect 9004 53068 9044 53108
rect 9100 52396 9140 52436
rect 9484 65584 9524 65624
rect 9868 77512 9908 77552
rect 10060 77512 10100 77552
rect 10348 83644 10388 83684
rect 10636 84400 10676 84440
rect 10444 83140 10484 83180
rect 10540 79108 10580 79148
rect 10732 79360 10772 79400
rect 10924 83392 10964 83432
rect 10828 79276 10868 79316
rect 10828 79108 10868 79148
rect 11020 82300 11060 82340
rect 11404 83812 11444 83852
rect 11020 79696 11060 79736
rect 11020 79108 11060 79148
rect 10924 79024 10964 79064
rect 10732 78100 10772 78140
rect 10348 78016 10388 78056
rect 10252 77596 10292 77636
rect 10348 77512 10388 77552
rect 10924 77596 10964 77636
rect 9964 76840 10004 76880
rect 10156 76504 10196 76544
rect 9964 76000 10004 76040
rect 10156 76000 10196 76040
rect 10348 76924 10388 76964
rect 10444 76252 10484 76292
rect 10348 75832 10388 75872
rect 10252 75580 10292 75620
rect 10156 75160 10196 75200
rect 10060 74992 10100 75032
rect 10252 74740 10292 74780
rect 10060 73060 10100 73100
rect 10156 72808 10196 72848
rect 9964 72388 10004 72428
rect 10444 75160 10484 75200
rect 10348 73144 10388 73184
rect 10732 76504 10772 76544
rect 10636 75664 10676 75704
rect 10636 74992 10676 75032
rect 10636 74656 10676 74696
rect 10348 72976 10388 73016
rect 10348 72640 10388 72680
rect 11020 76924 11060 76964
rect 10924 76504 10964 76544
rect 11020 75832 11060 75872
rect 10924 75328 10964 75368
rect 10828 74404 10868 74444
rect 10636 72640 10676 72680
rect 10348 71800 10388 71840
rect 10732 71548 10772 71588
rect 10540 70876 10580 70916
rect 9772 69028 9812 69068
rect 10060 69196 10100 69236
rect 10156 68944 10196 68984
rect 9676 68440 9716 68480
rect 9964 68440 10004 68480
rect 9868 68356 9908 68396
rect 9772 67852 9812 67892
rect 9772 67600 9812 67640
rect 9772 64576 9812 64616
rect 10060 67768 10100 67808
rect 10348 68944 10388 68984
rect 10252 68440 10292 68480
rect 10540 70120 10580 70160
rect 10444 67936 10484 67976
rect 10156 66928 10196 66968
rect 10732 69868 10772 69908
rect 10636 69196 10676 69236
rect 10732 69112 10772 69152
rect 10636 68944 10676 68984
rect 10732 68440 10772 68480
rect 10924 72976 10964 73016
rect 11212 81796 11252 81836
rect 11308 79948 11348 79988
rect 11404 79360 11444 79400
rect 11308 79108 11348 79148
rect 11308 78940 11348 78980
rect 11212 76420 11252 76460
rect 11116 73648 11156 73688
rect 11020 72892 11060 72932
rect 11020 72640 11060 72680
rect 11116 71548 11156 71588
rect 10924 69868 10964 69908
rect 10924 68440 10964 68480
rect 10828 67936 10868 67976
rect 10540 67768 10580 67808
rect 9484 61720 9524 61760
rect 9772 61720 9812 61760
rect 9772 61132 9812 61172
rect 9388 59704 9428 59744
rect 9676 59620 9716 59660
rect 9964 64324 10004 64364
rect 10060 63820 10100 63860
rect 10060 63400 10100 63440
rect 10060 63064 10100 63104
rect 9964 61552 10004 61592
rect 10060 60880 10100 60920
rect 9868 59872 9908 59912
rect 9292 58864 9332 58904
rect 9388 58696 9428 58736
rect 9964 59704 10004 59744
rect 10732 66424 10772 66464
rect 10924 67600 10964 67640
rect 10828 66340 10868 66380
rect 10348 66088 10388 66128
rect 10252 65500 10292 65540
rect 10444 65668 10484 65708
rect 10348 65248 10388 65288
rect 10540 65164 10580 65204
rect 10828 64576 10868 64616
rect 11212 70120 11252 70160
rect 11116 69280 11156 69320
rect 12172 84400 12212 84440
rect 11980 83224 12020 83264
rect 12748 81964 12788 82004
rect 11404 76672 11444 76712
rect 11692 79108 11732 79148
rect 11980 79780 12020 79820
rect 12268 79780 12308 79820
rect 11500 76000 11540 76040
rect 12172 79696 12212 79736
rect 11980 78016 12020 78056
rect 12940 81208 12980 81248
rect 12748 79360 12788 79400
rect 12172 76504 12212 76544
rect 11884 76252 11924 76292
rect 12172 76252 12212 76292
rect 11980 76168 12020 76208
rect 11692 75832 11732 75872
rect 11596 75160 11636 75200
rect 11404 74992 11444 75032
rect 11500 74656 11540 74696
rect 11500 73396 11540 73436
rect 11404 72976 11444 73016
rect 11212 68440 11252 68480
rect 11212 67516 11252 67556
rect 11596 72388 11636 72428
rect 11596 71968 11636 72008
rect 11884 74320 11924 74360
rect 11788 73984 11828 74024
rect 12076 75160 12116 75200
rect 12076 74656 12116 74696
rect 11980 74236 12020 74276
rect 11980 73816 12020 73856
rect 12268 76168 12308 76208
rect 12268 74488 12308 74528
rect 12268 74236 12308 74276
rect 11980 73564 12020 73604
rect 11788 73396 11828 73436
rect 11788 72724 11828 72764
rect 12076 72808 12116 72848
rect 11596 70624 11636 70664
rect 11980 71128 12020 71168
rect 11980 70960 12020 71000
rect 11884 69112 11924 69152
rect 11692 68272 11732 68312
rect 11596 68104 11636 68144
rect 11788 67768 11828 67808
rect 11116 65500 11156 65540
rect 11020 64660 11060 64700
rect 11500 66172 11540 66212
rect 11308 65500 11348 65540
rect 11404 65416 11444 65456
rect 11308 65164 11348 65204
rect 11212 64324 11252 64364
rect 10348 63820 10388 63860
rect 10540 63736 10580 63776
rect 10444 63652 10484 63692
rect 10636 63484 10676 63524
rect 10252 63064 10292 63104
rect 10252 61720 10292 61760
rect 10540 63148 10580 63188
rect 11020 63988 11060 64028
rect 10828 63652 10868 63692
rect 11020 63736 11060 63776
rect 10732 63148 10772 63188
rect 10732 62980 10772 63020
rect 10444 61804 10484 61844
rect 10348 61636 10388 61676
rect 10252 61300 10292 61340
rect 10540 61720 10580 61760
rect 10540 61300 10580 61340
rect 10540 61048 10580 61088
rect 10540 60796 10580 60836
rect 10348 60544 10388 60584
rect 10252 59620 10292 59660
rect 10060 59200 10100 59240
rect 9964 58864 10004 58904
rect 9868 58696 9908 58736
rect 9964 58528 10004 58568
rect 10156 58444 10196 58484
rect 9868 57940 9908 57980
rect 9484 56764 9524 56804
rect 9676 56344 9716 56384
rect 9484 56260 9524 56300
rect 9292 56092 9332 56132
rect 9676 55252 9716 55292
rect 9292 53488 9332 53528
rect 9676 54748 9716 54788
rect 9484 54496 9524 54536
rect 9676 54160 9716 54200
rect 9580 54076 9620 54116
rect 9388 53320 9428 53360
rect 9676 53992 9716 54032
rect 9580 53740 9620 53780
rect 9196 51640 9236 51680
rect 9676 53068 9716 53108
rect 10060 57100 10100 57140
rect 9868 56092 9908 56132
rect 10060 55672 10100 55712
rect 10444 60040 10484 60080
rect 10348 58780 10388 58820
rect 10444 58444 10484 58484
rect 10348 55672 10388 55712
rect 10252 55504 10292 55544
rect 9868 55000 9908 55040
rect 10156 54916 10196 54956
rect 10252 54832 10292 54872
rect 10156 54664 10196 54704
rect 10060 54244 10100 54284
rect 10060 53992 10100 54032
rect 9964 53740 10004 53780
rect 9868 52984 9908 53024
rect 9292 51052 9332 51092
rect 9100 50968 9140 51008
rect 9196 50716 9236 50756
rect 9292 49288 9332 49328
rect 9196 48112 9236 48152
rect 9292 47776 9332 47816
rect 9292 47440 9332 47480
rect 9580 52312 9620 52352
rect 9868 51808 9908 51848
rect 9772 50800 9812 50840
rect 9484 50380 9524 50420
rect 9484 50212 9524 50252
rect 9100 47104 9140 47144
rect 9292 46852 9332 46892
rect 9196 46600 9236 46640
rect 9196 45088 9236 45128
rect 9100 44416 9140 44456
rect 9100 44248 9140 44288
rect 9484 46180 9524 46220
rect 9676 48112 9716 48152
rect 9868 48028 9908 48068
rect 10156 53320 10196 53360
rect 10924 62896 10964 62936
rect 11308 63820 11348 63860
rect 10828 61048 10868 61088
rect 10636 60460 10676 60500
rect 10828 60712 10868 60752
rect 10636 59116 10676 59156
rect 11116 61804 11156 61844
rect 11020 61552 11060 61592
rect 11404 61804 11444 61844
rect 12364 73900 12404 73940
rect 13228 84820 13268 84860
rect 13324 84400 13364 84440
rect 14092 84484 14132 84524
rect 14476 84904 14516 84944
rect 14668 84568 14708 84608
rect 14860 84484 14900 84524
rect 15436 85576 15476 85616
rect 13708 84400 13748 84440
rect 13900 84400 13940 84440
rect 14284 84400 14324 84440
rect 15052 84400 15092 84440
rect 15244 84400 15284 84440
rect 14956 83728 14996 83768
rect 15724 85828 15764 85868
rect 13516 83476 13556 83516
rect 15148 83476 15188 83516
rect 13900 82804 13940 82844
rect 13228 80536 13268 80576
rect 13132 79276 13172 79316
rect 12940 78100 12980 78140
rect 13036 77176 13076 77216
rect 12844 76840 12884 76880
rect 12748 76588 12788 76628
rect 12748 76252 12788 76292
rect 12652 76084 12692 76124
rect 12748 74656 12788 74696
rect 12652 74488 12692 74528
rect 12556 74320 12596 74360
rect 12460 73396 12500 73436
rect 12748 74152 12788 74192
rect 12652 73816 12692 73856
rect 12364 71380 12404 71420
rect 12748 72136 12788 72176
rect 12268 69112 12308 69152
rect 12172 68104 12212 68144
rect 12076 66760 12116 66800
rect 12460 71296 12500 71336
rect 12652 70960 12692 71000
rect 11980 66088 12020 66128
rect 12268 65668 12308 65708
rect 11788 63904 11828 63944
rect 11692 61720 11732 61760
rect 11884 63400 11924 63440
rect 11500 61384 11540 61424
rect 11212 60796 11252 60836
rect 11308 60712 11348 60752
rect 11500 59956 11540 59996
rect 11404 59620 11444 59660
rect 10924 59200 10964 59240
rect 11020 58948 11060 58988
rect 10924 58444 10964 58484
rect 10924 57856 10964 57896
rect 11212 58444 11252 58484
rect 11788 58528 11828 58568
rect 10636 56680 10676 56720
rect 10828 56680 10868 56720
rect 11020 56596 11060 56636
rect 10924 56260 10964 56300
rect 11404 57352 11444 57392
rect 11020 55924 11060 55964
rect 11212 55588 11252 55628
rect 10636 55168 10676 55208
rect 10828 55168 10868 55208
rect 10540 54748 10580 54788
rect 10540 54160 10580 54200
rect 10252 53236 10292 53276
rect 10156 52900 10196 52940
rect 10540 53068 10580 53108
rect 10348 52564 10388 52604
rect 10732 53824 10772 53864
rect 10924 54160 10964 54200
rect 10828 53320 10868 53360
rect 11212 53908 11252 53948
rect 11884 57940 11924 57980
rect 11884 57688 11924 57728
rect 12364 63939 12404 63944
rect 12364 63904 12404 63939
rect 12268 61636 12308 61676
rect 12172 61300 12212 61340
rect 12556 69280 12596 69320
rect 12748 69112 12788 69152
rect 12748 68440 12788 68480
rect 12748 67768 12788 67808
rect 12556 65668 12596 65708
rect 12652 65248 12692 65288
rect 12652 63988 12692 64028
rect 12748 63232 12788 63272
rect 12748 63064 12788 63104
rect 12460 61468 12500 61508
rect 12460 61132 12500 61172
rect 12172 60628 12212 60668
rect 12076 60040 12116 60080
rect 12460 60460 12500 60500
rect 12652 60376 12692 60416
rect 12172 57940 12212 57980
rect 11980 57016 12020 57056
rect 12076 55588 12116 55628
rect 11404 54832 11444 54872
rect 10828 53068 10868 53108
rect 10732 52900 10772 52940
rect 10156 52396 10196 52436
rect 10732 52480 10772 52520
rect 10252 52312 10292 52352
rect 10444 52228 10484 52268
rect 10444 51892 10484 51932
rect 10156 49792 10196 49832
rect 10156 49540 10196 49580
rect 10060 48784 10100 48824
rect 10252 48784 10292 48824
rect 10252 48196 10292 48236
rect 10252 47944 10292 47984
rect 10348 47104 10388 47144
rect 10252 46852 10292 46892
rect 9580 46012 9620 46052
rect 9676 45844 9716 45884
rect 9580 45760 9620 45800
rect 9388 45508 9428 45548
rect 9292 44920 9332 44960
rect 9004 43744 9044 43784
rect 9100 42652 9140 42692
rect 9100 40468 9140 40508
rect 9004 40384 9044 40424
rect 10252 46348 10292 46388
rect 10060 46180 10100 46220
rect 9868 46012 9908 46052
rect 9868 45340 9908 45380
rect 9964 45172 10004 45212
rect 9868 45088 9908 45128
rect 9772 45004 9812 45044
rect 9676 44920 9716 44960
rect 9580 42820 9620 42860
rect 9772 42820 9812 42860
rect 9772 41896 9812 41936
rect 9676 41812 9716 41852
rect 9388 40300 9428 40340
rect 9964 43492 10004 43532
rect 10924 52648 10964 52688
rect 10924 52480 10964 52520
rect 10636 52312 10676 52352
rect 10924 52312 10964 52352
rect 10636 52060 10676 52100
rect 10636 49288 10676 49328
rect 11116 53320 11156 53360
rect 11116 53068 11156 53108
rect 11116 52816 11156 52856
rect 11308 53236 11348 53276
rect 11788 54916 11828 54956
rect 11500 53992 11540 54032
rect 11596 53824 11636 53864
rect 11500 53656 11540 53696
rect 11116 52312 11156 52352
rect 11020 52228 11060 52268
rect 11692 53320 11732 53360
rect 12076 53992 12116 54032
rect 11980 52900 12020 52940
rect 11788 52648 11828 52688
rect 11788 52480 11828 52520
rect 11884 52060 11924 52100
rect 10732 47776 10772 47816
rect 10924 47776 10964 47816
rect 10924 47356 10964 47396
rect 10828 47272 10868 47312
rect 10924 47188 10964 47228
rect 10828 46852 10868 46892
rect 11500 51808 11540 51848
rect 11212 50296 11252 50336
rect 11116 50212 11156 50252
rect 11404 50464 11444 50504
rect 11788 49624 11828 49664
rect 11308 49372 11348 49412
rect 11116 49120 11156 49160
rect 11596 49120 11636 49160
rect 11500 48868 11540 48908
rect 11500 48280 11540 48320
rect 11692 48532 11732 48572
rect 11404 47860 11444 47900
rect 11884 48448 11924 48488
rect 10252 44752 10292 44792
rect 10348 44500 10388 44540
rect 10252 44248 10292 44288
rect 10060 42652 10100 42692
rect 9964 41896 10004 41936
rect 10252 42232 10292 42272
rect 10156 41896 10196 41936
rect 10060 41812 10100 41852
rect 10060 41308 10100 41348
rect 9100 39544 9140 39584
rect 8908 38200 8948 38240
rect 8812 37612 8852 37652
rect 8332 36520 8372 36560
rect 8812 36520 8852 36560
rect 8812 36016 8852 36056
rect 8620 35932 8660 35972
rect 8236 35260 8276 35300
rect 8620 35260 8660 35300
rect 7852 35176 7892 35216
rect 8236 35008 8276 35048
rect 7852 34924 7892 34964
rect 7756 34336 7796 34376
rect 7660 34252 7700 34292
rect 7180 33328 7220 33368
rect 7180 32740 7220 32780
rect 7084 32320 7124 32360
rect 6988 32068 7028 32108
rect 7756 34084 7796 34124
rect 7660 33832 7700 33872
rect 7564 33748 7604 33788
rect 7468 32740 7508 32780
rect 6988 31564 7028 31604
rect 7276 31480 7316 31520
rect 6892 31312 6932 31352
rect 7084 31144 7124 31184
rect 6412 30388 6452 30428
rect 6412 30052 6452 30092
rect 6700 30304 6740 30344
rect 6220 29632 6260 29672
rect 5932 29380 5972 29420
rect 5740 28204 5780 28244
rect 4588 26776 4628 26816
rect 4492 25264 4532 25304
rect 4396 25180 4436 25220
rect 4396 24340 4436 24380
rect 3628 23164 3668 23204
rect 4204 23164 4244 23204
rect 3820 23080 3860 23120
rect 4108 22912 4148 22952
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 4012 22492 4052 22532
rect 3916 22408 3956 22448
rect 3340 22324 3380 22364
rect 3628 22240 3668 22280
rect 3820 22240 3860 22280
rect 3532 22156 3572 22196
rect 3532 21652 3572 21692
rect 3724 21652 3764 21692
rect 3340 21568 3380 21608
rect 3628 21568 3668 21608
rect 4108 22240 4148 22280
rect 4300 22576 4340 22616
rect 4588 23920 4628 23960
rect 4588 23584 4628 23624
rect 4492 23500 4532 23540
rect 4588 23416 4628 23456
rect 4492 23164 4532 23204
rect 4396 21988 4436 22028
rect 4204 21736 4244 21776
rect 4588 22324 4628 22364
rect 5164 27448 5204 27488
rect 5356 27448 5396 27488
rect 4876 26776 4916 26816
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 5068 26272 5108 26312
rect 5740 27784 5780 27824
rect 5740 27196 5780 27236
rect 5644 27028 5684 27068
rect 4780 25516 4820 25556
rect 5548 25348 5588 25388
rect 5068 25180 5108 25220
rect 5356 25180 5396 25220
rect 4972 25096 5012 25136
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 5452 24928 5492 24968
rect 5356 24592 5396 24632
rect 4876 24508 4916 24548
rect 4972 24256 5012 24296
rect 5068 23584 5108 23624
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 4780 22828 4820 22868
rect 4780 22660 4820 22700
rect 5932 27280 5972 27320
rect 6028 26776 6068 26816
rect 5836 26608 5876 26648
rect 5836 25348 5876 25388
rect 6028 25684 6068 25724
rect 5740 24844 5780 24884
rect 5644 23920 5684 23960
rect 6124 24676 6164 24716
rect 5836 24340 5876 24380
rect 6124 24340 6164 24380
rect 5548 23080 5588 23120
rect 6028 23752 6068 23792
rect 5932 23164 5972 23204
rect 5452 22660 5492 22700
rect 5644 22660 5684 22700
rect 5356 22492 5396 22532
rect 5452 22408 5492 22448
rect 5260 22072 5300 22112
rect 4396 21484 4436 21524
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 4108 20392 4148 20432
rect 4684 21736 4724 21776
rect 5356 21652 5396 21692
rect 4300 20224 4340 20264
rect 3532 19804 3572 19844
rect 4012 19804 4052 19844
rect 3340 18544 3380 18584
rect 3436 18040 3476 18080
rect 3340 17956 3380 17996
rect 2860 17872 2900 17912
rect 2764 17788 2804 17828
rect 2476 17032 2516 17072
rect 2284 16192 2324 16232
rect 2188 14176 2228 14216
rect 2092 11236 2132 11276
rect 1996 10900 2036 10940
rect 1804 9724 1844 9764
rect 1612 9472 1652 9512
rect 364 8632 404 8672
rect 1900 9388 1940 9428
rect 2476 15100 2516 15140
rect 2668 17200 2708 17240
rect 2668 17032 2708 17072
rect 2956 17788 2996 17828
rect 3052 17536 3092 17576
rect 2956 17368 2996 17408
rect 2860 16864 2900 16904
rect 2764 16192 2804 16232
rect 2860 15772 2900 15812
rect 2860 15100 2900 15140
rect 3436 17536 3476 17576
rect 3239 17116 3279 17156
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 4300 19888 4340 19928
rect 4684 20644 4724 20684
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 5452 21568 5492 21608
rect 5548 21400 5588 21440
rect 5452 20560 5492 20600
rect 5452 20308 5492 20348
rect 4684 20140 4724 20180
rect 4492 19888 4532 19928
rect 5068 19888 5108 19928
rect 4300 19300 4340 19340
rect 4780 19216 4820 19256
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 4108 18628 4148 18668
rect 5068 18628 5108 18668
rect 4204 18544 4244 18584
rect 4204 18376 4244 18416
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 3820 17620 3860 17660
rect 3916 17200 3956 17240
rect 3244 16864 3284 16904
rect 3436 16864 3476 16904
rect 3340 16696 3380 16736
rect 3724 17032 3764 17072
rect 4108 17284 4148 17324
rect 4972 18544 5012 18584
rect 4396 17956 4436 17996
rect 4300 17284 4340 17324
rect 4204 17200 4244 17240
rect 5164 17788 5204 17828
rect 4876 17704 4916 17744
rect 5068 17704 5108 17744
rect 4684 17536 4724 17576
rect 5356 18460 5396 18500
rect 5452 18124 5492 18164
rect 5452 17788 5492 17828
rect 5356 17704 5396 17744
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 4588 17116 4628 17156
rect 4012 16864 4052 16904
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 4492 17032 4532 17072
rect 4204 16780 4244 16820
rect 4300 16612 4340 16652
rect 3628 16444 3668 16484
rect 3532 16360 3572 16400
rect 3532 15940 3572 15980
rect 3916 16360 3956 16400
rect 3724 16108 3764 16148
rect 4204 16360 4244 16400
rect 4108 16192 4148 16232
rect 4012 15940 4052 15980
rect 4012 15520 4052 15560
rect 3340 15100 3380 15140
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 4012 14848 4052 14888
rect 2476 11068 2516 11108
rect 2476 10144 2516 10184
rect 2380 8212 2420 8252
rect 2956 14344 2996 14384
rect 3244 14596 3284 14636
rect 3148 14176 3188 14216
rect 2956 13252 2996 13292
rect 2860 12580 2900 12620
rect 2668 12412 2708 12452
rect 3148 13000 3188 13040
rect 2860 12160 2900 12200
rect 3148 12244 3188 12284
rect 3148 11908 3188 11948
rect 3052 11824 3092 11864
rect 2860 11236 2900 11276
rect 2956 10984 2996 11024
rect 3532 14680 3572 14720
rect 3724 14680 3764 14720
rect 3436 14596 3476 14636
rect 4012 14512 4052 14552
rect 3532 14008 3572 14048
rect 3820 14260 3860 14300
rect 3820 14008 3860 14048
rect 5356 16612 5396 16652
rect 4588 16360 4628 16400
rect 4876 16360 4916 16400
rect 4588 16192 4628 16232
rect 6028 22828 6068 22868
rect 5932 21988 5972 22028
rect 5836 21736 5876 21776
rect 5740 19888 5780 19928
rect 5644 19804 5684 19844
rect 5644 18628 5684 18668
rect 5644 18376 5684 18416
rect 5548 17620 5588 17660
rect 5452 16192 5492 16232
rect 4492 15940 4532 15980
rect 4396 15268 4436 15308
rect 4300 14848 4340 14888
rect 4396 14512 4436 14552
rect 4588 14428 4628 14468
rect 4108 14176 4148 14216
rect 4588 14176 4628 14216
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 5548 15604 5588 15644
rect 4972 15352 5012 15392
rect 5644 15436 5684 15476
rect 6316 29128 6356 29168
rect 6604 29800 6644 29840
rect 6988 30220 7028 30260
rect 7276 30640 7316 30680
rect 7372 30556 7412 30596
rect 7180 30136 7220 30176
rect 7084 30052 7124 30092
rect 6700 29128 6740 29168
rect 6988 29128 7028 29168
rect 7276 29380 7316 29420
rect 7180 29128 7220 29168
rect 7468 29128 7508 29168
rect 6892 28456 6932 28496
rect 6508 27700 6548 27740
rect 6316 27028 6356 27068
rect 6604 27364 6644 27404
rect 6508 27280 6548 27320
rect 6412 25684 6452 25724
rect 6604 27196 6644 27236
rect 6316 25012 6356 25052
rect 6220 23752 6260 23792
rect 6220 21568 6260 21608
rect 6124 21484 6164 21524
rect 6796 27616 6836 27656
rect 6988 28288 7028 28328
rect 7276 28288 7316 28328
rect 6892 26440 6932 26480
rect 7180 28204 7220 28244
rect 7084 25936 7124 25976
rect 6988 25432 7028 25472
rect 7084 25264 7124 25304
rect 6700 24592 6740 24632
rect 6892 23920 6932 23960
rect 6604 23248 6644 23288
rect 6796 23248 6836 23288
rect 6508 23164 6548 23204
rect 6892 22912 6932 22952
rect 6508 22660 6548 22700
rect 6604 22240 6644 22280
rect 6508 21568 6548 21608
rect 6412 20644 6452 20684
rect 6124 20224 6164 20264
rect 6124 19636 6164 19676
rect 6028 19300 6068 19340
rect 6028 19048 6068 19088
rect 6220 19468 6260 19508
rect 6412 19720 6452 19760
rect 6892 22156 6932 22196
rect 6796 22072 6836 22112
rect 6700 21568 6740 21608
rect 6892 21736 6932 21776
rect 6892 21484 6932 21524
rect 7084 23080 7124 23120
rect 6988 21400 7028 21440
rect 7276 27616 7316 27656
rect 7660 32740 7700 32780
rect 7756 32152 7796 32192
rect 8044 34084 8084 34124
rect 7948 32992 7988 33032
rect 8044 32908 8084 32948
rect 7948 32740 7988 32780
rect 7660 31144 7700 31184
rect 7852 30808 7892 30848
rect 7852 30640 7892 30680
rect 8044 32320 8084 32360
rect 8044 31312 8084 31352
rect 7660 29128 7700 29168
rect 8140 31228 8180 31268
rect 8140 30976 8180 31016
rect 8524 34924 8564 34964
rect 8524 34588 8564 34628
rect 8332 32992 8372 33032
rect 8044 30220 8084 30260
rect 7852 29800 7892 29840
rect 7564 28456 7604 28496
rect 8524 32740 8564 32780
rect 8428 32404 8468 32444
rect 8524 31312 8564 31352
rect 9964 39712 10004 39752
rect 9868 39628 9908 39668
rect 9676 38536 9716 38576
rect 9676 38200 9716 38240
rect 9196 37360 9236 37400
rect 9196 36016 9236 36056
rect 9100 35176 9140 35216
rect 9196 35092 9236 35132
rect 8812 33664 8852 33704
rect 9196 34084 9236 34124
rect 9004 33664 9044 33704
rect 8812 32068 8852 32108
rect 8812 31480 8852 31520
rect 8716 31144 8756 31184
rect 8620 30976 8660 31016
rect 8332 30472 8372 30512
rect 8236 29716 8276 29756
rect 8236 29296 8276 29336
rect 8524 30136 8564 30176
rect 8620 30052 8660 30092
rect 8236 29128 8276 29168
rect 8044 27616 8084 27656
rect 7756 27196 7796 27236
rect 7948 27112 7988 27152
rect 7468 26860 7508 26900
rect 7372 26776 7412 26816
rect 7276 26608 7316 26648
rect 7852 26440 7892 26480
rect 7756 25264 7796 25304
rect 7564 25180 7604 25220
rect 7564 24760 7604 24800
rect 8428 27448 8468 27488
rect 8236 27196 8276 27236
rect 8524 26860 8564 26900
rect 8332 26776 8372 26816
rect 8332 26104 8372 26144
rect 8332 25768 8372 25808
rect 7372 24592 7412 24632
rect 7756 24592 7796 24632
rect 7948 24592 7988 24632
rect 7948 24172 7988 24212
rect 7276 23920 7316 23960
rect 7468 23920 7508 23960
rect 7852 23920 7892 23960
rect 7276 23668 7316 23708
rect 7180 22996 7220 23036
rect 7948 23332 7988 23372
rect 7564 23164 7604 23204
rect 7468 22912 7508 22952
rect 7468 22660 7508 22700
rect 7276 22408 7316 22448
rect 7372 22324 7412 22364
rect 7180 22240 7220 22280
rect 7276 21988 7316 22028
rect 7180 21820 7220 21860
rect 7948 23080 7988 23120
rect 8524 26272 8564 26312
rect 8428 25180 8468 25220
rect 8524 24760 8564 24800
rect 7660 21904 7700 21944
rect 7372 21820 7412 21860
rect 7564 21820 7604 21860
rect 7468 21568 7508 21608
rect 7468 21400 7508 21440
rect 7372 20140 7412 20180
rect 6700 19300 6740 19340
rect 6796 19132 6836 19172
rect 7276 19048 7316 19088
rect 5836 18628 5876 18668
rect 6220 18712 6260 18752
rect 5932 18460 5972 18500
rect 5836 18124 5876 18164
rect 5836 17872 5876 17912
rect 6028 17536 6068 17576
rect 6028 15856 6068 15896
rect 5836 15436 5876 15476
rect 5932 15016 5972 15056
rect 5260 14680 5300 14720
rect 5260 14512 5300 14552
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 5164 14176 5204 14216
rect 4012 13924 4052 13964
rect 4300 13924 4340 13964
rect 4108 13840 4148 13880
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 3340 12664 3380 12704
rect 3340 12496 3380 12536
rect 3532 12496 3572 12536
rect 4012 13252 4052 13292
rect 3916 13168 3956 13208
rect 4108 13000 4148 13040
rect 3916 12580 3956 12620
rect 3820 12496 3860 12536
rect 4012 12496 4052 12536
rect 3436 12328 3476 12368
rect 3340 12244 3380 12284
rect 3244 11656 3284 11696
rect 3436 11824 3476 11864
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 3916 11908 3956 11948
rect 3724 11824 3764 11864
rect 3340 11488 3380 11528
rect 4108 11656 4148 11696
rect 4300 12664 4340 12704
rect 4396 12412 4436 12452
rect 4300 12076 4340 12116
rect 4684 13672 4724 13712
rect 4588 13168 4628 13208
rect 4684 12580 4724 12620
rect 4588 12328 4628 12368
rect 5252 14092 5292 14132
rect 4972 13756 5012 13796
rect 5164 13588 5204 13628
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 4876 12580 4916 12620
rect 5260 12580 5300 12620
rect 4972 12412 5012 12452
rect 5260 12244 5300 12284
rect 4492 11740 4532 11780
rect 4780 11824 4820 11864
rect 4972 11824 5012 11864
rect 4684 11656 4724 11696
rect 4492 11488 4532 11528
rect 2764 10060 2804 10100
rect 2956 10060 2996 10100
rect 2860 9472 2900 9512
rect 3244 9472 3284 9512
rect 2860 9304 2900 9344
rect 2572 7792 2612 7832
rect 3436 11320 3476 11360
rect 3724 11236 3764 11276
rect 3532 11068 3572 11108
rect 3436 10144 3476 10184
rect 4204 11152 4244 11192
rect 4108 10984 4148 11024
rect 3724 10816 3764 10856
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 3820 10312 3860 10352
rect 3628 10060 3668 10100
rect 4300 10732 4340 10772
rect 3916 9976 3956 10016
rect 3436 9472 3476 9512
rect 3916 9556 3956 9596
rect 3628 9472 3668 9512
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 6028 14680 6068 14720
rect 6220 18124 6260 18164
rect 6412 18544 6452 18584
rect 6700 18712 6740 18752
rect 6796 18544 6836 18584
rect 6988 18544 7028 18584
rect 6412 18292 6452 18332
rect 6412 17956 6452 17996
rect 6316 17788 6356 17828
rect 5836 14344 5876 14384
rect 5740 14008 5780 14048
rect 5644 13924 5684 13964
rect 5836 13840 5876 13880
rect 5644 13168 5684 13208
rect 5644 12832 5684 12872
rect 5644 12664 5684 12704
rect 5548 12496 5588 12536
rect 5740 12496 5780 12536
rect 5452 12328 5492 12368
rect 5452 11152 5492 11192
rect 5164 10984 5204 11024
rect 5356 10984 5396 11024
rect 4780 10732 4820 10772
rect 3436 9220 3476 9260
rect 3052 8548 3092 8588
rect 2956 8380 2996 8420
rect 2956 7960 2996 8000
rect 3340 8632 3380 8672
rect 3148 8380 3188 8420
rect 3244 8296 3284 8336
rect 3148 3676 3188 3716
rect 2956 1240 2996 1280
rect 2572 904 2612 944
rect 2764 568 2804 608
rect 3635 9220 3675 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3628 8884 3668 8924
rect 3916 8884 3956 8924
rect 3724 8800 3764 8840
rect 3827 8800 3867 8840
rect 3628 8296 3668 8336
rect 3532 8128 3572 8168
rect 4012 8632 4052 8672
rect 3916 8548 3956 8588
rect 3916 8128 3956 8168
rect 3532 7960 3572 8000
rect 4396 9472 4436 9512
rect 4300 9304 4340 9344
rect 4492 9220 4532 9260
rect 4492 8968 4532 9008
rect 4204 8464 4244 8504
rect 4108 8296 4148 8336
rect 4108 8128 4148 8168
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 4204 7540 4244 7580
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 3340 3172 3380 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4396 8632 4436 8672
rect 4492 8380 4532 8420
rect 5740 10984 5780 11024
rect 6028 14344 6068 14384
rect 6124 14260 6164 14300
rect 6412 14260 6452 14300
rect 6124 14008 6164 14048
rect 6316 13924 6356 13964
rect 6412 13756 6452 13796
rect 6028 13588 6068 13628
rect 6124 13504 6164 13544
rect 6124 12832 6164 12872
rect 5932 12664 5972 12704
rect 5932 12328 5972 12368
rect 6604 18124 6644 18164
rect 6604 17536 6644 17576
rect 6892 17704 6932 17744
rect 7084 17704 7124 17744
rect 7180 17536 7220 17576
rect 7564 21316 7604 21356
rect 7564 19048 7604 19088
rect 7564 18712 7604 18752
rect 7660 18376 7700 18416
rect 7852 22240 7892 22280
rect 8140 22072 8180 22112
rect 7948 21736 7988 21776
rect 8044 21568 8084 21608
rect 8716 29800 8756 29840
rect 8716 27364 8756 27404
rect 9004 31396 9044 31436
rect 9196 31396 9236 31436
rect 9196 31144 9236 31184
rect 8908 30220 8948 30260
rect 8908 29968 8948 30008
rect 9100 29800 9140 29840
rect 9388 37360 9428 37400
rect 9388 36520 9428 36560
rect 9772 36688 9812 36728
rect 10156 39712 10196 39752
rect 10156 39040 10196 39080
rect 10252 38956 10292 38996
rect 10252 38536 10292 38576
rect 10252 38200 10292 38240
rect 9868 36520 9908 36560
rect 9676 35848 9716 35888
rect 9772 35764 9812 35804
rect 9772 35260 9812 35300
rect 9388 34420 9428 34460
rect 9868 35176 9908 35216
rect 9676 35008 9716 35048
rect 9868 35008 9908 35048
rect 9676 34756 9716 34796
rect 9580 34336 9620 34376
rect 9388 34252 9428 34292
rect 9484 34084 9524 34124
rect 9772 34504 9812 34544
rect 9772 34000 9812 34040
rect 10444 38704 10484 38744
rect 10924 46348 10964 46388
rect 10828 45760 10868 45800
rect 11020 45592 11060 45632
rect 10924 45424 10964 45464
rect 10732 45004 10772 45044
rect 10924 43660 10964 43700
rect 10732 42736 10772 42776
rect 10732 41896 10772 41936
rect 11212 46432 11252 46472
rect 11212 45256 11252 45296
rect 11404 45172 11444 45212
rect 11308 43408 11348 43448
rect 11116 40972 11156 41012
rect 11212 40636 11252 40676
rect 11596 46516 11636 46556
rect 11596 45676 11636 45716
rect 11980 46600 12020 46640
rect 12364 57016 12404 57056
rect 12460 56344 12500 56384
rect 12460 55588 12500 55628
rect 12460 53656 12500 53696
rect 13420 80200 13460 80240
rect 13420 79360 13460 79400
rect 13804 81292 13844 81332
rect 13708 79528 13748 79568
rect 13324 76924 13364 76964
rect 13132 76672 13172 76712
rect 13708 76840 13748 76880
rect 13516 76672 13556 76712
rect 13420 76252 13460 76292
rect 13324 76168 13364 76208
rect 12940 75496 12980 75536
rect 13036 75160 13076 75200
rect 13132 74404 13172 74444
rect 12940 73900 12980 73940
rect 13228 73816 13268 73856
rect 13132 73564 13172 73604
rect 13036 73396 13076 73436
rect 13228 72220 13268 72260
rect 13132 72136 13172 72176
rect 13036 71464 13076 71504
rect 13228 71968 13268 72008
rect 12940 67600 12980 67640
rect 13420 74068 13460 74108
rect 13420 73900 13460 73940
rect 13420 71968 13460 72008
rect 13612 76084 13652 76124
rect 14284 82216 14324 82256
rect 15724 83056 15764 83096
rect 15340 81880 15380 81920
rect 14284 79780 14324 79820
rect 14092 79696 14132 79736
rect 14188 79276 14228 79316
rect 14092 78184 14132 78224
rect 14572 79360 14612 79400
rect 14380 78100 14420 78140
rect 14572 78100 14612 78140
rect 14764 78100 14804 78140
rect 14092 76672 14132 76712
rect 14092 75580 14132 75620
rect 13900 75160 13940 75200
rect 13804 74152 13844 74192
rect 13708 73396 13748 73436
rect 13612 72724 13652 72764
rect 13804 73060 13844 73100
rect 14284 75244 14324 75284
rect 14572 75244 14612 75284
rect 14092 74908 14132 74948
rect 13900 72136 13940 72176
rect 13708 72052 13748 72092
rect 13996 71968 14036 72008
rect 13900 71800 13940 71840
rect 13708 71548 13748 71588
rect 13708 70876 13748 70916
rect 13516 69952 13556 69992
rect 13132 69112 13172 69152
rect 13708 69112 13748 69152
rect 13036 66928 13076 66968
rect 13036 66424 13076 66464
rect 12940 65500 12980 65540
rect 12844 60292 12884 60332
rect 13036 61216 13076 61256
rect 13420 67600 13460 67640
rect 14380 74320 14420 74360
rect 15916 83476 15956 83516
rect 15532 79780 15572 79820
rect 15916 79780 15956 79820
rect 15340 79276 15380 79316
rect 15244 78856 15284 78896
rect 15052 78016 15092 78056
rect 14764 76168 14804 76208
rect 14188 73984 14228 74024
rect 14284 73816 14324 73856
rect 14284 73564 14324 73604
rect 14188 71800 14228 71840
rect 14092 71296 14132 71336
rect 13900 69952 13940 69992
rect 13324 63904 13364 63944
rect 13420 63568 13460 63608
rect 13324 61720 13364 61760
rect 13324 60460 13364 60500
rect 12940 60124 12980 60164
rect 12748 60040 12788 60080
rect 12844 59956 12884 59996
rect 13324 60040 13364 60080
rect 12748 58528 12788 58568
rect 12748 58024 12788 58064
rect 12940 59788 12980 59828
rect 13420 58780 13460 58820
rect 13420 58612 13460 58652
rect 13132 57856 13172 57896
rect 13612 66592 13652 66632
rect 13612 66088 13652 66128
rect 14188 70876 14228 70916
rect 14092 70540 14132 70580
rect 13996 69364 14036 69404
rect 14668 73648 14708 73688
rect 15244 78100 15284 78140
rect 15148 76588 15188 76628
rect 15436 77344 15476 77384
rect 15340 76336 15380 76376
rect 15052 76168 15092 76208
rect 15244 76000 15284 76040
rect 15724 77260 15764 77300
rect 15628 76840 15668 76880
rect 14956 74572 14996 74612
rect 14860 73900 14900 73940
rect 15340 75496 15380 75536
rect 15052 73984 15092 74024
rect 14764 71548 14804 71588
rect 14476 71464 14516 71504
rect 15724 75916 15764 75956
rect 15628 75496 15668 75536
rect 15628 75244 15668 75284
rect 15628 74656 15668 74696
rect 15340 74488 15380 74528
rect 15244 73900 15284 73940
rect 15340 73648 15380 73688
rect 14956 72136 14996 72176
rect 14380 69952 14420 69992
rect 14188 68944 14228 68984
rect 14092 68272 14132 68312
rect 14092 67096 14132 67136
rect 14284 67264 14324 67304
rect 14860 71044 14900 71084
rect 14860 70876 14900 70916
rect 14860 70540 14900 70580
rect 14764 70456 14804 70496
rect 14668 69028 14708 69068
rect 15148 72892 15188 72932
rect 15148 72304 15188 72344
rect 15244 72220 15284 72260
rect 15148 72136 15188 72176
rect 15052 71800 15092 71840
rect 15052 71548 15092 71588
rect 14956 69868 14996 69908
rect 14956 69700 14996 69740
rect 14764 68440 14804 68480
rect 14572 68020 14612 68060
rect 15148 71296 15188 71336
rect 15148 70456 15188 70496
rect 15148 69700 15188 69740
rect 15340 72136 15380 72176
rect 15820 74320 15860 74360
rect 15820 74152 15860 74192
rect 15628 72976 15668 73016
rect 15532 71968 15572 72008
rect 15340 71800 15380 71840
rect 15532 71499 15572 71504
rect 15532 71464 15572 71499
rect 15724 71632 15764 71672
rect 15340 70456 15380 70496
rect 15436 69952 15476 69992
rect 15148 68944 15188 68984
rect 15052 67684 15092 67724
rect 14572 67600 14612 67640
rect 14764 67600 14804 67640
rect 14476 67096 14516 67136
rect 13996 66340 14036 66380
rect 13900 65500 13940 65540
rect 13804 65416 13844 65456
rect 13996 64576 14036 64616
rect 13612 64156 13652 64196
rect 13996 63904 14036 63944
rect 13804 63064 13844 63104
rect 13708 62980 13748 63020
rect 13612 62812 13652 62852
rect 13900 61216 13940 61256
rect 13804 60292 13844 60332
rect 13708 59872 13748 59912
rect 13804 59704 13844 59744
rect 13708 59620 13748 59660
rect 13804 59200 13844 59240
rect 13708 58696 13748 58736
rect 13516 57268 13556 57308
rect 13228 57100 13268 57140
rect 13420 56932 13460 56972
rect 13804 58444 13844 58484
rect 14188 66340 14228 66380
rect 14572 66844 14612 66884
rect 14284 64324 14324 64364
rect 14764 66928 14804 66968
rect 15340 68440 15380 68480
rect 15340 68272 15380 68312
rect 15628 70456 15668 70496
rect 15724 69952 15764 69992
rect 15532 68188 15572 68228
rect 15244 67096 15284 67136
rect 14956 66844 14996 66884
rect 15148 66844 15188 66884
rect 14380 63820 14420 63860
rect 14476 63232 14516 63272
rect 14092 61720 14132 61760
rect 14092 61552 14132 61592
rect 13996 59620 14036 59660
rect 13708 56932 13748 56972
rect 13612 56680 13652 56720
rect 13900 56680 13940 56720
rect 13228 56344 13268 56384
rect 14668 63904 14708 63944
rect 14572 61720 14612 61760
rect 14572 61384 14612 61424
rect 14572 61216 14612 61256
rect 14284 60460 14324 60500
rect 14284 59704 14324 59744
rect 13708 56092 13748 56132
rect 12652 53992 12692 54032
rect 12748 53488 12788 53528
rect 12460 53236 12500 53276
rect 12364 53068 12404 53108
rect 12364 52900 12404 52940
rect 12652 53320 12692 53360
rect 12556 52648 12596 52688
rect 12748 52564 12788 52604
rect 12268 52312 12308 52352
rect 12460 52060 12500 52100
rect 12268 51136 12308 51176
rect 12172 50296 12212 50336
rect 12172 48280 12212 48320
rect 12172 47272 12212 47312
rect 12364 50296 12404 50336
rect 12556 51808 12596 51848
rect 12748 51808 12788 51848
rect 13228 54832 13268 54872
rect 12940 54160 12980 54200
rect 12940 53152 12980 53192
rect 12940 52900 12980 52940
rect 13516 53824 13556 53864
rect 13228 53488 13268 53528
rect 13420 53488 13460 53528
rect 13132 53320 13172 53360
rect 13228 53236 13268 53276
rect 13132 52984 13172 53024
rect 13036 52816 13076 52856
rect 13036 52396 13076 52436
rect 12940 52144 12980 52184
rect 13036 51976 13076 52016
rect 12460 48280 12500 48320
rect 12652 50380 12692 50420
rect 13036 51556 13076 51596
rect 13228 52900 13268 52940
rect 13324 52312 13364 52352
rect 13612 53404 13652 53444
rect 13804 53992 13844 54032
rect 13713 52564 13753 52604
rect 13612 52480 13652 52520
rect 13516 52144 13556 52184
rect 13516 51976 13556 52016
rect 13804 51472 13844 51512
rect 13420 51052 13460 51092
rect 13228 50548 13268 50588
rect 13036 50212 13076 50252
rect 12940 49624 12980 49664
rect 12844 49540 12884 49580
rect 12940 49461 12980 49496
rect 12940 49456 12980 49461
rect 12364 48028 12404 48068
rect 12460 47944 12500 47984
rect 12556 46852 12596 46892
rect 11692 45592 11732 45632
rect 11788 44248 11828 44288
rect 11596 43492 11636 43532
rect 11500 41644 11540 41684
rect 11692 43156 11732 43196
rect 11788 41560 11828 41600
rect 11404 39880 11444 39920
rect 10828 38452 10868 38492
rect 10732 38368 10772 38408
rect 10636 38116 10676 38156
rect 10732 37948 10772 37988
rect 10348 36688 10388 36728
rect 10060 36520 10100 36560
rect 10060 35848 10100 35888
rect 10348 35680 10388 35720
rect 10156 35512 10196 35552
rect 9964 34756 10004 34796
rect 9964 34420 10004 34460
rect 10252 35176 10292 35216
rect 10732 36856 10772 36896
rect 10540 35932 10580 35972
rect 10444 34924 10484 34964
rect 10348 34840 10388 34880
rect 10252 34420 10292 34460
rect 10156 34084 10196 34124
rect 10060 34000 10100 34040
rect 8908 28540 8948 28580
rect 8716 25348 8756 25388
rect 8620 24340 8660 24380
rect 8620 24172 8660 24212
rect 9100 26440 9140 26480
rect 8524 23080 8564 23120
rect 8524 22912 8564 22952
rect 8332 21904 8372 21944
rect 7852 21148 7892 21188
rect 8332 20896 8372 20936
rect 8524 20896 8564 20936
rect 8716 23080 8756 23120
rect 9004 23080 9044 23120
rect 9484 30220 9524 30260
rect 9676 32068 9716 32108
rect 9388 28792 9428 28832
rect 9292 26272 9332 26312
rect 9196 24004 9236 24044
rect 9292 23920 9332 23960
rect 9196 23836 9236 23876
rect 9580 23920 9620 23960
rect 9868 32320 9908 32360
rect 9868 28456 9908 28496
rect 10156 32824 10196 32864
rect 10060 32320 10100 32360
rect 10348 33916 10388 33956
rect 10924 37612 10964 37652
rect 11020 36856 11060 36896
rect 11020 36688 11060 36728
rect 10924 36520 10964 36560
rect 10732 35428 10772 35468
rect 10732 34840 10772 34880
rect 10636 34420 10676 34460
rect 10732 34336 10772 34376
rect 10636 34168 10676 34208
rect 10540 33496 10580 33536
rect 10828 33664 10868 33704
rect 10732 33580 10772 33620
rect 10636 32908 10676 32948
rect 10732 32824 10772 32864
rect 10156 31312 10196 31352
rect 10924 32992 10964 33032
rect 10924 32824 10964 32864
rect 11212 38200 11252 38240
rect 11596 41308 11636 41348
rect 11212 37108 11252 37148
rect 11308 36436 11348 36476
rect 11308 36184 11348 36224
rect 11500 36772 11540 36812
rect 11500 36604 11540 36644
rect 11500 36436 11540 36476
rect 11404 35932 11444 35972
rect 11212 34756 11252 34796
rect 11500 35512 11540 35552
rect 11404 34504 11444 34544
rect 11212 34168 11252 34208
rect 11404 33832 11444 33872
rect 11212 32908 11252 32948
rect 11020 32740 11060 32780
rect 10348 29800 10388 29840
rect 10828 30640 10868 30680
rect 10540 29884 10580 29924
rect 10252 28456 10292 28496
rect 10252 28288 10292 28328
rect 10060 27364 10100 27404
rect 10060 27196 10100 27236
rect 9964 26104 10004 26144
rect 10444 28288 10484 28328
rect 9964 24424 10004 24464
rect 9772 24088 9812 24128
rect 9964 23920 10004 23960
rect 10156 23920 10196 23960
rect 9676 23836 9716 23876
rect 9676 23668 9716 23708
rect 9484 23584 9524 23624
rect 9580 23416 9620 23456
rect 9388 23332 9428 23372
rect 9292 23248 9332 23288
rect 9772 23080 9812 23120
rect 8908 22576 8948 22616
rect 9196 22492 9236 22532
rect 9388 22828 9428 22868
rect 8812 21820 8852 21860
rect 9868 22828 9908 22868
rect 9580 22576 9620 22616
rect 9772 22492 9812 22532
rect 9484 22240 9524 22280
rect 9868 22240 9908 22280
rect 10156 22576 10196 22616
rect 9676 21652 9716 21692
rect 8716 21148 8756 21188
rect 9196 21148 9236 21188
rect 8620 20560 8660 20600
rect 8620 20392 8660 20432
rect 7948 20224 7988 20264
rect 8044 20056 8084 20096
rect 8140 19888 8180 19928
rect 8044 19300 8084 19340
rect 7948 18628 7988 18668
rect 8524 20224 8564 20264
rect 8332 19972 8372 20012
rect 8668 19972 8708 20012
rect 8572 19888 8612 19928
rect 8812 19720 8852 19760
rect 8908 19636 8948 19676
rect 8332 19048 8372 19088
rect 7948 18376 7988 18416
rect 7852 18208 7892 18248
rect 7756 17872 7796 17912
rect 7564 17536 7604 17576
rect 7468 17368 7508 17408
rect 6892 16696 6932 16736
rect 7084 16696 7124 16736
rect 6988 16360 7028 16400
rect 6604 14932 6644 14972
rect 6988 15520 7028 15560
rect 6988 15184 7028 15224
rect 6796 14344 6836 14384
rect 6796 14092 6836 14132
rect 6700 14008 6740 14048
rect 6604 13840 6644 13880
rect 6700 13504 6740 13544
rect 6508 13168 6548 13208
rect 6412 12832 6452 12872
rect 6220 11908 6260 11948
rect 6412 11908 6452 11948
rect 6124 11488 6164 11528
rect 6220 11404 6260 11444
rect 6988 13840 7028 13880
rect 6892 13084 6932 13124
rect 7660 17032 7700 17072
rect 7660 16696 7700 16736
rect 7564 16528 7604 16568
rect 7276 16360 7316 16400
rect 7468 15436 7508 15476
rect 7372 15268 7412 15308
rect 7276 14680 7316 14720
rect 7180 14176 7220 14216
rect 7084 13084 7124 13124
rect 7180 12916 7220 12956
rect 7084 12832 7124 12872
rect 6604 11656 6644 11696
rect 6892 11656 6932 11696
rect 7372 13000 7412 13040
rect 7564 15016 7604 15056
rect 7852 16780 7892 16820
rect 7756 14260 7796 14300
rect 8140 17872 8180 17912
rect 8044 17536 8084 17576
rect 8140 17368 8180 17408
rect 7948 15352 7988 15392
rect 8140 16780 8180 16820
rect 8620 18628 8660 18668
rect 8428 18124 8468 18164
rect 8524 17872 8564 17912
rect 8428 17620 8468 17660
rect 8716 18544 8756 18584
rect 9100 20056 9140 20096
rect 9388 19888 9428 19928
rect 9292 19552 9332 19592
rect 9100 19132 9140 19172
rect 9004 17620 9044 17660
rect 9772 21568 9812 21608
rect 9772 21148 9812 21188
rect 9580 20728 9620 20768
rect 9580 20560 9620 20600
rect 9484 18880 9524 18920
rect 9196 18124 9236 18164
rect 9196 17956 9236 17996
rect 9484 17872 9524 17912
rect 9388 17704 9428 17744
rect 9292 17620 9332 17660
rect 8716 17368 8756 17408
rect 9004 17200 9044 17240
rect 8908 16360 8948 16400
rect 8332 16192 8372 16232
rect 8236 15772 8276 15812
rect 8044 15100 8084 15140
rect 7948 15016 7988 15056
rect 8140 14932 8180 14972
rect 7948 14680 7988 14720
rect 8044 14428 8084 14468
rect 8236 14176 8276 14216
rect 7948 14092 7988 14132
rect 7852 13924 7892 13964
rect 7660 13504 7700 13544
rect 7468 12832 7508 12872
rect 7372 12664 7412 12704
rect 6604 11404 6644 11444
rect 6604 11236 6644 11276
rect 5932 11152 5972 11192
rect 5356 10564 5396 10604
rect 4876 10144 4916 10184
rect 5260 10144 5300 10184
rect 5644 10312 5684 10352
rect 5452 10144 5492 10184
rect 5159 9976 5199 10016
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 4684 9724 4724 9764
rect 5836 10900 5876 10940
rect 6028 10060 6068 10100
rect 5932 9976 5972 10016
rect 4876 8968 4916 9008
rect 5164 9472 5204 9512
rect 4972 8884 5012 8924
rect 4780 8800 4820 8840
rect 5548 8800 5588 8840
rect 4684 8716 4724 8756
rect 4876 8632 4916 8672
rect 4780 8548 4820 8588
rect 4684 8380 4724 8420
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4972 7960 5012 8000
rect 4780 7540 4820 7580
rect 4684 7456 4724 7496
rect 4492 7372 4532 7412
rect 4108 1912 4148 1952
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 3532 820 3572 860
rect 3340 64 3380 104
rect 3916 316 3956 356
rect 4300 484 4340 524
rect 5836 9808 5876 9848
rect 6508 11152 6548 11192
rect 6316 10984 6356 11024
rect 6412 10648 6452 10688
rect 7468 12160 7508 12200
rect 7276 11908 7316 11948
rect 7180 11404 7220 11444
rect 7084 11236 7124 11276
rect 6604 10732 6644 10772
rect 6316 9976 6356 10016
rect 6412 9472 6452 9512
rect 6220 9304 6260 9344
rect 5836 8380 5876 8420
rect 5836 8212 5876 8252
rect 5740 7372 5780 7412
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 5740 2080 5780 2120
rect 5356 988 5396 1028
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 5644 736 5684 776
rect 5452 568 5492 608
rect 5068 232 5108 272
rect 4876 148 4916 188
rect 6124 8800 6164 8840
rect 6316 8716 6356 8756
rect 7180 10984 7220 11024
rect 6988 10312 7028 10352
rect 7084 9808 7124 9848
rect 6988 9724 7028 9764
rect 6988 9472 7028 9512
rect 6892 9304 6932 9344
rect 6988 9136 7028 9176
rect 6316 8380 6356 8420
rect 6028 8128 6068 8168
rect 6316 7624 6356 7664
rect 6604 7624 6644 7664
rect 7084 8716 7124 8756
rect 7276 10228 7316 10268
rect 8044 13504 8084 13544
rect 7852 13168 7892 13208
rect 8524 15520 8564 15560
rect 8428 14932 8468 14972
rect 8524 14428 8564 14468
rect 8428 13924 8468 13964
rect 7948 13000 7988 13040
rect 8140 12916 8180 12956
rect 7852 12832 7892 12872
rect 7564 12076 7604 12116
rect 7564 11656 7604 11696
rect 8140 12496 8180 12536
rect 7948 12076 7988 12116
rect 7756 11488 7796 11528
rect 7564 10144 7604 10184
rect 7468 9220 7508 9260
rect 7372 9052 7412 9092
rect 7276 8380 7316 8420
rect 7180 8296 7220 8336
rect 7180 8128 7220 8168
rect 6988 5776 7028 5816
rect 6412 3760 6452 3800
rect 6124 2164 6164 2204
rect 5932 1492 5972 1532
rect 6316 1408 6356 1448
rect 6028 1240 6068 1280
rect 6892 2836 6932 2876
rect 6508 2080 6548 2120
rect 6892 2080 6932 2120
rect 7852 11404 7892 11444
rect 7756 7708 7796 7748
rect 7468 7540 7508 7580
rect 7756 7456 7796 7496
rect 8332 12580 8372 12620
rect 8236 11824 8276 11864
rect 8332 11740 8372 11780
rect 8140 10648 8180 10688
rect 8044 9472 8084 9512
rect 8140 8800 8180 8840
rect 8908 15604 8948 15644
rect 8908 15268 8948 15308
rect 8716 15100 8756 15140
rect 8812 14848 8852 14888
rect 8716 14428 8756 14468
rect 8908 13504 8948 13544
rect 9100 16108 9140 16148
rect 8716 13252 8756 13292
rect 9196 14680 9236 14720
rect 9100 12664 9140 12704
rect 9004 12580 9044 12620
rect 8812 11824 8852 11864
rect 8908 11740 8948 11780
rect 8428 10900 8468 10940
rect 8620 11068 8660 11108
rect 8812 10900 8852 10940
rect 8716 9724 8756 9764
rect 8044 7876 8084 7916
rect 8428 7456 8468 7496
rect 7852 3760 7892 3800
rect 8428 6448 8468 6488
rect 9004 11572 9044 11612
rect 9196 11572 9236 11612
rect 9484 17032 9524 17072
rect 9484 16528 9524 16568
rect 9676 20056 9716 20096
rect 9676 19636 9716 19676
rect 9676 18964 9716 19004
rect 10348 27448 10388 27488
rect 10348 24004 10388 24044
rect 10348 23164 10388 23204
rect 10252 22492 10292 22532
rect 10348 21484 10388 21524
rect 10348 21064 10388 21104
rect 10252 19720 10292 19760
rect 10348 19636 10388 19676
rect 11116 31480 11156 31520
rect 11308 32740 11348 32780
rect 11212 30976 11252 31016
rect 11116 30640 11156 30680
rect 11020 29884 11060 29924
rect 10924 29464 10964 29504
rect 11692 38704 11732 38744
rect 12076 46432 12116 46472
rect 12652 46348 12692 46388
rect 12652 45928 12692 45968
rect 12460 45760 12500 45800
rect 11980 42652 12020 42692
rect 11980 42400 12020 42440
rect 11980 41560 12020 41600
rect 12364 41728 12404 41768
rect 12556 43996 12596 44036
rect 12556 43492 12596 43532
rect 13132 49456 13172 49496
rect 12940 48616 12980 48656
rect 13036 48112 13076 48152
rect 13420 49876 13460 49916
rect 13420 48700 13460 48740
rect 13324 48112 13364 48152
rect 12940 46348 12980 46388
rect 12844 46012 12884 46052
rect 12940 44584 12980 44624
rect 12844 43912 12884 43952
rect 12076 41308 12116 41348
rect 11884 40300 11924 40340
rect 12172 39712 12212 39752
rect 13228 46096 13268 46136
rect 13420 46348 13460 46388
rect 13324 46012 13364 46052
rect 13420 45424 13460 45464
rect 13324 44584 13364 44624
rect 13708 50968 13748 51008
rect 13996 56008 14036 56048
rect 13996 53992 14036 54032
rect 14188 57016 14228 57056
rect 14380 56764 14420 56804
rect 14284 56344 14324 56384
rect 14188 54916 14228 54956
rect 14188 53992 14228 54032
rect 13708 50800 13748 50840
rect 13900 50800 13940 50840
rect 13900 49624 13940 49664
rect 14476 55336 14516 55376
rect 14380 54412 14420 54452
rect 14188 52480 14228 52520
rect 14284 52144 14324 52184
rect 14188 51640 14228 51680
rect 14092 51136 14132 51176
rect 14092 50968 14132 51008
rect 14092 49876 14132 49916
rect 13612 47944 13652 47984
rect 13996 49372 14036 49412
rect 13900 48700 13940 48740
rect 14188 49372 14228 49412
rect 14188 48616 14228 48656
rect 14092 48112 14132 48152
rect 13900 47944 13940 47984
rect 13804 47272 13844 47312
rect 14092 46852 14132 46892
rect 13900 45928 13940 45968
rect 13804 45004 13844 45044
rect 14092 45760 14132 45800
rect 14476 53320 14516 53360
rect 15724 67600 15764 67640
rect 15724 67180 15764 67220
rect 15628 66844 15668 66884
rect 15532 65416 15572 65456
rect 15436 65332 15476 65372
rect 15148 64240 15188 64280
rect 14956 63904 14996 63944
rect 16108 79360 16148 79400
rect 16108 79024 16148 79064
rect 16012 78184 16052 78224
rect 16012 77764 16052 77804
rect 16300 80284 16340 80324
rect 16492 79444 16532 79484
rect 16396 79360 16436 79400
rect 16972 85576 17012 85616
rect 17356 84484 17396 84524
rect 18028 85408 18068 85448
rect 17932 85072 17972 85112
rect 17740 84568 17780 84608
rect 17164 84400 17204 84440
rect 17548 84400 17588 84440
rect 18316 84484 18356 84524
rect 19084 85912 19124 85952
rect 19276 85912 19316 85952
rect 19276 85744 19316 85784
rect 18892 84904 18932 84944
rect 18808 84652 18848 84692
rect 18890 84652 18930 84692
rect 18972 84652 19012 84692
rect 19054 84652 19094 84692
rect 19136 84652 19176 84692
rect 18700 84484 18740 84524
rect 18124 84400 18164 84440
rect 18508 84400 18548 84440
rect 19564 85408 19604 85448
rect 19468 84400 19508 84440
rect 19276 83728 19316 83768
rect 19852 84736 19892 84776
rect 16684 80368 16724 80408
rect 16876 79360 16916 79400
rect 16300 77764 16340 77804
rect 16204 77680 16244 77720
rect 16588 79024 16628 79064
rect 16396 77428 16436 77468
rect 17068 77680 17108 77720
rect 17740 77680 17780 77720
rect 16204 76924 16244 76964
rect 16108 76672 16148 76712
rect 16108 75916 16148 75956
rect 16012 75496 16052 75536
rect 16012 75328 16052 75368
rect 15916 72976 15956 73016
rect 15916 71464 15956 71504
rect 16684 76840 16724 76880
rect 16204 75244 16244 75284
rect 16108 74404 16148 74444
rect 16108 74152 16148 74192
rect 16300 73816 16340 73856
rect 16204 73564 16244 73604
rect 16300 73060 16340 73100
rect 16780 76504 16820 76544
rect 17260 77428 17300 77468
rect 17740 76924 17780 76964
rect 17548 76840 17588 76880
rect 16972 76168 17012 76208
rect 17452 76588 17492 76628
rect 17068 75748 17108 75788
rect 17068 75580 17108 75620
rect 17260 75580 17300 75620
rect 16876 75244 16916 75284
rect 16972 75160 17012 75200
rect 16972 74404 17012 74444
rect 16588 73648 16628 73688
rect 16108 71968 16148 72008
rect 16204 70624 16244 70664
rect 16108 70540 16148 70580
rect 16396 72304 16436 72344
rect 16108 69868 16148 69908
rect 16204 69784 16244 69824
rect 16108 69196 16148 69236
rect 16204 68188 16244 68228
rect 15916 67852 15956 67892
rect 16300 67516 16340 67556
rect 15916 67264 15956 67304
rect 16396 67264 16436 67304
rect 15820 66844 15860 66884
rect 15724 64576 15764 64616
rect 14860 63820 14900 63860
rect 15628 63820 15668 63860
rect 14764 62224 14804 62264
rect 15148 63064 15188 63104
rect 15532 63064 15572 63104
rect 15052 62980 15092 63020
rect 15052 62812 15092 62852
rect 14956 62224 14996 62264
rect 14956 60796 14996 60836
rect 14860 60712 14900 60752
rect 14668 60544 14708 60584
rect 14668 60376 14708 60416
rect 14668 59956 14708 59996
rect 15628 62308 15668 62348
rect 15628 61720 15668 61760
rect 15148 61048 15188 61088
rect 15052 60376 15092 60416
rect 15628 60124 15668 60164
rect 15052 60040 15092 60080
rect 15436 60040 15476 60080
rect 14764 58192 14804 58232
rect 14668 57856 14708 57896
rect 14956 57100 14996 57140
rect 14668 56932 14708 56972
rect 14668 56512 14708 56552
rect 14668 56344 14708 56384
rect 14668 56092 14708 56132
rect 14668 53908 14708 53948
rect 14860 54328 14900 54368
rect 14764 52732 14804 52772
rect 14668 51724 14708 51764
rect 14860 51724 14900 51764
rect 14572 50968 14612 51008
rect 14572 50800 14612 50840
rect 14476 50548 14516 50588
rect 14380 49708 14420 49748
rect 14380 49540 14420 49580
rect 14284 48196 14324 48236
rect 14284 47860 14324 47900
rect 14476 49456 14516 49496
rect 14380 46768 14420 46808
rect 14764 50380 14804 50420
rect 14956 50044 14996 50084
rect 15436 59368 15476 59408
rect 15820 61300 15860 61340
rect 16300 65584 16340 65624
rect 16300 64576 16340 64616
rect 16300 61888 16340 61928
rect 16204 61552 16244 61592
rect 16204 60544 16244 60584
rect 16108 60040 16148 60080
rect 16012 59956 16052 59996
rect 15916 59620 15956 59660
rect 16113 59620 16153 59660
rect 15340 58780 15380 58820
rect 15244 57856 15284 57896
rect 15436 56848 15476 56888
rect 15724 59116 15764 59156
rect 15628 58192 15668 58232
rect 15628 58024 15668 58064
rect 15916 59368 15956 59408
rect 16204 58948 16244 58988
rect 16012 58024 16052 58064
rect 15628 57436 15668 57476
rect 15628 57016 15668 57056
rect 15148 54160 15188 54200
rect 15340 54160 15380 54200
rect 15148 53824 15188 53864
rect 15340 53908 15380 53948
rect 15724 55840 15764 55880
rect 15820 55588 15860 55628
rect 15724 55504 15764 55544
rect 15244 53488 15284 53528
rect 15148 51808 15188 51848
rect 15148 50632 15188 50672
rect 14764 49708 14804 49748
rect 14668 49540 14708 49580
rect 14764 46684 14804 46724
rect 14572 46348 14612 46388
rect 13708 44836 13748 44876
rect 13900 44668 13940 44708
rect 13804 44584 13844 44624
rect 13708 44500 13748 44540
rect 13228 43996 13268 44036
rect 12844 43324 12884 43364
rect 12748 43240 12788 43280
rect 12748 42736 12788 42776
rect 12844 41980 12884 42020
rect 12748 41896 12788 41936
rect 12652 40384 12692 40424
rect 12652 40132 12692 40172
rect 12460 39712 12500 39752
rect 12556 39544 12596 39584
rect 12460 39040 12500 39080
rect 12076 38368 12116 38408
rect 11884 38032 11924 38072
rect 11884 37360 11924 37400
rect 11788 37276 11828 37316
rect 11692 36268 11732 36308
rect 11692 35932 11732 35972
rect 12172 37276 12212 37316
rect 12364 36520 12404 36560
rect 11980 36184 12020 36224
rect 12172 36016 12212 36056
rect 11980 35848 12020 35888
rect 13420 44164 13460 44204
rect 13420 43576 13460 43616
rect 13324 43408 13364 43448
rect 13228 43324 13268 43364
rect 13228 42736 13268 42776
rect 13036 41980 13076 42020
rect 12940 40216 12980 40256
rect 12844 39964 12884 40004
rect 13996 44584 14036 44624
rect 14092 44500 14132 44540
rect 14284 44416 14324 44456
rect 14380 44248 14420 44288
rect 14284 44164 14324 44204
rect 13996 43912 14036 43952
rect 14188 43912 14228 43952
rect 14092 43576 14132 43616
rect 13612 43240 13652 43280
rect 14476 43408 14516 43448
rect 14380 43240 14420 43280
rect 13996 42736 14036 42776
rect 14764 46012 14804 46052
rect 15052 49540 15092 49580
rect 15244 49708 15284 49748
rect 15244 49456 15284 49496
rect 15436 53572 15476 53612
rect 16108 55504 16148 55544
rect 15916 55168 15956 55208
rect 15916 55000 15956 55040
rect 15628 53824 15668 53864
rect 15628 53656 15668 53696
rect 15532 51640 15572 51680
rect 15532 51388 15572 51428
rect 15820 53320 15860 53360
rect 15724 53152 15764 53192
rect 15628 50716 15668 50756
rect 15820 52900 15860 52940
rect 16012 53908 16052 53948
rect 16300 57940 16340 57980
rect 16300 57016 16340 57056
rect 16972 72304 17012 72344
rect 16684 71464 16724 71504
rect 16588 69952 16628 69992
rect 16876 69112 16916 69152
rect 16684 68944 16724 68984
rect 16972 68944 17012 68984
rect 16588 68440 16628 68480
rect 16972 68272 17012 68312
rect 16780 68020 16820 68060
rect 16588 67600 16628 67640
rect 16972 67684 17012 67724
rect 16684 67516 16724 67556
rect 16780 67264 16820 67304
rect 16876 67180 16916 67220
rect 16684 67012 16724 67052
rect 16876 66928 16916 66968
rect 16588 66676 16628 66716
rect 17260 74320 17300 74360
rect 17164 74068 17204 74108
rect 17164 73060 17204 73100
rect 17260 72808 17300 72848
rect 17260 71968 17300 72008
rect 17164 71296 17204 71336
rect 17164 70792 17204 70832
rect 17164 70540 17204 70580
rect 17356 71548 17396 71588
rect 17644 76168 17684 76208
rect 17548 76000 17588 76040
rect 17548 75748 17588 75788
rect 17740 75580 17780 75620
rect 17452 71464 17492 71504
rect 17356 70792 17396 70832
rect 17356 70624 17396 70664
rect 18988 83308 19028 83348
rect 18808 83140 18848 83180
rect 18890 83140 18930 83180
rect 18972 83140 19012 83180
rect 19054 83140 19094 83180
rect 19136 83140 19176 83180
rect 19660 83392 19700 83432
rect 19468 83308 19508 83348
rect 18988 82804 19028 82844
rect 19372 81712 19412 81752
rect 18808 81628 18848 81668
rect 18890 81628 18930 81668
rect 18972 81628 19012 81668
rect 19054 81628 19094 81668
rect 19136 81628 19176 81668
rect 19084 81460 19124 81500
rect 18988 81124 19028 81164
rect 18892 81040 18932 81080
rect 18412 78268 18452 78308
rect 19180 81376 19220 81416
rect 19372 81292 19412 81332
rect 19660 82300 19700 82340
rect 19564 81712 19604 81752
rect 19660 81376 19700 81416
rect 19276 80704 19316 80744
rect 19180 80536 19220 80576
rect 19084 80284 19124 80324
rect 18808 80116 18848 80156
rect 18890 80116 18930 80156
rect 18972 80116 19012 80156
rect 19054 80116 19094 80156
rect 19136 80116 19176 80156
rect 19468 80536 19508 80576
rect 19372 80200 19412 80240
rect 19372 79948 19412 79988
rect 18988 79780 19028 79820
rect 19276 79696 19316 79736
rect 19180 79360 19220 79400
rect 19276 79108 19316 79148
rect 18700 79024 18740 79064
rect 18988 78772 19028 78812
rect 18808 78604 18848 78644
rect 18890 78604 18930 78644
rect 18972 78604 19012 78644
rect 19054 78604 19094 78644
rect 19136 78604 19176 78644
rect 19180 78436 19220 78476
rect 18508 77512 18548 77552
rect 18988 78268 19028 78308
rect 19372 78100 19412 78140
rect 19276 77596 19316 77636
rect 18988 77428 19028 77468
rect 19564 80032 19604 80072
rect 19756 80452 19796 80492
rect 19660 79696 19700 79736
rect 19564 78772 19604 78812
rect 19756 79528 19796 79568
rect 20524 84400 20564 84440
rect 20048 83896 20088 83936
rect 20130 83896 20170 83936
rect 20212 83896 20252 83936
rect 20294 83896 20334 83936
rect 20376 83896 20416 83936
rect 20048 82384 20088 82424
rect 20130 82384 20170 82424
rect 20212 82384 20252 82424
rect 20294 82384 20334 82424
rect 20376 82384 20416 82424
rect 19948 81376 19988 81416
rect 20048 80872 20088 80912
rect 20130 80872 20170 80912
rect 20212 80872 20252 80912
rect 20294 80872 20334 80912
rect 20376 80872 20416 80912
rect 19948 79696 19988 79736
rect 19852 79192 19892 79232
rect 19660 78688 19700 78728
rect 19564 78352 19604 78392
rect 20048 79360 20088 79400
rect 20130 79360 20170 79400
rect 20212 79360 20252 79400
rect 20294 79360 20334 79400
rect 20376 79360 20416 79400
rect 19948 78520 19988 78560
rect 19660 77680 19700 77720
rect 19084 77260 19124 77300
rect 18808 77092 18848 77132
rect 18890 77092 18930 77132
rect 18972 77092 19012 77132
rect 19054 77092 19094 77132
rect 19136 77092 19176 77132
rect 18124 76504 18164 76544
rect 18220 76000 18260 76040
rect 18028 74572 18068 74612
rect 18220 75244 18260 75284
rect 18604 76756 18644 76796
rect 18796 76672 18836 76712
rect 18700 76588 18740 76628
rect 18988 76420 19028 76460
rect 19180 76168 19220 76208
rect 19372 76420 19412 76460
rect 19468 76336 19508 76376
rect 19852 77428 19892 77468
rect 20048 77848 20088 77888
rect 20130 77848 20170 77888
rect 20212 77848 20252 77888
rect 20294 77848 20334 77888
rect 20376 77848 20416 77888
rect 20044 77008 20084 77048
rect 19852 76756 19892 76796
rect 19756 76252 19796 76292
rect 19372 76084 19412 76124
rect 19660 76084 19700 76124
rect 18808 75580 18848 75620
rect 18890 75580 18930 75620
rect 18972 75580 19012 75620
rect 19054 75580 19094 75620
rect 19136 75580 19176 75620
rect 18508 75412 18548 75452
rect 18796 75244 18836 75284
rect 18124 73228 18164 73268
rect 17932 73060 17972 73100
rect 18604 74992 18644 75032
rect 18604 74740 18644 74780
rect 18604 73648 18644 73688
rect 19084 74992 19124 75032
rect 19554 75832 19594 75872
rect 19564 75664 19604 75704
rect 19756 75748 19796 75788
rect 19948 76504 19988 76544
rect 20140 76504 20180 76544
rect 19948 76336 19988 76376
rect 20048 76336 20088 76376
rect 20130 76336 20170 76376
rect 20212 76336 20252 76376
rect 20294 76336 20334 76376
rect 20376 76336 20416 76376
rect 19948 75916 19988 75956
rect 20044 75664 20084 75704
rect 20044 75496 20084 75536
rect 19852 75076 19892 75116
rect 20140 74992 20180 75032
rect 19852 74404 19892 74444
rect 18808 74068 18848 74108
rect 18890 74068 18930 74108
rect 18972 74068 19012 74108
rect 19054 74068 19094 74108
rect 19136 74068 19176 74108
rect 19276 74068 19316 74108
rect 18892 73900 18932 73940
rect 18412 73564 18452 73604
rect 18700 73564 18740 73604
rect 19180 73648 19220 73688
rect 18988 73060 19028 73100
rect 17836 72052 17876 72092
rect 17740 71800 17780 71840
rect 17740 70960 17780 71000
rect 17644 70792 17684 70832
rect 17356 70204 17396 70244
rect 17260 69784 17300 69824
rect 17740 70540 17780 70580
rect 17740 69952 17780 69992
rect 17932 70624 17972 70664
rect 17932 69952 17972 69992
rect 17356 68944 17396 68984
rect 17836 69280 17876 69320
rect 17740 69196 17780 69236
rect 17740 68944 17780 68984
rect 17740 68440 17780 68480
rect 17932 68440 17972 68480
rect 17260 67936 17300 67976
rect 17260 67684 17300 67724
rect 17260 67348 17300 67388
rect 17644 68104 17684 68144
rect 17548 67600 17588 67640
rect 17068 66676 17108 66716
rect 16684 66088 16724 66128
rect 16684 65584 16724 65624
rect 16684 64576 16724 64616
rect 16876 65920 16916 65960
rect 16492 62560 16532 62600
rect 16780 62980 16820 63020
rect 16780 62560 16820 62600
rect 16588 61300 16628 61340
rect 16588 60712 16628 60752
rect 16684 60544 16724 60584
rect 16588 60040 16628 60080
rect 16396 56596 16436 56636
rect 16492 56260 16532 56300
rect 16492 55756 16532 55796
rect 16300 55000 16340 55040
rect 16204 53824 16244 53864
rect 16108 53572 16148 53612
rect 16108 52816 16148 52856
rect 15916 52060 15956 52100
rect 15916 51892 15956 51932
rect 15724 50632 15764 50672
rect 15532 50464 15572 50504
rect 15724 50464 15764 50504
rect 15436 50380 15476 50420
rect 15628 50296 15668 50336
rect 15532 50128 15572 50168
rect 15340 49204 15380 49244
rect 14956 48700 14996 48740
rect 16396 53656 16436 53696
rect 17068 65416 17108 65456
rect 17356 66088 17396 66128
rect 17548 66088 17588 66128
rect 17068 64576 17108 64616
rect 16972 64492 17012 64532
rect 17932 67936 17972 67976
rect 18412 72976 18452 73016
rect 18124 72808 18164 72848
rect 18124 70036 18164 70076
rect 18604 72556 18644 72596
rect 18412 71968 18452 72008
rect 18988 72892 19028 72932
rect 18796 72808 18836 72848
rect 19180 72808 19220 72848
rect 18808 72556 18848 72596
rect 18890 72556 18930 72596
rect 18972 72556 19012 72596
rect 19054 72556 19094 72596
rect 19136 72556 19176 72596
rect 18796 72388 18836 72428
rect 18988 72388 19028 72428
rect 19372 73144 19412 73184
rect 19756 74236 19796 74276
rect 20048 74824 20088 74864
rect 20130 74824 20170 74864
rect 20212 74824 20252 74864
rect 20294 74824 20334 74864
rect 20376 74824 20416 74864
rect 20044 74236 20084 74276
rect 19948 73900 19988 73940
rect 19564 72976 19604 73016
rect 19468 72640 19508 72680
rect 18220 69784 18260 69824
rect 18124 69700 18164 69740
rect 18124 68608 18164 68648
rect 18508 71800 18548 71840
rect 18124 68020 18164 68060
rect 17932 66088 17972 66128
rect 17644 65584 17684 65624
rect 17740 65500 17780 65540
rect 17740 64660 17780 64700
rect 17932 65584 17972 65624
rect 18412 68440 18452 68480
rect 19372 72220 19412 72260
rect 18892 71716 18932 71756
rect 19756 73732 19796 73772
rect 20048 73312 20088 73352
rect 20130 73312 20170 73352
rect 20212 73312 20252 73352
rect 20294 73312 20334 73352
rect 20376 73312 20416 73352
rect 19756 72724 19796 72764
rect 19660 72304 19700 72344
rect 19756 72220 19796 72260
rect 19564 71968 19604 72008
rect 19468 71632 19508 71672
rect 18988 71296 19028 71336
rect 18892 71212 18932 71252
rect 18808 71044 18848 71084
rect 18890 71044 18930 71084
rect 18972 71044 19012 71084
rect 19054 71044 19094 71084
rect 19136 71044 19176 71084
rect 19180 70876 19220 70916
rect 19372 71212 19412 71252
rect 19660 71296 19700 71336
rect 19756 70708 19796 70748
rect 19372 70204 19412 70244
rect 18808 69532 18848 69572
rect 18890 69532 18930 69572
rect 18972 69532 19012 69572
rect 19054 69532 19094 69572
rect 19136 69532 19176 69572
rect 19660 70036 19700 70076
rect 19468 69364 19508 69404
rect 19372 69280 19412 69320
rect 18892 69112 18932 69152
rect 18700 69028 18740 69068
rect 18892 68524 18932 68564
rect 18700 68440 18740 68480
rect 19756 69448 19796 69488
rect 19756 69280 19796 69320
rect 19564 68356 19604 68396
rect 19084 68272 19124 68312
rect 19372 68272 19412 68312
rect 18808 68020 18848 68060
rect 18890 68020 18930 68060
rect 18972 68020 19012 68060
rect 19054 68020 19094 68060
rect 19136 68020 19176 68060
rect 18508 67684 18548 67724
rect 18124 65668 18164 65708
rect 18316 65500 18356 65540
rect 18124 65451 18164 65456
rect 18124 65416 18164 65451
rect 18124 64324 18164 64364
rect 17260 63232 17300 63272
rect 17644 63232 17684 63272
rect 16972 63148 17012 63188
rect 17164 63064 17204 63104
rect 17164 62896 17204 62936
rect 16876 59956 16916 59996
rect 16972 59620 17012 59660
rect 16876 59536 16916 59576
rect 17164 60628 17204 60668
rect 17548 63064 17588 63104
rect 17260 60544 17300 60584
rect 17644 62896 17684 62936
rect 18028 64156 18068 64196
rect 17932 63736 17972 63776
rect 18028 63316 18068 63356
rect 18028 63064 18068 63104
rect 17740 62392 17780 62432
rect 17452 61300 17492 61340
rect 17356 60460 17396 60500
rect 17164 60292 17204 60332
rect 17452 60292 17492 60332
rect 17068 59032 17108 59072
rect 16972 58780 17012 58820
rect 16780 58528 16820 58568
rect 16780 57856 16820 57896
rect 16684 56932 16724 56972
rect 16684 56512 16724 56552
rect 17260 60040 17300 60080
rect 17644 59956 17684 59996
rect 17260 59116 17300 59156
rect 17164 58024 17204 58064
rect 17548 59032 17588 59072
rect 17836 61048 17876 61088
rect 18028 62392 18068 62432
rect 18220 60460 18260 60500
rect 18124 60292 18164 60332
rect 18220 59872 18260 59912
rect 18124 59704 18164 59744
rect 17644 58528 17684 58568
rect 17548 58108 17588 58148
rect 18028 57940 18068 57980
rect 16876 56764 16916 56804
rect 16780 56344 16820 56384
rect 16972 56344 17012 56384
rect 16876 56260 16916 56300
rect 17548 57856 17588 57896
rect 17644 57772 17684 57812
rect 17164 57688 17204 57728
rect 17548 56932 17588 56972
rect 17836 57856 17876 57896
rect 18124 57772 18164 57812
rect 17740 57688 17780 57728
rect 17740 57520 17780 57560
rect 18124 57268 18164 57308
rect 17932 57184 17972 57224
rect 18028 57100 18068 57140
rect 18508 66928 18548 66968
rect 19660 67600 19700 67640
rect 18808 66508 18848 66548
rect 18890 66508 18930 66548
rect 18972 66508 19012 66548
rect 19054 66508 19094 66548
rect 19136 66508 19176 66548
rect 19756 67096 19796 67136
rect 19948 72220 19988 72260
rect 20048 71800 20088 71840
rect 20130 71800 20170 71840
rect 20212 71800 20252 71840
rect 20294 71800 20334 71840
rect 20376 71800 20416 71840
rect 19948 71380 19988 71420
rect 19948 70792 19988 70832
rect 20044 70624 20084 70664
rect 20140 70540 20180 70580
rect 20048 70288 20088 70328
rect 20130 70288 20170 70328
rect 20212 70288 20252 70328
rect 20294 70288 20334 70328
rect 20376 70288 20416 70328
rect 20044 70036 20084 70076
rect 20140 69700 20180 69740
rect 20044 69616 20084 69656
rect 20044 69448 20084 69488
rect 19948 69112 19988 69152
rect 20044 68944 20084 68984
rect 20048 68776 20088 68816
rect 20130 68776 20170 68816
rect 20212 68776 20252 68816
rect 20294 68776 20334 68816
rect 20376 68776 20416 68816
rect 20044 68272 20084 68312
rect 19948 67936 19988 67976
rect 20140 67432 20180 67472
rect 20048 67264 20088 67304
rect 20130 67264 20170 67304
rect 20212 67264 20252 67304
rect 20294 67264 20334 67304
rect 20376 67264 20416 67304
rect 20620 84064 20660 84104
rect 21388 82720 21428 82760
rect 21388 82216 21428 82256
rect 20620 80536 20660 80576
rect 20620 76504 20660 76544
rect 20716 75748 20756 75788
rect 20620 75328 20660 75368
rect 20716 74320 20756 74360
rect 20620 72052 20660 72092
rect 20620 70960 20660 71000
rect 21388 70792 21428 70832
rect 20620 69700 20660 69740
rect 21388 68944 21428 68984
rect 20620 67936 20660 67976
rect 19948 66928 19988 66968
rect 19468 66592 19508 66632
rect 19180 65920 19220 65960
rect 19372 65500 19412 65540
rect 18700 65416 18740 65456
rect 19660 66256 19700 66296
rect 19948 66256 19988 66296
rect 19756 66172 19796 66212
rect 19564 65920 19604 65960
rect 18988 65248 19028 65288
rect 18808 64996 18848 65036
rect 18890 64996 18930 65036
rect 18972 64996 19012 65036
rect 19054 64996 19094 65036
rect 19136 64996 19176 65036
rect 19276 64912 19316 64952
rect 18988 64492 19028 64532
rect 18604 64156 18644 64196
rect 19756 65332 19796 65372
rect 20048 65752 20088 65792
rect 20130 65752 20170 65792
rect 20212 65752 20252 65792
rect 20294 65752 20334 65792
rect 20376 65752 20416 65792
rect 19948 65584 19988 65624
rect 20044 65248 20084 65288
rect 19852 64828 19892 64868
rect 19564 64576 19604 64616
rect 19660 64492 19700 64532
rect 19468 64072 19508 64112
rect 19372 63988 19412 64028
rect 18508 63904 18548 63944
rect 18508 62980 18548 63020
rect 19564 63904 19604 63944
rect 18808 63484 18848 63524
rect 18890 63484 18930 63524
rect 18972 63484 19012 63524
rect 19054 63484 19094 63524
rect 19136 63484 19176 63524
rect 19756 64408 19796 64448
rect 19948 64240 19988 64280
rect 20048 64240 20088 64280
rect 20130 64240 20170 64280
rect 20212 64240 20252 64280
rect 20294 64240 20334 64280
rect 20376 64240 20416 64280
rect 19756 63820 19796 63860
rect 19948 63568 19988 63608
rect 18508 62224 18548 62264
rect 19660 63232 19700 63272
rect 19660 62644 19700 62684
rect 18700 62224 18740 62264
rect 18604 61804 18644 61844
rect 18808 61972 18848 62012
rect 18890 61972 18930 62012
rect 18972 61972 19012 62012
rect 19054 61972 19094 62012
rect 19136 61972 19176 62012
rect 19084 61720 19124 61760
rect 18604 61636 18644 61676
rect 18988 61048 19028 61088
rect 19180 61552 19220 61592
rect 18604 60712 18644 60752
rect 19180 60628 19220 60668
rect 18604 60544 18644 60584
rect 18508 59284 18548 59324
rect 18412 58696 18452 58736
rect 18316 58024 18356 58064
rect 18808 60460 18848 60500
rect 18890 60460 18930 60500
rect 18972 60460 19012 60500
rect 19054 60460 19094 60500
rect 19136 60460 19176 60500
rect 19852 62560 19892 62600
rect 20524 62896 20564 62936
rect 20048 62728 20088 62768
rect 20130 62728 20170 62768
rect 20212 62728 20252 62768
rect 20294 62728 20334 62768
rect 20376 62728 20416 62768
rect 20044 62308 20084 62348
rect 19564 61384 19604 61424
rect 19372 61132 19412 61172
rect 19948 61888 19988 61928
rect 19468 60880 19508 60920
rect 19372 60040 19412 60080
rect 19180 59536 19220 59576
rect 18808 58948 18848 58988
rect 18890 58948 18930 58988
rect 18972 58948 19012 58988
rect 19054 58948 19094 58988
rect 19136 58948 19176 58988
rect 19372 59284 19412 59324
rect 20048 61216 20088 61256
rect 20130 61216 20170 61256
rect 20212 61216 20252 61256
rect 20294 61216 20334 61256
rect 20376 61216 20416 61256
rect 20044 60796 20084 60836
rect 21004 60544 21044 60584
rect 20236 60208 20276 60248
rect 19756 59788 19796 59828
rect 19948 59872 19988 59912
rect 20048 59704 20088 59744
rect 20130 59704 20170 59744
rect 20212 59704 20252 59744
rect 20294 59704 20334 59744
rect 20376 59704 20416 59744
rect 19948 59536 19988 59576
rect 19852 59368 19892 59408
rect 19756 59284 19796 59324
rect 18796 58696 18836 58736
rect 18892 57940 18932 57980
rect 19084 57856 19124 57896
rect 18988 57772 19028 57812
rect 17740 56848 17780 56888
rect 17932 56848 17972 56888
rect 17356 56260 17396 56300
rect 17164 55756 17204 55796
rect 17452 55756 17492 55796
rect 16972 55504 17012 55544
rect 16684 54580 16724 54620
rect 16588 54160 16628 54200
rect 16684 54076 16724 54116
rect 17740 56344 17780 56384
rect 18028 56680 18068 56720
rect 18700 57604 18740 57644
rect 18808 57436 18848 57476
rect 18890 57436 18930 57476
rect 18972 57436 19012 57476
rect 19054 57436 19094 57476
rect 19136 57436 19176 57476
rect 19372 57100 19412 57140
rect 19276 57016 19316 57056
rect 19276 56848 19316 56888
rect 18988 56512 19028 56552
rect 18220 56008 18260 56048
rect 17548 55588 17588 55628
rect 17644 55504 17684 55544
rect 17452 54916 17492 54956
rect 16780 53656 16820 53696
rect 17548 54748 17588 54788
rect 17164 54580 17204 54620
rect 17836 55000 17876 55040
rect 17260 54160 17300 54200
rect 17164 53908 17204 53948
rect 17548 54160 17588 54200
rect 17452 53824 17492 53864
rect 17260 53656 17300 53696
rect 16972 53488 17012 53528
rect 17164 53488 17204 53528
rect 16684 53068 16724 53108
rect 16588 52984 16628 53024
rect 16684 52900 16724 52940
rect 16492 52648 16532 52688
rect 16588 52480 16628 52520
rect 16492 52396 16532 52436
rect 16300 52060 16340 52100
rect 16396 51976 16436 52016
rect 16300 51724 16340 51764
rect 16204 51640 16244 51680
rect 16396 51640 16436 51680
rect 16300 51556 16340 51596
rect 16204 50296 16244 50336
rect 15628 49204 15668 49244
rect 16012 49204 16052 49244
rect 15532 49120 15572 49160
rect 15052 48448 15092 48488
rect 14956 47944 14996 47984
rect 14956 47020 14996 47060
rect 14668 44584 14708 44624
rect 14668 44332 14708 44372
rect 14668 43828 14708 43868
rect 13228 41644 13268 41684
rect 13324 41476 13364 41516
rect 13516 41476 13556 41516
rect 13420 41392 13460 41432
rect 12940 39628 12980 39668
rect 13420 38704 13460 38744
rect 13036 38620 13076 38660
rect 13324 38200 13364 38240
rect 12844 38116 12884 38156
rect 13420 38116 13460 38156
rect 13324 37864 13364 37904
rect 12748 37780 12788 37820
rect 12844 37276 12884 37316
rect 12748 36688 12788 36728
rect 13516 37360 13556 37400
rect 13420 36940 13460 36980
rect 13324 36520 13364 36560
rect 13228 36436 13268 36476
rect 11788 35428 11828 35468
rect 12172 35176 12212 35216
rect 12076 35092 12116 35132
rect 11692 34924 11732 34964
rect 11980 34924 12020 34964
rect 11692 34504 11732 34544
rect 11980 34672 12020 34712
rect 12460 35512 12500 35552
rect 12364 34924 12404 34964
rect 12268 34672 12308 34712
rect 12652 35680 12692 35720
rect 12652 35428 12692 35468
rect 12844 34924 12884 34964
rect 12748 34336 12788 34376
rect 12940 34420 12980 34460
rect 12364 34168 12404 34208
rect 12460 34084 12500 34124
rect 12268 34000 12308 34040
rect 11788 33748 11828 33788
rect 12364 33748 12404 33788
rect 11404 32152 11444 32192
rect 10732 28876 10772 28916
rect 10732 27448 10772 27488
rect 10636 26440 10676 26480
rect 10636 23920 10676 23960
rect 10540 20056 10580 20096
rect 10828 25516 10868 25556
rect 10732 21568 10772 21608
rect 10732 20728 10772 20768
rect 11020 23752 11060 23792
rect 11020 23332 11060 23372
rect 10924 22072 10964 22112
rect 10924 21820 10964 21860
rect 11788 32740 11828 32780
rect 11692 30472 11732 30512
rect 11596 29800 11636 29840
rect 11596 29212 11636 29252
rect 11500 28708 11540 28748
rect 11308 28372 11348 28412
rect 11404 28288 11444 28328
rect 12172 33244 12212 33284
rect 11980 33076 12020 33116
rect 12748 34000 12788 34040
rect 12556 33916 12596 33956
rect 12652 33160 12692 33200
rect 12652 32404 12692 32444
rect 12940 33748 12980 33788
rect 13132 35092 13172 35132
rect 13900 41644 13940 41684
rect 13804 41392 13844 41432
rect 14476 41728 14516 41768
rect 14476 41224 14516 41264
rect 13996 40300 14036 40340
rect 14476 40216 14516 40256
rect 14380 39964 14420 40004
rect 14188 39124 14228 39164
rect 13996 39040 14036 39080
rect 13900 38620 13940 38660
rect 13804 36940 13844 36980
rect 13708 36604 13748 36644
rect 13612 35008 13652 35048
rect 13228 34924 13268 34964
rect 12844 33580 12884 33620
rect 12652 31564 12692 31604
rect 12364 31144 12404 31184
rect 11980 30052 12020 30092
rect 12172 29800 12212 29840
rect 11980 28708 12020 28748
rect 11884 28624 11924 28664
rect 11212 27448 11252 27488
rect 11308 26104 11348 26144
rect 11884 28120 11924 28160
rect 12364 29548 12404 29588
rect 12268 29212 12308 29252
rect 12940 32488 12980 32528
rect 12172 28288 12212 28328
rect 11788 26104 11828 26144
rect 11596 25852 11636 25892
rect 11500 25180 11540 25220
rect 11212 24424 11252 24464
rect 11596 24340 11636 24380
rect 11692 24088 11732 24128
rect 11308 23752 11348 23792
rect 11596 23584 11636 23624
rect 11308 23416 11348 23456
rect 11500 23416 11540 23456
rect 11212 23248 11252 23288
rect 11116 23080 11156 23120
rect 11116 21820 11156 21860
rect 11692 22996 11732 23036
rect 11404 21148 11444 21188
rect 10924 21064 10964 21104
rect 11020 20896 11060 20936
rect 10636 19972 10676 20012
rect 11596 20896 11636 20936
rect 12076 27616 12116 27656
rect 12172 27532 12212 27572
rect 12076 25936 12116 25976
rect 11980 24760 12020 24800
rect 12076 24676 12116 24716
rect 11884 22744 11924 22784
rect 12172 21400 12212 21440
rect 12076 21064 12116 21104
rect 11404 20812 11444 20852
rect 11212 20308 11252 20348
rect 11020 20140 11060 20180
rect 11980 20896 12020 20936
rect 11753 20743 11793 20768
rect 11753 20728 11793 20743
rect 12364 28120 12404 28160
rect 12364 27196 12404 27236
rect 12556 28624 12596 28664
rect 12652 28540 12692 28580
rect 12556 27532 12596 27572
rect 12556 27364 12596 27404
rect 12460 26944 12500 26984
rect 12364 26524 12404 26564
rect 12652 27196 12692 27236
rect 13708 34420 13748 34460
rect 13420 33244 13460 33284
rect 13228 33076 13268 33116
rect 13420 32992 13460 33032
rect 13612 32992 13652 33032
rect 13228 32908 13268 32948
rect 13516 32908 13556 32948
rect 13420 32656 13460 32696
rect 13804 33328 13844 33368
rect 13516 32488 13556 32528
rect 13708 32404 13748 32444
rect 13228 32320 13268 32360
rect 13324 32152 13364 32192
rect 13132 31480 13172 31520
rect 13420 31564 13460 31604
rect 13324 31480 13364 31520
rect 13036 28624 13076 28664
rect 13228 28624 13268 28664
rect 12940 28288 12980 28328
rect 12748 26692 12788 26732
rect 12844 26608 12884 26648
rect 12652 26356 12692 26396
rect 12556 25516 12596 25556
rect 12460 25432 12500 25472
rect 12844 26104 12884 26144
rect 12748 25684 12788 25724
rect 13132 25852 13172 25892
rect 12940 25600 12980 25640
rect 13036 25348 13076 25388
rect 12364 22408 12404 22448
rect 11500 20308 11540 20348
rect 11980 20308 12020 20348
rect 11788 20224 11828 20264
rect 10924 20056 10964 20096
rect 11404 20056 11444 20096
rect 11116 19972 11156 20012
rect 10732 19888 10772 19928
rect 10540 19804 10580 19844
rect 11500 19888 11540 19928
rect 10732 19636 10772 19676
rect 10444 19552 10484 19592
rect 9964 19300 10004 19340
rect 10060 19300 10100 19340
rect 9964 18880 10004 18920
rect 9868 18460 9908 18500
rect 9772 18376 9812 18416
rect 9676 17704 9716 17744
rect 9676 17032 9716 17072
rect 9964 17704 10004 17744
rect 9868 17032 9908 17072
rect 9580 16444 9620 16484
rect 9580 16024 9620 16064
rect 9580 15772 9620 15812
rect 9580 14848 9620 14888
rect 9580 14680 9620 14720
rect 9772 16444 9812 16484
rect 10156 18544 10196 18584
rect 10348 18544 10388 18584
rect 10156 18124 10196 18164
rect 11212 19552 11252 19592
rect 10540 18544 10580 18584
rect 10636 18376 10676 18416
rect 10924 18544 10964 18584
rect 10828 17872 10868 17912
rect 11020 17788 11060 17828
rect 10924 17704 10964 17744
rect 11212 18880 11252 18920
rect 11212 18712 11252 18752
rect 10636 17620 10676 17660
rect 10924 17452 10964 17492
rect 10924 16696 10964 16736
rect 10060 16444 10100 16484
rect 10732 16360 10772 16400
rect 9868 16024 9908 16064
rect 10156 15856 10196 15896
rect 9772 15772 9812 15812
rect 10060 15772 10100 15812
rect 9964 14848 10004 14888
rect 10540 15520 10580 15560
rect 10828 16192 10868 16232
rect 9388 14176 9428 14216
rect 9580 14092 9620 14132
rect 9772 13000 9812 13040
rect 9964 14512 10004 14552
rect 9964 14008 10004 14048
rect 9964 13504 10004 13544
rect 9868 12916 9908 12956
rect 9964 12748 10004 12788
rect 9580 12244 9620 12284
rect 9580 11488 9620 11528
rect 9292 11236 9332 11276
rect 9388 11068 9428 11108
rect 9580 10984 9620 11024
rect 9004 10228 9044 10268
rect 9004 9808 9044 9848
rect 8908 8464 8948 8504
rect 8812 8296 8852 8336
rect 8908 7960 8948 8000
rect 8716 7708 8756 7748
rect 8812 7540 8852 7580
rect 8716 4768 8756 4808
rect 7084 1996 7124 2036
rect 6700 1828 6740 1868
rect 7084 1324 7124 1364
rect 6508 1240 6548 1280
rect 6796 1240 6836 1280
rect 6700 1156 6740 1196
rect 6604 1072 6644 1112
rect 6412 904 6452 944
rect 6412 400 6452 440
rect 6220 148 6260 188
rect 7660 2332 7700 2372
rect 7276 2080 7316 2120
rect 7756 1996 7796 2036
rect 7276 1492 7316 1532
rect 7564 1408 7604 1448
rect 7468 1240 7508 1280
rect 7372 1156 7412 1196
rect 7084 484 7124 524
rect 6988 64 7028 104
rect 7948 1828 7988 1868
rect 8140 1828 8180 1868
rect 7852 904 7892 944
rect 8332 1660 8372 1700
rect 8812 2164 8852 2204
rect 9772 10228 9812 10268
rect 9772 9976 9812 10016
rect 10156 14008 10196 14048
rect 10348 12916 10388 12956
rect 10636 13168 10676 13208
rect 10636 12580 10676 12620
rect 10060 11992 10100 12032
rect 10060 11488 10100 11528
rect 9964 9472 10004 9512
rect 9676 9304 9716 9344
rect 9388 8800 9428 8840
rect 9292 8716 9332 8756
rect 9292 8464 9332 8504
rect 9196 8380 9236 8420
rect 9292 4432 9332 4472
rect 9580 8716 9620 8756
rect 9484 8296 9524 8336
rect 9004 1996 9044 2036
rect 10924 14680 10964 14720
rect 10828 14596 10868 14636
rect 10828 13000 10868 13040
rect 10252 11152 10292 11192
rect 10156 11068 10196 11108
rect 10252 10396 10292 10436
rect 10636 11908 10676 11948
rect 10540 10564 10580 10604
rect 10444 10228 10484 10268
rect 10348 10060 10388 10100
rect 9964 7876 10004 7916
rect 9676 7456 9716 7496
rect 9964 6952 10004 6992
rect 9964 6784 10004 6824
rect 9580 2500 9620 2540
rect 9388 1996 9428 2036
rect 9772 4096 9812 4136
rect 9676 1912 9716 1952
rect 8428 1492 8468 1532
rect 8140 1324 8180 1364
rect 8332 1240 8372 1280
rect 8236 1072 8276 1112
rect 8236 736 8276 776
rect 8524 904 8564 944
rect 8716 904 8756 944
rect 8908 1660 8948 1700
rect 8812 736 8852 776
rect 9196 904 9236 944
rect 9100 484 9140 524
rect 9388 1156 9428 1196
rect 10156 7456 10196 7496
rect 10156 6952 10196 6992
rect 10252 6280 10292 6320
rect 9772 1660 9812 1700
rect 9484 652 9524 692
rect 10444 4096 10484 4136
rect 10828 11656 10868 11696
rect 10828 11152 10868 11192
rect 11596 19468 11636 19508
rect 11692 19384 11732 19424
rect 11692 17620 11732 17660
rect 11884 17200 11924 17240
rect 11212 16612 11252 16652
rect 11308 16528 11348 16568
rect 11212 16360 11252 16400
rect 11116 16276 11156 16316
rect 11212 15856 11252 15896
rect 11116 14596 11156 14636
rect 11020 11656 11060 11696
rect 11020 11068 11060 11108
rect 10924 10984 10964 11024
rect 11596 16192 11636 16232
rect 11596 14932 11636 14972
rect 11308 14764 11348 14804
rect 11500 14680 11540 14720
rect 11404 14260 11444 14300
rect 11212 14008 11252 14048
rect 11404 13084 11444 13124
rect 11404 12748 11444 12788
rect 11308 12412 11348 12452
rect 11596 13924 11636 13964
rect 11308 12076 11348 12116
rect 11500 11992 11540 12032
rect 11212 11824 11252 11864
rect 11212 11152 11252 11192
rect 11308 11068 11348 11108
rect 11404 10984 11444 11024
rect 11212 10312 11252 10352
rect 10828 9976 10868 10016
rect 10924 9556 10964 9596
rect 11020 8968 11060 9008
rect 11404 10144 11444 10184
rect 11308 8800 11348 8840
rect 11212 8632 11252 8672
rect 11116 8128 11156 8168
rect 11596 11656 11636 11696
rect 11788 16024 11828 16064
rect 11884 14260 11924 14300
rect 11788 12748 11828 12788
rect 12076 17368 12116 17408
rect 12076 17032 12116 17072
rect 12364 20308 12404 20348
rect 12652 25096 12692 25136
rect 12652 23752 12692 23792
rect 12556 23500 12596 23540
rect 12652 22912 12692 22952
rect 13996 38536 14036 38576
rect 13996 38200 14036 38240
rect 14188 37780 14228 37820
rect 14284 37696 14324 37736
rect 14188 37360 14228 37400
rect 14092 36688 14132 36728
rect 14476 38116 14516 38156
rect 14380 36520 14420 36560
rect 14284 36100 14324 36140
rect 14092 35176 14132 35216
rect 14380 35176 14420 35216
rect 14668 42064 14708 42104
rect 14668 40132 14708 40172
rect 14668 39964 14708 40004
rect 14668 39040 14708 39080
rect 14668 38368 14708 38408
rect 14668 38200 14708 38240
rect 14572 37864 14612 37904
rect 14860 44584 14900 44624
rect 15148 46516 15188 46556
rect 15916 48196 15956 48236
rect 16012 47944 16052 47984
rect 15340 46432 15380 46472
rect 15052 46348 15092 46388
rect 15244 46348 15284 46388
rect 15340 46264 15380 46304
rect 15244 45844 15284 45884
rect 15628 45760 15668 45800
rect 15532 45508 15572 45548
rect 15244 45424 15284 45464
rect 15052 45256 15092 45296
rect 15244 45256 15284 45296
rect 15244 44416 15284 44456
rect 15148 44248 15188 44288
rect 15052 44164 15092 44204
rect 14956 43912 14996 43952
rect 14956 41980 14996 42020
rect 14860 41896 14900 41936
rect 15436 44248 15476 44288
rect 15340 43408 15380 43448
rect 15916 46348 15956 46388
rect 15820 45760 15860 45800
rect 15820 45424 15860 45464
rect 16396 51220 16436 51260
rect 16396 50212 16436 50252
rect 16396 49876 16436 49916
rect 16396 49204 16436 49244
rect 16300 48868 16340 48908
rect 16300 48448 16340 48488
rect 16492 48616 16532 48656
rect 16396 48112 16436 48152
rect 16204 47944 16244 47984
rect 16300 47440 16340 47480
rect 16204 46852 16244 46892
rect 16108 45928 16148 45968
rect 16012 45760 16052 45800
rect 16108 45508 16148 45548
rect 16684 52060 16724 52100
rect 17068 53320 17108 53360
rect 17068 53068 17108 53108
rect 16876 52816 16916 52856
rect 16972 52648 17012 52688
rect 16876 52144 16916 52184
rect 16780 51892 16820 51932
rect 16780 51556 16820 51596
rect 16684 50968 16724 51008
rect 17164 52648 17204 52688
rect 17068 52480 17108 52520
rect 17068 51724 17108 51764
rect 16780 48616 16820 48656
rect 16684 48280 16724 48320
rect 16972 50632 17012 50672
rect 17644 53992 17684 54032
rect 18412 55924 18452 55964
rect 18124 55000 18164 55040
rect 18808 55924 18848 55964
rect 18890 55924 18930 55964
rect 18972 55924 19012 55964
rect 19054 55924 19094 55964
rect 19136 55924 19176 55964
rect 18220 54160 18260 54200
rect 17932 53992 17972 54032
rect 17740 53488 17780 53528
rect 17740 52984 17780 53024
rect 17548 52816 17588 52856
rect 17548 52648 17588 52688
rect 18508 55000 18548 55040
rect 18316 53908 18356 53948
rect 18028 53320 18068 53360
rect 18808 54412 18848 54452
rect 18890 54412 18930 54452
rect 18972 54412 19012 54452
rect 19054 54412 19094 54452
rect 19136 54412 19176 54452
rect 18892 53992 18932 54032
rect 19756 58612 19796 58652
rect 19564 57352 19604 57392
rect 19660 57268 19700 57308
rect 19948 59116 19988 59156
rect 20716 58864 20756 58904
rect 20048 58192 20088 58232
rect 20130 58192 20170 58232
rect 20212 58192 20252 58232
rect 20294 58192 20334 58232
rect 20376 58192 20416 58232
rect 20716 58108 20756 58148
rect 20620 57856 20660 57896
rect 19948 57772 19988 57812
rect 20044 57688 20084 57728
rect 20236 57604 20276 57644
rect 19948 57184 19988 57224
rect 19564 57100 19604 57140
rect 19468 56932 19508 56972
rect 19948 57016 19988 57056
rect 19756 56932 19796 56972
rect 20048 56680 20088 56720
rect 20130 56680 20170 56720
rect 20212 56680 20252 56720
rect 20294 56680 20334 56720
rect 20376 56680 20416 56720
rect 19468 56370 19508 56384
rect 19468 56344 19508 56370
rect 19468 55756 19508 55796
rect 19372 55504 19412 55544
rect 19660 55504 19700 55544
rect 19564 55000 19604 55040
rect 19372 54748 19412 54788
rect 18412 53320 18452 53360
rect 18700 53320 18740 53360
rect 19276 53320 19316 53360
rect 18220 52900 18260 52940
rect 18028 52816 18068 52856
rect 18220 52732 18260 52772
rect 17356 51724 17396 51764
rect 17260 51556 17300 51596
rect 17164 51472 17204 51512
rect 17740 51724 17780 51764
rect 17548 51640 17588 51680
rect 17452 51136 17492 51176
rect 17356 50464 17396 50504
rect 16972 50212 17012 50252
rect 16972 49204 17012 49244
rect 16972 47944 17012 47984
rect 17356 50296 17396 50336
rect 17164 49456 17204 49496
rect 17644 50968 17684 51008
rect 17644 50716 17684 50756
rect 17548 50464 17588 50504
rect 17644 50128 17684 50168
rect 17644 49624 17684 49664
rect 17452 49540 17492 49580
rect 17548 49204 17588 49244
rect 17356 49120 17396 49160
rect 18028 52480 18068 52520
rect 18808 52900 18848 52940
rect 18890 52900 18930 52940
rect 18972 52900 19012 52940
rect 19054 52900 19094 52940
rect 19136 52900 19176 52940
rect 18700 52816 18740 52856
rect 18220 52396 18260 52436
rect 17932 52312 17972 52352
rect 18508 52312 18548 52352
rect 18316 51724 18356 51764
rect 18220 51640 18260 51680
rect 18028 51136 18068 51176
rect 17836 50800 17876 50840
rect 18220 50632 18260 50672
rect 18124 50128 18164 50168
rect 18124 49540 18164 49580
rect 18028 49288 18068 49328
rect 17548 48616 17588 48656
rect 17452 48280 17492 48320
rect 16588 47356 16628 47396
rect 16876 47356 16916 47396
rect 16684 47020 16724 47060
rect 16588 46348 16628 46388
rect 16588 46012 16628 46052
rect 16300 45172 16340 45212
rect 16780 46432 16820 46472
rect 16780 46264 16820 46304
rect 16780 45592 16820 45632
rect 16204 44416 16244 44456
rect 17068 46432 17108 46472
rect 17068 46264 17108 46304
rect 17068 45795 17108 45800
rect 17068 45760 17108 45795
rect 16972 45004 17012 45044
rect 17452 46432 17492 46472
rect 17260 46264 17300 46304
rect 17164 44416 17204 44456
rect 16780 44248 16820 44288
rect 15724 41980 15764 42020
rect 15916 42736 15956 42776
rect 16300 42736 16340 42776
rect 16300 41896 16340 41936
rect 16588 43408 16628 43448
rect 16876 43240 16916 43280
rect 16780 43156 16820 43196
rect 16684 42820 16724 42860
rect 16492 41896 16532 41936
rect 16396 41812 16436 41852
rect 15628 41728 15668 41768
rect 15436 41476 15476 41516
rect 14956 40468 14996 40508
rect 14860 40384 14900 40424
rect 15148 40300 15188 40340
rect 15052 40216 15092 40256
rect 14956 40132 14996 40172
rect 14860 39712 14900 39752
rect 15052 40048 15092 40088
rect 14956 38704 14996 38744
rect 14860 37612 14900 37652
rect 14956 35932 14996 35972
rect 13996 34168 14036 34208
rect 14572 34168 14612 34208
rect 14092 34084 14132 34124
rect 14092 33916 14132 33956
rect 14476 33580 14516 33620
rect 14284 33412 14324 33452
rect 14092 33244 14132 33284
rect 13996 32152 14036 32192
rect 14284 32152 14324 32192
rect 14380 32068 14420 32108
rect 13420 28540 13460 28580
rect 13708 29800 13748 29840
rect 13996 29800 14036 29840
rect 13900 29716 13940 29756
rect 13804 29044 13844 29084
rect 13804 28288 13844 28328
rect 13324 27532 13364 27572
rect 13516 26608 13556 26648
rect 14092 29296 14132 29336
rect 13996 29212 14036 29252
rect 13996 28288 14036 28328
rect 13996 27616 14036 27656
rect 13900 26608 13940 26648
rect 13804 26524 13844 26564
rect 13420 26440 13460 26480
rect 13708 26440 13748 26480
rect 13324 26356 13364 26396
rect 13612 26104 13652 26144
rect 13324 25684 13364 25724
rect 13228 25096 13268 25136
rect 12940 24928 12980 24968
rect 13036 24760 13076 24800
rect 13228 24760 13268 24800
rect 13516 25348 13556 25388
rect 13420 25264 13460 25304
rect 13804 25348 13844 25388
rect 14572 33244 14612 33284
rect 14956 35008 14996 35048
rect 15244 40132 15284 40172
rect 15532 39880 15572 39920
rect 15340 38116 15380 38156
rect 15148 37780 15188 37820
rect 15436 37696 15476 37736
rect 15436 37528 15476 37568
rect 15436 36688 15476 36728
rect 15340 36520 15380 36560
rect 15244 36100 15284 36140
rect 15244 35344 15284 35384
rect 15052 34420 15092 34460
rect 14956 34336 14996 34376
rect 14956 33244 14996 33284
rect 15436 35260 15476 35300
rect 15436 34504 15476 34544
rect 16108 41728 16148 41768
rect 15820 40552 15860 40592
rect 16012 40468 16052 40508
rect 15916 40389 15956 40424
rect 15916 40384 15956 40389
rect 15820 39628 15860 39668
rect 15724 38704 15764 38744
rect 16108 39880 16148 39920
rect 16108 39628 16148 39668
rect 15916 38536 15956 38576
rect 16108 38536 16148 38576
rect 16300 38704 16340 38744
rect 16492 38704 16532 38744
rect 16300 38536 16340 38576
rect 15820 37864 15860 37904
rect 15820 37696 15860 37736
rect 15916 37612 15956 37652
rect 15724 36688 15764 36728
rect 15916 36604 15956 36644
rect 15724 36436 15764 36476
rect 15628 35260 15668 35300
rect 15628 35008 15668 35048
rect 15244 33916 15284 33956
rect 14572 31228 14612 31268
rect 14572 30640 14612 30680
rect 14476 29296 14516 29336
rect 14380 28036 14420 28076
rect 14476 27868 14516 27908
rect 14572 27448 14612 27488
rect 14092 26524 14132 26564
rect 13996 26104 14036 26144
rect 14092 25348 14132 25388
rect 13996 25264 14036 25304
rect 14092 25096 14132 25136
rect 13516 24592 13556 24632
rect 12844 24424 12884 24464
rect 13516 24172 13556 24212
rect 13228 23920 13268 23960
rect 12844 23164 12884 23204
rect 13132 23164 13172 23204
rect 12748 22576 12788 22616
rect 13420 23080 13460 23120
rect 13036 22912 13076 22952
rect 12556 22492 12596 22532
rect 12940 22492 12980 22532
rect 13996 24340 14036 24380
rect 13612 23836 13652 23876
rect 13900 23836 13940 23876
rect 14092 24256 14132 24296
rect 13612 23080 13652 23120
rect 13228 22744 13268 22784
rect 13420 22744 13460 22784
rect 13132 22576 13172 22616
rect 12652 22324 12692 22364
rect 12556 21568 12596 21608
rect 12364 19384 12404 19424
rect 12556 19216 12596 19256
rect 12268 18880 12308 18920
rect 12172 15016 12212 15056
rect 12076 14596 12116 14636
rect 12172 14344 12212 14384
rect 12076 13168 12116 13208
rect 11788 12076 11828 12116
rect 11692 11068 11732 11108
rect 11596 10984 11636 11024
rect 11596 10648 11636 10688
rect 11596 10396 11636 10436
rect 10924 7456 10964 7496
rect 10924 7120 10964 7160
rect 11500 7876 11540 7916
rect 11884 11908 11924 11948
rect 12076 12244 12116 12284
rect 12652 19048 12692 19088
rect 12556 18376 12596 18416
rect 12460 17200 12500 17240
rect 12364 15016 12404 15056
rect 12364 13924 12404 13964
rect 12268 12412 12308 12452
rect 12172 11824 12212 11864
rect 12364 11740 12404 11780
rect 12172 11656 12212 11696
rect 12076 11572 12116 11612
rect 11980 10648 12020 10688
rect 11884 10312 11924 10352
rect 11692 9472 11732 9512
rect 11788 8800 11828 8840
rect 11692 8632 11732 8672
rect 11692 8044 11732 8084
rect 11500 6448 11540 6488
rect 11500 6280 11540 6320
rect 11788 7876 11828 7916
rect 11500 6028 11540 6068
rect 9868 1156 9908 1196
rect 10060 1660 10100 1700
rect 9964 820 10004 860
rect 9868 736 9908 776
rect 9772 232 9812 272
rect 10348 1156 10388 1196
rect 10252 736 10292 776
rect 10540 1828 10580 1868
rect 10924 1828 10964 1868
rect 10828 1408 10868 1448
rect 10732 1324 10772 1364
rect 10540 904 10580 944
rect 10636 820 10676 860
rect 11884 6028 11924 6068
rect 12076 8380 12116 8420
rect 12940 20896 12980 20936
rect 12844 20056 12884 20096
rect 12844 19720 12884 19760
rect 13132 22072 13172 22112
rect 13324 20896 13364 20936
rect 13132 20728 13172 20768
rect 13132 20392 13172 20432
rect 13036 20224 13076 20264
rect 13036 19720 13076 19760
rect 13228 20056 13268 20096
rect 13228 19384 13268 19424
rect 12844 19300 12884 19340
rect 13420 20728 13460 20768
rect 13516 19888 13556 19928
rect 13708 21904 13748 21944
rect 13804 21316 13844 21356
rect 13804 20392 13844 20432
rect 14284 25180 14324 25220
rect 14188 23248 14228 23288
rect 14092 21820 14132 21860
rect 14572 26440 14612 26480
rect 14476 25096 14516 25136
rect 14476 24592 14516 24632
rect 14764 31480 14804 31520
rect 14764 30808 14804 30848
rect 15148 32152 15188 32192
rect 14860 30136 14900 30176
rect 14860 29884 14900 29924
rect 14764 29716 14804 29756
rect 15052 30220 15092 30260
rect 15244 31480 15284 31520
rect 15340 31228 15380 31268
rect 15532 31312 15572 31352
rect 15532 30556 15572 30596
rect 15436 30304 15476 30344
rect 15340 29632 15380 29672
rect 15052 29380 15092 29420
rect 14956 29296 14996 29336
rect 14764 27196 14804 27236
rect 15244 29548 15284 29588
rect 15148 29212 15188 29252
rect 15052 28960 15092 29000
rect 15436 29464 15476 29504
rect 15340 29044 15380 29084
rect 14956 27112 14996 27152
rect 14860 26776 14900 26816
rect 14764 26692 14804 26732
rect 15244 28288 15284 28328
rect 15244 27532 15284 27572
rect 15244 26860 15284 26900
rect 15148 26776 15188 26816
rect 14956 26440 14996 26480
rect 15436 27868 15476 27908
rect 15820 35932 15860 35972
rect 15724 33832 15764 33872
rect 15724 33664 15764 33704
rect 15724 32320 15764 32360
rect 16396 38200 16436 38240
rect 15916 34336 15956 34376
rect 16300 37696 16340 37736
rect 16492 38116 16532 38156
rect 16396 36520 16436 36560
rect 16684 39712 16724 39752
rect 16588 37192 16628 37232
rect 16588 36772 16628 36812
rect 16588 35680 16628 35720
rect 16204 35176 16244 35216
rect 17260 44248 17300 44288
rect 17452 45508 17492 45548
rect 17164 43828 17204 43868
rect 17740 47944 17780 47984
rect 17644 47020 17684 47060
rect 17740 46348 17780 46388
rect 17740 46096 17780 46136
rect 17740 45508 17780 45548
rect 17644 44332 17684 44372
rect 17644 44164 17684 44204
rect 17548 42736 17588 42776
rect 17260 41896 17300 41936
rect 17164 40384 17204 40424
rect 17452 39712 17492 39752
rect 17260 38704 17300 38744
rect 18412 51640 18452 51680
rect 18412 50296 18452 50336
rect 18412 49288 18452 49328
rect 18796 52480 18836 52520
rect 18700 51892 18740 51932
rect 18604 51724 18644 51764
rect 18604 51556 18644 51596
rect 18604 49456 18644 49496
rect 18508 48952 18548 48992
rect 18808 51388 18848 51428
rect 18890 51388 18930 51428
rect 18972 51388 19012 51428
rect 19054 51388 19094 51428
rect 19136 51388 19176 51428
rect 18892 51220 18932 51260
rect 19468 53488 19508 53528
rect 19660 53320 19700 53360
rect 19468 53152 19508 53192
rect 19852 55756 19892 55796
rect 19852 55336 19892 55376
rect 20140 55336 20180 55376
rect 20048 55168 20088 55208
rect 20130 55168 20170 55208
rect 20212 55168 20252 55208
rect 20294 55168 20334 55208
rect 20376 55168 20416 55208
rect 19948 54832 19988 54872
rect 19852 54160 19892 54200
rect 19948 53992 19988 54032
rect 19852 53572 19892 53612
rect 20048 53656 20088 53696
rect 20130 53656 20170 53696
rect 20212 53656 20252 53696
rect 20294 53656 20334 53696
rect 20376 53656 20416 53696
rect 19756 53068 19796 53108
rect 19564 52984 19604 53024
rect 20236 53320 20276 53360
rect 20044 53068 20084 53108
rect 19948 52900 19988 52940
rect 19660 52732 19700 52772
rect 19852 52732 19892 52772
rect 19660 52480 19700 52520
rect 19948 52648 19988 52688
rect 20140 52565 20180 52604
rect 20140 52564 20180 52565
rect 20048 52144 20088 52184
rect 20130 52144 20170 52184
rect 20212 52144 20252 52184
rect 20294 52144 20334 52184
rect 20376 52144 20416 52184
rect 20140 51556 20180 51596
rect 19948 51220 19988 51260
rect 19564 51052 19604 51092
rect 19084 50968 19124 51008
rect 19372 50968 19412 51008
rect 20140 50800 20180 50840
rect 19948 50632 19988 50672
rect 20048 50632 20088 50672
rect 20130 50632 20170 50672
rect 20212 50632 20252 50672
rect 20294 50632 20334 50672
rect 20376 50632 20416 50672
rect 18988 50380 19028 50420
rect 18796 50128 18836 50168
rect 19180 50296 19220 50336
rect 19372 50296 19412 50336
rect 19372 50128 19412 50168
rect 18808 49876 18848 49916
rect 18890 49876 18930 49916
rect 18972 49876 19012 49916
rect 19054 49876 19094 49916
rect 19136 49876 19176 49916
rect 18892 48868 18932 48908
rect 19084 48868 19124 48908
rect 18700 48616 18740 48656
rect 18508 48448 18548 48488
rect 18604 48364 18644 48404
rect 18808 48364 18848 48404
rect 18890 48364 18930 48404
rect 18972 48364 19012 48404
rect 19054 48364 19094 48404
rect 19136 48364 19176 48404
rect 18412 48196 18452 48236
rect 18220 47944 18260 47984
rect 19372 49876 19412 49916
rect 19276 47944 19316 47984
rect 18124 47692 18164 47732
rect 18028 47272 18068 47312
rect 17932 46264 17972 46304
rect 19276 47104 19316 47144
rect 18604 47020 18644 47060
rect 18808 46852 18848 46892
rect 18890 46852 18930 46892
rect 18972 46852 19012 46892
rect 19054 46852 19094 46892
rect 19136 46852 19176 46892
rect 18604 46432 18644 46472
rect 19756 50128 19796 50168
rect 19660 50044 19700 50084
rect 19660 49876 19700 49916
rect 19852 49456 19892 49496
rect 19852 48952 19892 48992
rect 20140 50296 20180 50336
rect 21196 58192 21236 58232
rect 21004 57688 21044 57728
rect 20812 56176 20852 56216
rect 20812 55840 20852 55880
rect 20716 53320 20756 53360
rect 20812 52564 20852 52604
rect 20908 51472 20948 51512
rect 20812 51052 20852 51092
rect 20236 50212 20276 50252
rect 20620 50212 20660 50252
rect 20524 49960 20564 50000
rect 20044 49288 20084 49328
rect 20620 49792 20660 49832
rect 20048 49120 20088 49160
rect 20130 49120 20170 49160
rect 20212 49120 20252 49160
rect 20294 49120 20334 49160
rect 20376 49120 20416 49160
rect 20524 49120 20564 49160
rect 19468 48700 19508 48740
rect 19468 48280 19508 48320
rect 20044 48616 20084 48656
rect 20620 48616 20660 48656
rect 19852 48532 19892 48572
rect 19564 48196 19604 48236
rect 19564 48028 19604 48068
rect 18604 46264 18644 46304
rect 18124 46096 18164 46136
rect 18412 46096 18452 46136
rect 17932 45592 17972 45632
rect 18220 45760 18260 45800
rect 18028 45508 18068 45548
rect 18412 45424 18452 45464
rect 17932 45340 17972 45380
rect 17836 44080 17876 44120
rect 18316 44080 18356 44120
rect 18316 43912 18356 43952
rect 17932 43492 17972 43532
rect 18508 43912 18548 43952
rect 19948 47944 19988 47984
rect 19852 47860 19892 47900
rect 19852 46936 19892 46976
rect 20048 47608 20088 47648
rect 20130 47608 20170 47648
rect 20212 47608 20252 47648
rect 20294 47608 20334 47648
rect 20376 47608 20416 47648
rect 18808 45340 18848 45380
rect 18890 45340 18930 45380
rect 18972 45340 19012 45380
rect 19054 45340 19094 45380
rect 19136 45340 19176 45380
rect 18700 44416 18740 44456
rect 18988 45172 19028 45212
rect 18892 45004 18932 45044
rect 19468 44668 19508 44708
rect 19660 45508 19700 45548
rect 21388 56344 21428 56384
rect 21388 55840 21428 55880
rect 21196 51304 21236 51344
rect 20908 46600 20948 46640
rect 20044 46437 20084 46472
rect 20044 46432 20084 46437
rect 20236 46348 20276 46388
rect 19756 45004 19796 45044
rect 20048 46096 20088 46136
rect 20130 46096 20170 46136
rect 20212 46096 20252 46136
rect 20294 46096 20334 46136
rect 20376 46096 20416 46136
rect 20048 44584 20088 44624
rect 20130 44584 20170 44624
rect 20212 44584 20252 44624
rect 20294 44584 20334 44624
rect 20376 44584 20416 44624
rect 19948 44164 19988 44204
rect 18808 43828 18848 43868
rect 18890 43828 18930 43868
rect 18972 43828 19012 43868
rect 19054 43828 19094 43868
rect 19136 43828 19176 43868
rect 18316 43156 18356 43196
rect 20048 43072 20088 43112
rect 20130 43072 20170 43112
rect 20212 43072 20252 43112
rect 20294 43072 20334 43112
rect 20376 43072 20416 43112
rect 20236 42736 20276 42776
rect 19756 42568 19796 42608
rect 20044 42568 20084 42608
rect 19564 42484 19604 42524
rect 18124 42400 18164 42440
rect 17932 42064 17972 42104
rect 18124 41980 18164 42020
rect 17740 41896 17780 41936
rect 17836 40636 17876 40676
rect 18028 40384 18068 40424
rect 17644 38452 17684 38492
rect 17068 37276 17108 37316
rect 16972 36940 17012 36980
rect 16684 35344 16724 35384
rect 16108 32320 16148 32360
rect 16300 32152 16340 32192
rect 16972 36772 17012 36812
rect 17068 36604 17108 36644
rect 16972 36520 17012 36560
rect 16684 34840 16724 34880
rect 16876 34588 16916 34628
rect 16684 34420 16724 34460
rect 16972 34336 17012 34376
rect 17548 36940 17588 36980
rect 17356 35848 17396 35888
rect 18808 42316 18848 42356
rect 18890 42316 18930 42356
rect 18972 42316 19012 42356
rect 19054 42316 19094 42356
rect 19136 42316 19176 42356
rect 18700 41896 18740 41936
rect 18988 41896 19028 41936
rect 19468 41728 19508 41768
rect 19276 41140 19316 41180
rect 19468 41056 19508 41096
rect 19660 41980 19700 42020
rect 20524 42232 20564 42272
rect 19852 42064 19892 42104
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 19852 41392 19892 41432
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 19372 40720 19412 40760
rect 19564 40720 19604 40760
rect 19180 39964 19220 40004
rect 19564 39796 19604 39836
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 19276 38788 19316 38828
rect 18700 38704 18740 38744
rect 18988 38704 19028 38744
rect 18604 38116 18644 38156
rect 19276 38116 19316 38156
rect 18220 38032 18260 38072
rect 18220 37864 18260 37904
rect 18604 37864 18644 37904
rect 18124 36856 18164 36896
rect 18220 36772 18260 36812
rect 18124 35932 18164 35972
rect 17260 35008 17300 35048
rect 17164 34420 17204 34460
rect 17260 33244 17300 33284
rect 16492 32152 16532 32192
rect 16204 31480 16244 31520
rect 16204 30640 16244 30680
rect 16396 31060 16436 31100
rect 16204 30472 16244 30512
rect 15820 29968 15860 30008
rect 16300 29968 16340 30008
rect 15724 29632 15764 29672
rect 15916 29800 15956 29840
rect 15820 29464 15860 29504
rect 15916 29128 15956 29168
rect 15628 28624 15668 28664
rect 15532 27616 15572 27656
rect 15820 27784 15860 27824
rect 15436 27196 15476 27236
rect 16108 28288 16148 28328
rect 16108 28120 16148 28160
rect 15916 27448 15956 27488
rect 16300 29296 16340 29336
rect 16204 27364 16244 27404
rect 15724 26188 15764 26228
rect 15148 25516 15188 25556
rect 14764 24508 14804 24548
rect 14860 24424 14900 24464
rect 15244 24676 15284 24716
rect 14476 23752 14516 23792
rect 14476 23248 14516 23288
rect 15148 23920 15188 23960
rect 15436 25180 15476 25220
rect 15436 24760 15476 24800
rect 15340 23920 15380 23960
rect 15244 23584 15284 23624
rect 15244 22996 15284 23036
rect 14476 22492 14516 22532
rect 15148 22492 15188 22532
rect 14380 22240 14420 22280
rect 14572 22240 14612 22280
rect 14764 22240 14804 22280
rect 14284 21904 14324 21944
rect 14284 21736 14324 21776
rect 13708 19972 13748 20012
rect 12940 19048 12980 19088
rect 12844 18292 12884 18332
rect 12844 17872 12884 17912
rect 13708 19300 13748 19340
rect 13612 19048 13652 19088
rect 13324 18880 13364 18920
rect 13228 18544 13268 18584
rect 13228 18208 13268 18248
rect 13228 17620 13268 17660
rect 13132 17536 13172 17576
rect 12940 17368 12980 17408
rect 13132 17116 13172 17156
rect 13804 18880 13844 18920
rect 13900 18292 13940 18332
rect 13708 18040 13748 18080
rect 13516 17872 13556 17912
rect 13900 17704 13940 17744
rect 13516 17368 13556 17408
rect 13708 17200 13748 17240
rect 13516 16948 13556 16988
rect 12940 16108 12980 16148
rect 13036 16024 13076 16064
rect 13036 15604 13076 15644
rect 12844 15520 12884 15560
rect 12748 15184 12788 15224
rect 12652 12748 12692 12788
rect 12556 12412 12596 12452
rect 12844 15100 12884 15140
rect 12844 14008 12884 14048
rect 13420 15016 13460 15056
rect 13612 16696 13652 16736
rect 13804 17116 13844 17156
rect 13516 14932 13556 14972
rect 13708 16360 13748 16400
rect 13612 14764 13652 14804
rect 13132 13756 13172 13796
rect 12940 13084 12980 13124
rect 12940 12580 12980 12620
rect 12844 12412 12884 12452
rect 13036 12496 13076 12536
rect 13036 12076 13076 12116
rect 12940 11992 12980 12032
rect 12940 11320 12980 11360
rect 12748 11236 12788 11276
rect 12748 11068 12788 11108
rect 12652 10312 12692 10352
rect 12556 10144 12596 10184
rect 13036 11236 13076 11276
rect 13516 13168 13556 13208
rect 13420 11320 13460 11360
rect 12460 9472 12500 9512
rect 12556 9136 12596 9176
rect 12460 8632 12500 8672
rect 12460 8380 12500 8420
rect 12364 7288 12404 7328
rect 12076 6784 12116 6824
rect 12172 6448 12212 6488
rect 12076 6280 12116 6320
rect 12748 8044 12788 8084
rect 12652 7288 12692 7328
rect 12748 7120 12788 7160
rect 12460 5524 12500 5564
rect 12076 5104 12116 5144
rect 11980 2752 12020 2792
rect 11308 1660 11348 1700
rect 11884 2332 11924 2372
rect 11692 1828 11732 1868
rect 12076 1828 12116 1868
rect 11596 1156 11636 1196
rect 11212 1072 11252 1112
rect 11212 904 11252 944
rect 11884 1324 11924 1364
rect 12172 1240 12212 1280
rect 11980 1072 12020 1112
rect 11020 736 11060 776
rect 12556 988 12596 1028
rect 13036 9976 13076 10016
rect 12940 9556 12980 9596
rect 12940 8632 12980 8672
rect 12940 8380 12980 8420
rect 12748 5020 12788 5060
rect 13228 10816 13268 10856
rect 13132 7204 13172 7244
rect 13324 10732 13364 10772
rect 13324 8464 13364 8504
rect 14668 21904 14708 21944
rect 14572 21820 14612 21860
rect 15052 22240 15092 22280
rect 14860 21568 14900 21608
rect 14476 20644 14516 20684
rect 14188 19468 14228 19508
rect 14092 19300 14132 19340
rect 14188 19132 14228 19172
rect 14380 19048 14420 19088
rect 14092 17368 14132 17408
rect 14092 17200 14132 17240
rect 14092 15688 14132 15728
rect 14092 14932 14132 14972
rect 13996 14848 14036 14888
rect 13900 13672 13940 13712
rect 13516 9976 13556 10016
rect 13708 12748 13748 12788
rect 13612 9808 13652 9848
rect 13996 13168 14036 13208
rect 13996 12664 14036 12704
rect 13900 11404 13940 11444
rect 15436 22240 15476 22280
rect 15340 22072 15380 22112
rect 15820 25852 15860 25892
rect 15724 24760 15764 24800
rect 15724 24592 15764 24632
rect 16012 25096 16052 25136
rect 15916 24760 15956 24800
rect 16108 24844 16148 24884
rect 15820 24004 15860 24044
rect 16492 30220 16532 30260
rect 17356 32992 17396 33032
rect 16780 32656 16820 32696
rect 16780 32404 16820 32444
rect 16780 31144 16820 31184
rect 16684 31060 16724 31100
rect 16876 30640 16916 30680
rect 17356 32152 17396 32192
rect 17356 31648 17396 31688
rect 17548 34504 17588 34544
rect 17740 35848 17780 35888
rect 17740 35344 17780 35384
rect 17644 34168 17684 34208
rect 17548 34084 17588 34124
rect 18124 34336 18164 34376
rect 18028 34084 18068 34124
rect 17740 33832 17780 33872
rect 17548 32656 17588 32696
rect 17164 31396 17204 31436
rect 17452 31312 17492 31352
rect 17356 30976 17396 31016
rect 17260 30808 17300 30848
rect 16588 29884 16628 29924
rect 16588 29632 16628 29672
rect 16492 29128 16532 29168
rect 16588 28204 16628 28244
rect 17068 30220 17108 30260
rect 16780 29716 16820 29756
rect 16684 27952 16724 27992
rect 16684 27784 16724 27824
rect 17164 30052 17204 30092
rect 17068 29212 17108 29252
rect 16972 29044 17012 29084
rect 17068 28876 17108 28916
rect 16876 28120 16916 28160
rect 16396 26608 16436 26648
rect 16588 27196 16628 27236
rect 16684 26776 16724 26816
rect 16492 26524 16532 26564
rect 16684 26524 16724 26564
rect 16396 25768 16436 25808
rect 16300 25096 16340 25136
rect 16012 24340 16052 24380
rect 15916 23920 15956 23960
rect 16108 24004 16148 24044
rect 16204 23080 16244 23120
rect 15724 22492 15764 22532
rect 15724 22324 15764 22364
rect 15628 22072 15668 22112
rect 15340 21652 15380 21692
rect 15244 21568 15284 21608
rect 15436 21484 15476 21524
rect 15340 20896 15380 20936
rect 15148 20560 15188 20600
rect 15724 21484 15764 21524
rect 16012 22660 16052 22700
rect 16108 22324 16148 22364
rect 16012 22072 16052 22112
rect 15628 21148 15668 21188
rect 15340 20476 15380 20516
rect 15628 20476 15668 20516
rect 14860 19468 14900 19508
rect 14764 19300 14804 19340
rect 14668 18880 14708 18920
rect 14668 18712 14708 18752
rect 14572 18376 14612 18416
rect 14476 18292 14516 18332
rect 14380 18208 14420 18248
rect 14284 14848 14324 14888
rect 15340 19384 15380 19424
rect 14956 18712 14996 18752
rect 15052 18628 15092 18668
rect 14668 17200 14708 17240
rect 14764 17116 14804 17156
rect 14476 14512 14516 14552
rect 14380 13168 14420 13208
rect 14284 12664 14324 12704
rect 14284 12412 14324 12452
rect 14284 11656 14324 11696
rect 14764 16696 14804 16736
rect 14668 16360 14708 16400
rect 14668 16024 14708 16064
rect 14668 13672 14708 13712
rect 14668 13084 14708 13124
rect 14572 11572 14612 11612
rect 13804 11236 13844 11276
rect 13996 11152 14036 11192
rect 13900 11068 13940 11108
rect 13900 10816 13940 10856
rect 13804 9724 13844 9764
rect 13420 8128 13460 8168
rect 13420 7960 13460 8000
rect 13708 9472 13748 9512
rect 13612 9388 13652 9428
rect 13612 8548 13652 8588
rect 14092 11068 14132 11108
rect 13996 8548 14036 8588
rect 13900 8128 13940 8168
rect 13612 7960 13652 8000
rect 13708 7288 13748 7328
rect 13516 7120 13556 7160
rect 13228 7036 13268 7076
rect 13324 6952 13364 6992
rect 13036 3844 13076 3884
rect 12940 3088 12980 3128
rect 14380 9976 14420 10016
rect 14284 9472 14324 9512
rect 15052 18376 15092 18416
rect 15244 17704 15284 17744
rect 15436 18124 15476 18164
rect 15628 17956 15668 17996
rect 16012 21400 16052 21440
rect 15916 19636 15956 19676
rect 15820 19216 15860 19256
rect 15148 17032 15188 17072
rect 15052 16948 15092 16988
rect 15052 16360 15092 16400
rect 15532 16696 15572 16736
rect 15340 16528 15380 16568
rect 14956 16024 14996 16064
rect 14956 15520 14996 15560
rect 15436 16360 15476 16400
rect 15628 16192 15668 16232
rect 15148 14512 15188 14552
rect 15532 14092 15572 14132
rect 15436 14008 15476 14048
rect 15244 13168 15284 13208
rect 15916 18544 15956 18584
rect 16012 18292 16052 18332
rect 15916 17956 15956 17996
rect 15820 17032 15860 17072
rect 15820 16696 15860 16736
rect 15820 15520 15860 15560
rect 16012 17872 16052 17912
rect 15916 14596 15956 14636
rect 16204 20560 16244 20600
rect 16204 20308 16244 20348
rect 16204 19216 16244 19256
rect 16204 18628 16244 18668
rect 16108 15436 16148 15476
rect 16012 14344 16052 14384
rect 15916 14260 15956 14300
rect 16492 24592 16532 24632
rect 16588 24172 16628 24212
rect 16588 23920 16628 23960
rect 16396 23836 16436 23876
rect 16396 23248 16436 23288
rect 16492 22996 16532 23036
rect 17068 27532 17108 27572
rect 16876 26776 16916 26816
rect 16876 26608 16916 26648
rect 16972 26440 17012 26480
rect 16876 26020 16916 26060
rect 16876 25684 16916 25724
rect 16780 25012 16820 25052
rect 16396 22660 16436 22700
rect 16492 21652 16532 21692
rect 16396 21568 16436 21608
rect 16396 17200 16436 17240
rect 16684 22324 16724 22364
rect 16876 23248 16916 23288
rect 17068 26272 17108 26312
rect 17068 26104 17108 26144
rect 18028 32824 18068 32864
rect 17740 31396 17780 31436
rect 17836 31228 17876 31268
rect 17836 30640 17876 30680
rect 17932 30472 17972 30512
rect 17836 30388 17876 30428
rect 17740 30220 17780 30260
rect 17548 30052 17588 30092
rect 17356 29632 17396 29672
rect 17548 29380 17588 29420
rect 17740 29800 17780 29840
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 18700 37696 18740 37736
rect 19276 37444 19316 37484
rect 19468 39460 19508 39500
rect 19468 38704 19508 38744
rect 19468 38368 19508 38408
rect 19660 39628 19700 39668
rect 19660 38956 19700 38996
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 20044 39880 20084 39920
rect 19852 39712 19892 39752
rect 19852 39040 19892 39080
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 20044 38116 20084 38156
rect 20236 38032 20276 38072
rect 19852 37948 19892 37988
rect 20044 37444 20084 37484
rect 19660 37276 19700 37316
rect 19372 37108 19412 37148
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 19468 36268 19508 36308
rect 19756 36940 19796 36980
rect 18988 36100 19028 36140
rect 20236 37360 20276 37400
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 20140 36688 20180 36728
rect 19948 36184 19988 36224
rect 18316 35260 18356 35300
rect 18220 33748 18260 33788
rect 18220 33412 18260 33452
rect 19180 35344 19220 35384
rect 18988 35092 19028 35132
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 20044 36016 20084 36056
rect 19564 35932 19604 35972
rect 19852 35764 19892 35804
rect 19468 34672 19508 34712
rect 19372 34504 19412 34544
rect 19756 35680 19796 35720
rect 19660 35008 19700 35048
rect 19852 35596 19892 35636
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 20524 35344 20564 35384
rect 18412 33664 18452 33704
rect 18412 32740 18452 32780
rect 18316 32656 18356 32696
rect 18124 31228 18164 31268
rect 18124 30388 18164 30428
rect 18316 30052 18356 30092
rect 18124 29464 18164 29504
rect 18028 29296 18068 29336
rect 17932 29128 17972 29168
rect 17836 29044 17876 29084
rect 17356 28624 17396 28664
rect 17260 28372 17300 28412
rect 17356 28120 17396 28160
rect 17548 28288 17588 28328
rect 17260 27112 17300 27152
rect 17452 27112 17492 27152
rect 17356 26860 17396 26900
rect 17260 26272 17300 26312
rect 17260 25936 17300 25976
rect 17260 25432 17300 25472
rect 17932 28876 17972 28916
rect 17740 26524 17780 26564
rect 17740 25600 17780 25640
rect 17644 25432 17684 25472
rect 17452 25348 17492 25388
rect 17253 25264 17260 25304
rect 17260 25264 17293 25304
rect 17356 25264 17396 25304
rect 17356 24424 17396 24464
rect 17164 23584 17204 23624
rect 17356 23920 17396 23960
rect 17548 25180 17588 25220
rect 17548 23920 17588 23960
rect 17452 23164 17492 23204
rect 16876 22996 16916 23036
rect 17260 22912 17300 22952
rect 16972 21904 17012 21944
rect 17068 21652 17108 21692
rect 16684 20812 16724 20852
rect 16876 21568 16916 21608
rect 17164 21568 17204 21608
rect 17260 21484 17300 21524
rect 16972 21316 17012 21356
rect 17164 21232 17204 21272
rect 16876 20560 16916 20600
rect 16684 18628 16724 18668
rect 16780 18208 16820 18248
rect 16588 17788 16628 17828
rect 16396 16948 16436 16988
rect 16972 19972 17012 20012
rect 17068 19720 17108 19760
rect 17068 19132 17108 19172
rect 17260 20812 17300 20852
rect 17644 23080 17684 23120
rect 17644 21568 17684 21608
rect 17452 20980 17492 21020
rect 17356 20560 17396 20600
rect 17548 20560 17588 20600
rect 17452 20056 17492 20096
rect 17260 19888 17300 19928
rect 17260 19636 17300 19676
rect 17932 25768 17972 25808
rect 18220 29380 18260 29420
rect 18604 33832 18644 33872
rect 19276 33916 19316 33956
rect 19660 34252 19700 34292
rect 19564 33916 19604 33956
rect 19468 33580 19508 33620
rect 18700 33328 18740 33368
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 19180 33076 19220 33116
rect 18604 32908 18644 32948
rect 18796 32824 18836 32864
rect 18604 32152 18644 32192
rect 18988 32488 19028 32528
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 19084 31564 19124 31604
rect 20044 34168 20084 34208
rect 19852 34084 19892 34124
rect 19372 32824 19412 32864
rect 19372 31480 19412 31520
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 19948 33832 19988 33872
rect 20044 33748 20084 33788
rect 19852 33076 19892 33116
rect 19756 32992 19796 33032
rect 19948 32992 19988 33032
rect 19852 32740 19892 32780
rect 19660 32572 19700 32612
rect 19564 31144 19604 31184
rect 19372 30556 19412 30596
rect 18988 30388 19028 30428
rect 18508 29464 18548 29504
rect 18412 29296 18452 29336
rect 18508 29128 18548 29168
rect 18316 28876 18356 28916
rect 18316 28624 18356 28664
rect 18220 27532 18260 27572
rect 19468 30388 19508 30428
rect 18700 30220 18740 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 19372 29800 19412 29840
rect 19276 29296 19316 29336
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18700 28624 18740 28664
rect 18604 28540 18644 28580
rect 18988 28540 19028 28580
rect 18700 27616 18740 27656
rect 19084 28036 19124 28076
rect 19084 27532 19124 27572
rect 18412 27196 18452 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 18124 26608 18164 26648
rect 18124 26104 18164 26144
rect 18028 25600 18068 25640
rect 18028 25432 18068 25472
rect 17932 25348 17972 25388
rect 17932 24508 17972 24548
rect 17932 24340 17972 24380
rect 18124 25180 18164 25220
rect 18412 26356 18452 26396
rect 19756 30892 19796 30932
rect 20428 32656 20468 32696
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 21004 32656 21044 32696
rect 20044 32236 20084 32276
rect 20524 31648 20564 31688
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 20620 30640 20660 30680
rect 19756 30136 19796 30176
rect 19660 29716 19700 29756
rect 19852 30052 19892 30092
rect 19852 29800 19892 29840
rect 20044 29884 20084 29924
rect 19948 29632 19988 29672
rect 19852 29296 19892 29336
rect 19756 29128 19796 29168
rect 19660 29044 19700 29084
rect 19564 28960 19604 29000
rect 19660 28876 19700 28916
rect 19564 28792 19604 28832
rect 19756 28540 19796 28580
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 20716 29968 20756 30008
rect 20044 29128 20084 29168
rect 19852 28456 19892 28496
rect 19660 28288 19700 28328
rect 19660 27868 19700 27908
rect 19948 28372 19988 28412
rect 19756 27364 19796 27404
rect 19372 26860 19412 26900
rect 18700 26272 18740 26312
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 20044 27784 20084 27824
rect 20716 27700 20756 27740
rect 20524 26944 20564 26984
rect 19468 26692 19508 26732
rect 18988 26440 19028 26480
rect 18892 26272 18932 26312
rect 18892 26104 18932 26144
rect 19276 26356 19316 26396
rect 19180 25852 19220 25892
rect 19564 26608 19604 26648
rect 19948 26608 19988 26648
rect 20812 26608 20852 26648
rect 20524 26524 20564 26564
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 18316 25516 18356 25556
rect 18220 24760 18260 24800
rect 18124 23080 18164 23120
rect 18412 25180 18452 25220
rect 18220 22912 18260 22952
rect 17932 22408 17972 22448
rect 18023 20728 18063 20768
rect 17932 19552 17972 19592
rect 17836 19384 17876 19424
rect 17548 19216 17588 19256
rect 16972 18460 17012 18500
rect 16972 17452 17012 17492
rect 16300 14092 16340 14132
rect 15724 13840 15764 13880
rect 15532 13084 15572 13124
rect 15148 12664 15188 12704
rect 14956 12496 14996 12536
rect 15148 12328 15188 12368
rect 14860 11908 14900 11948
rect 15148 11824 15188 11864
rect 15148 11656 15188 11696
rect 14668 10900 14708 10940
rect 15052 11068 15092 11108
rect 14956 9808 14996 9848
rect 14860 9724 14900 9764
rect 14668 9640 14708 9680
rect 14572 9304 14612 9344
rect 14668 8800 14708 8840
rect 14476 8128 14516 8168
rect 14860 8128 14900 8168
rect 14092 6868 14132 6908
rect 13420 6532 13460 6572
rect 13996 6448 14036 6488
rect 13996 6280 14036 6320
rect 13804 2668 13844 2708
rect 14380 6952 14420 6992
rect 14668 6196 14708 6236
rect 14860 7120 14900 7160
rect 15340 11572 15380 11612
rect 15916 13840 15956 13880
rect 16012 13756 16052 13796
rect 16300 13756 16340 13796
rect 15820 13168 15860 13208
rect 15724 13000 15764 13040
rect 16204 13168 16244 13208
rect 16108 13084 16148 13124
rect 15820 12664 15860 12704
rect 15628 12244 15668 12284
rect 15532 11488 15572 11528
rect 15724 11656 15764 11696
rect 15724 10984 15764 11024
rect 15724 10144 15764 10184
rect 15244 9976 15284 10016
rect 15340 8800 15380 8840
rect 15436 8632 15476 8672
rect 15532 8464 15572 8504
rect 15052 7540 15092 7580
rect 14956 6616 14996 6656
rect 15436 7120 15476 7160
rect 15532 7036 15572 7076
rect 16012 12412 16052 12452
rect 16012 12244 16052 12284
rect 15916 11152 15956 11192
rect 15916 10984 15956 11024
rect 16396 13252 16436 13292
rect 16588 16192 16628 16232
rect 16684 15856 16724 15896
rect 16588 15520 16628 15560
rect 16588 14260 16628 14300
rect 16492 13168 16532 13208
rect 16300 12664 16340 12704
rect 16588 12580 16628 12620
rect 16396 12412 16436 12452
rect 16012 10900 16052 10940
rect 16108 10228 16148 10268
rect 16012 8632 16052 8672
rect 15916 7204 15956 7244
rect 15532 6700 15572 6740
rect 14764 5020 14804 5060
rect 15532 5020 15572 5060
rect 15148 3592 15188 3632
rect 14380 2668 14420 2708
rect 13900 2080 13940 2120
rect 12748 1660 12788 1700
rect 12652 736 12692 776
rect 13900 1492 13940 1532
rect 13132 1408 13172 1448
rect 13708 1240 13748 1280
rect 13036 1156 13076 1196
rect 13420 1156 13460 1196
rect 12940 820 12980 860
rect 12940 484 12980 524
rect 13324 400 13364 440
rect 13132 316 13172 356
rect 13612 904 13652 944
rect 13804 1156 13844 1196
rect 14284 2416 14324 2456
rect 14572 2416 14612 2456
rect 15148 2416 15188 2456
rect 14572 2080 14612 2120
rect 14284 1828 14324 1868
rect 14476 1660 14516 1700
rect 14476 1324 14516 1364
rect 14092 988 14132 1028
rect 14284 904 14324 944
rect 14380 316 14420 356
rect 14668 1828 14708 1868
rect 15244 2080 15284 2120
rect 14860 1660 14900 1700
rect 14668 904 14708 944
rect 14764 484 14804 524
rect 14956 1156 14996 1196
rect 15052 820 15092 860
rect 15148 400 15188 440
rect 15436 1744 15476 1784
rect 15436 1408 15476 1448
rect 15628 1828 15668 1868
rect 15532 1324 15572 1364
rect 15628 1240 15668 1280
rect 15532 652 15572 692
rect 15820 6700 15860 6740
rect 15916 4096 15956 4136
rect 15916 3172 15956 3212
rect 15820 1828 15860 1868
rect 15820 1492 15860 1532
rect 15820 1324 15860 1364
rect 16012 1828 16052 1868
rect 16300 10900 16340 10940
rect 16204 10144 16244 10184
rect 16588 12328 16628 12368
rect 16492 12244 16532 12284
rect 16396 9556 16436 9596
rect 16588 11404 16628 11444
rect 16588 11236 16628 11276
rect 17164 18376 17204 18416
rect 17260 18124 17300 18164
rect 17164 17956 17204 17996
rect 17260 17872 17300 17912
rect 17452 17872 17492 17912
rect 17164 17284 17204 17324
rect 17356 17788 17396 17828
rect 17260 16276 17300 16316
rect 16876 16192 16916 16232
rect 16972 15856 17012 15896
rect 16780 15520 16820 15560
rect 16780 14848 16820 14888
rect 16780 14680 16820 14720
rect 16972 15688 17012 15728
rect 17260 15100 17300 15140
rect 17644 19048 17684 19088
rect 17548 17284 17588 17324
rect 17644 17032 17684 17072
rect 17644 16276 17684 16316
rect 17644 15772 17684 15812
rect 17548 15688 17588 15728
rect 17452 15520 17492 15560
rect 17452 15268 17492 15308
rect 17356 14848 17396 14888
rect 17068 14512 17108 14552
rect 17836 19048 17876 19088
rect 17836 17536 17876 17576
rect 18220 19972 18260 20012
rect 18124 19720 18164 19760
rect 18124 19468 18164 19508
rect 18028 17620 18068 17660
rect 18220 18040 18260 18080
rect 18124 16696 18164 16736
rect 18220 16612 18260 16652
rect 17932 15856 17972 15896
rect 17740 15352 17780 15392
rect 17644 15268 17684 15308
rect 17740 15184 17780 15224
rect 17932 15100 17972 15140
rect 17836 15016 17876 15056
rect 17164 14344 17204 14384
rect 16780 12412 16820 12452
rect 16972 12664 17012 12704
rect 17068 12412 17108 12452
rect 16780 11992 16820 12032
rect 16972 11656 17012 11696
rect 17548 14512 17588 14552
rect 17548 14344 17588 14384
rect 17452 14260 17492 14300
rect 17356 14043 17396 14048
rect 17356 14008 17396 14043
rect 17260 13168 17300 13208
rect 17836 14260 17876 14300
rect 18220 15688 18260 15728
rect 18124 15520 18164 15560
rect 18604 24844 18644 24884
rect 18604 23920 18644 23960
rect 18508 23080 18548 23120
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 19084 25516 19124 25556
rect 19180 25432 19220 25472
rect 18892 25180 18932 25220
rect 19564 25852 19604 25892
rect 19756 26104 19796 26144
rect 19468 25432 19508 25472
rect 19660 25432 19700 25472
rect 19852 25432 19892 25472
rect 19468 25096 19508 25136
rect 19756 25348 19796 25388
rect 19276 24844 19316 24884
rect 19372 24760 19412 24800
rect 19660 24760 19700 24800
rect 18988 24592 19028 24632
rect 19084 24508 19124 24548
rect 18988 24340 19028 24380
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 19276 23752 19316 23792
rect 19121 23248 19161 23288
rect 19564 24256 19604 24296
rect 19660 23920 19700 23960
rect 19564 23752 19604 23792
rect 19852 24844 19892 24884
rect 20044 25096 20084 25136
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20524 24928 20564 24968
rect 20044 24760 20084 24800
rect 20044 24424 20084 24464
rect 20524 24424 20564 24464
rect 18412 22660 18452 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 18700 21652 18740 21692
rect 18604 20560 18644 20600
rect 19180 21568 19220 21608
rect 19852 23248 19892 23288
rect 19660 22828 19700 22868
rect 19564 21736 19604 21776
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 18796 20392 18836 20432
rect 18508 20140 18548 20180
rect 19564 21568 19604 21608
rect 19852 23080 19892 23120
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 20140 23248 20180 23288
rect 19852 22408 19892 22448
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 20812 24256 20852 24296
rect 21388 29296 21428 29336
rect 21388 22912 21428 22952
rect 20812 22576 20852 22616
rect 20620 21904 20660 21944
rect 19852 21652 19892 21692
rect 19948 21568 19988 21608
rect 19468 20896 19508 20936
rect 20140 21568 20180 21608
rect 19180 20728 19220 20768
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 19948 20308 19988 20348
rect 18412 19888 18452 19928
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 18604 19132 18644 19172
rect 19276 19132 19316 19172
rect 18412 17368 18452 17408
rect 18028 14344 18068 14384
rect 17740 14008 17780 14048
rect 17836 13840 17876 13880
rect 18220 15184 18260 15224
rect 17164 12244 17204 12284
rect 17548 12664 17588 12704
rect 17068 11572 17108 11612
rect 17260 11656 17300 11696
rect 17356 11572 17396 11612
rect 17644 12412 17684 12452
rect 16972 11152 17012 11192
rect 16876 10984 16916 11024
rect 17740 11320 17780 11360
rect 16684 9808 16724 9848
rect 17068 10816 17108 10856
rect 16972 10228 17012 10268
rect 16972 9976 17012 10016
rect 16588 9472 16628 9512
rect 16492 7288 16532 7328
rect 17164 10648 17204 10688
rect 17260 10480 17300 10520
rect 17644 10984 17684 11024
rect 17548 10816 17588 10856
rect 17452 10480 17492 10520
rect 17164 8800 17204 8840
rect 17740 10816 17780 10856
rect 17740 10480 17780 10520
rect 21196 21232 21236 21272
rect 21100 20896 21140 20936
rect 21100 20140 21140 20180
rect 19660 19804 19700 19844
rect 19852 19888 19892 19928
rect 20044 20056 20084 20096
rect 19948 19720 19988 19760
rect 19948 19300 19988 19340
rect 19660 19132 19700 19172
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 20044 18712 20084 18752
rect 20236 18712 20276 18752
rect 19084 18628 19124 18668
rect 19756 18628 19796 18668
rect 19180 18376 19220 18416
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 18796 17956 18836 17996
rect 19468 17956 19508 17996
rect 18892 17704 18932 17744
rect 19276 17704 19316 17744
rect 19852 18376 19892 18416
rect 19180 17452 19220 17492
rect 19276 17116 19316 17156
rect 18700 16948 18740 16988
rect 18604 16780 18644 16820
rect 18604 16612 18644 16652
rect 18892 16780 18932 16820
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 18796 16192 18836 16232
rect 18700 16108 18740 16148
rect 18700 15940 18740 15980
rect 19468 16360 19508 16400
rect 19180 16276 19220 16316
rect 19084 16192 19124 16232
rect 18988 15940 19028 15980
rect 19948 18040 19988 18080
rect 20044 17704 20084 17744
rect 19948 17620 19988 17660
rect 19660 17452 19700 17492
rect 19852 17284 19892 17324
rect 19660 16948 19700 16988
rect 19372 16192 19412 16232
rect 19756 16192 19796 16232
rect 19276 16024 19316 16064
rect 19276 15856 19316 15896
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 19468 15856 19508 15896
rect 19852 15772 19892 15812
rect 19660 15436 19700 15476
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 20044 16444 20084 16484
rect 20044 16024 20084 16064
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 20908 19888 20948 19928
rect 20812 19552 20852 19592
rect 19564 15268 19604 15308
rect 20044 15268 20084 15308
rect 18700 14596 18740 14636
rect 18604 14428 18644 14468
rect 17932 12496 17972 12536
rect 17932 11908 17972 11948
rect 18028 11236 18068 11276
rect 17932 11152 17972 11192
rect 17836 10312 17876 10352
rect 18028 10648 18068 10688
rect 18604 12580 18644 12620
rect 18508 12496 18548 12536
rect 18220 11488 18260 11528
rect 19372 14680 19412 14720
rect 19660 14680 19700 14720
rect 18988 13756 19028 13796
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 19276 13504 19316 13544
rect 19084 13336 19124 13376
rect 19276 13252 19316 13292
rect 18796 12496 18836 12536
rect 19660 14428 19700 14468
rect 19468 12748 19508 12788
rect 19852 14764 19892 14804
rect 19948 14680 19988 14720
rect 19564 12664 19604 12704
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 18220 11236 18260 11276
rect 18508 10984 18548 11024
rect 18220 10816 18260 10856
rect 18124 10480 18164 10520
rect 17356 9808 17396 9848
rect 17644 9472 17684 9512
rect 17644 8632 17684 8672
rect 17260 8128 17300 8168
rect 17644 8464 17684 8504
rect 17164 7036 17204 7076
rect 16684 6532 16724 6572
rect 16492 6448 16532 6488
rect 16396 6196 16436 6236
rect 16396 1828 16436 1868
rect 16204 1660 16244 1700
rect 15916 904 15956 944
rect 16108 1156 16148 1196
rect 16588 1408 16628 1448
rect 16876 6364 16916 6404
rect 16780 1828 16820 1868
rect 16972 6280 17012 6320
rect 17164 6196 17204 6236
rect 17356 3592 17396 3632
rect 17260 2080 17300 2120
rect 17644 2080 17684 2120
rect 17548 1828 17588 1868
rect 17932 10144 17972 10184
rect 18028 9976 18068 10016
rect 17932 9808 17972 9848
rect 17836 8800 17876 8840
rect 18028 9724 18068 9764
rect 18316 10480 18356 10520
rect 18604 10396 18644 10436
rect 19372 12076 19412 12116
rect 19372 11824 19412 11864
rect 18892 11236 18932 11276
rect 18892 10816 18932 10856
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18892 10228 18932 10268
rect 18604 9976 18644 10016
rect 18124 9640 18164 9680
rect 18508 9304 18548 9344
rect 18028 6532 18068 6572
rect 17932 6448 17972 6488
rect 19276 9724 19316 9764
rect 19564 12496 19604 12536
rect 19564 12328 19604 12368
rect 19468 9808 19508 9848
rect 19084 9640 19124 9680
rect 19372 9640 19412 9680
rect 19367 9472 19407 9512
rect 19564 9472 19604 9512
rect 19084 9220 19124 9260
rect 19852 12664 19892 12704
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 21100 16276 21140 16316
rect 21004 16192 21044 16232
rect 20812 14848 20852 14888
rect 20044 13924 20084 13964
rect 20716 13672 20756 13712
rect 20044 13252 20084 13292
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 20236 12580 20276 12620
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 19948 10228 19988 10268
rect 20140 10144 20180 10184
rect 20812 12496 20852 12536
rect 20716 10144 20756 10184
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 19660 9388 19700 9428
rect 19468 9220 19508 9260
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 19372 8968 19412 9008
rect 19084 8884 19124 8924
rect 18892 7960 18932 8000
rect 19180 7876 19220 7916
rect 19084 7708 19124 7748
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18988 7372 19028 7412
rect 18796 7288 18836 7328
rect 18700 7120 18740 7160
rect 20044 9472 20084 9512
rect 20140 9388 20180 9428
rect 19852 8968 19892 9008
rect 19756 8884 19796 8924
rect 20236 9304 20276 9344
rect 20524 9136 20564 9176
rect 19564 8632 19604 8672
rect 19564 7960 19604 8000
rect 19372 7288 19412 7328
rect 18604 6952 18644 6992
rect 20236 8884 20276 8924
rect 19756 8128 19796 8168
rect 19756 7792 19796 7832
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19948 8128 19988 8168
rect 20140 8128 20180 8168
rect 20716 8128 20756 8168
rect 19948 7960 19988 8000
rect 21292 20560 21332 20600
rect 21388 20056 21428 20096
rect 21292 15940 21332 15980
rect 21196 15772 21236 15812
rect 21388 15352 21428 15392
rect 21196 13420 21236 13460
rect 21196 10480 21236 10520
rect 21100 9724 21140 9764
rect 21196 8884 21236 8924
rect 21100 8128 21140 8168
rect 20044 7876 20084 7916
rect 19564 6952 19604 6992
rect 18700 6700 18740 6740
rect 19564 6700 19604 6740
rect 18604 6364 18644 6404
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 19756 6784 19796 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 19948 6364 19988 6404
rect 19468 5440 19508 5480
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 19948 5020 19988 5060
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 18028 2080 18068 2120
rect 18412 2080 18452 2120
rect 17836 1828 17876 1868
rect 18028 1240 18068 1280
rect 17644 148 17684 188
rect 17932 316 17972 356
rect 18508 1660 18548 1700
rect 18508 1324 18548 1364
rect 18412 1240 18452 1280
rect 18796 2248 18836 2288
rect 19180 2080 19220 2120
rect 19564 2080 19604 2120
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 18988 1660 19028 1700
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 19372 1492 19412 1532
rect 21292 1744 21332 1784
rect 18412 988 18452 1028
rect 18316 316 18356 356
rect 18700 1072 18740 1112
rect 19180 904 19220 944
rect 21388 1408 21428 1448
rect 20524 1324 20564 1364
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 20524 400 20564 440
<< metal3 >>
rect 19075 85952 19133 85953
rect 18990 85912 19084 85952
rect 19124 85912 19133 85952
rect 19075 85911 19133 85912
rect 19267 85952 19325 85953
rect 19267 85912 19276 85952
rect 19316 85912 19410 85952
rect 19267 85911 19325 85912
rect 7171 85828 7180 85868
rect 7220 85828 15724 85868
rect 15764 85828 15773 85868
rect 21424 85784 21504 85804
rect 19267 85744 19276 85784
rect 19316 85744 21504 85784
rect 21424 85724 21504 85744
rect 6499 85616 6557 85617
rect 16003 85616 16061 85617
rect 6403 85576 6412 85616
rect 6452 85576 6508 85616
rect 6548 85576 6557 85616
rect 15427 85576 15436 85616
rect 15476 85576 16012 85616
rect 16052 85576 16061 85616
rect 6499 85575 6557 85576
rect 16003 85575 16061 85576
rect 16867 85616 16925 85617
rect 16867 85576 16876 85616
rect 16916 85576 16972 85616
rect 17012 85576 17021 85616
rect 16867 85575 16925 85576
rect 21424 85448 21504 85468
rect 8515 85408 8524 85448
rect 8564 85408 18028 85448
rect 18068 85408 18077 85448
rect 19555 85408 19564 85448
rect 19604 85408 21504 85448
rect 21424 85388 21504 85408
rect 2371 85196 2429 85197
rect 2371 85156 2380 85196
rect 2420 85156 5644 85196
rect 5684 85156 5693 85196
rect 2371 85155 2429 85156
rect 17923 85112 17981 85113
rect 1027 85072 1036 85112
rect 1076 85072 6028 85112
rect 6068 85072 6077 85112
rect 17838 85072 17932 85112
rect 17972 85072 17981 85112
rect 17923 85071 17981 85072
rect 19843 85112 19901 85113
rect 21424 85112 21504 85132
rect 19843 85072 19852 85112
rect 19892 85072 21504 85112
rect 19843 85071 19901 85072
rect 21424 85052 21504 85072
rect 4099 84988 4108 85028
rect 4148 84988 4396 85028
rect 4436 84988 4445 85028
rect 16387 84944 16445 84945
rect 20611 84944 20669 84945
rect 14467 84904 14476 84944
rect 14516 84904 16396 84944
rect 16436 84904 16445 84944
rect 18883 84904 18892 84944
rect 18932 84904 20620 84944
rect 20660 84904 20669 84944
rect 16387 84903 16445 84904
rect 20611 84903 20669 84904
rect 3427 84820 3436 84860
rect 3476 84820 3724 84860
rect 3764 84820 3773 84860
rect 7747 84820 7756 84860
rect 7796 84820 13228 84860
rect 13268 84820 13277 84860
rect 21424 84776 21504 84796
rect 19843 84736 19852 84776
rect 19892 84736 21504 84776
rect 21424 84716 21504 84736
rect 3679 84652 3688 84692
rect 3728 84652 3770 84692
rect 3810 84652 3852 84692
rect 3892 84652 3934 84692
rect 3974 84652 4016 84692
rect 4056 84652 4065 84692
rect 5059 84652 5068 84692
rect 5108 84652 8524 84692
rect 8564 84652 8573 84692
rect 18799 84652 18808 84692
rect 18848 84652 18890 84692
rect 18930 84652 18972 84692
rect 19012 84652 19054 84692
rect 19094 84652 19136 84692
rect 19176 84652 19185 84692
rect 13891 84608 13949 84609
rect 20707 84608 20765 84609
rect 5251 84568 5260 84608
rect 5300 84568 7796 84608
rect 6883 84524 6941 84525
rect 7756 84524 7796 84568
rect 13891 84568 13900 84608
rect 13940 84568 14668 84608
rect 14708 84568 14717 84608
rect 17731 84568 17740 84608
rect 17780 84568 20716 84608
rect 20756 84568 20765 84608
rect 13891 84567 13949 84568
rect 20707 84567 20765 84568
rect 14275 84524 14333 84525
rect 14947 84524 15005 84525
rect 6595 84484 6604 84524
rect 6644 84484 6892 84524
rect 6932 84484 6941 84524
rect 7747 84484 7756 84524
rect 7796 84484 7805 84524
rect 14083 84484 14092 84524
rect 14132 84484 14284 84524
rect 14324 84484 14333 84524
rect 14851 84484 14860 84524
rect 14900 84484 14956 84524
rect 14996 84484 15005 84524
rect 6883 84483 6941 84484
rect 14275 84483 14333 84484
rect 14947 84483 15005 84484
rect 16771 84524 16829 84525
rect 17731 84524 17789 84525
rect 18595 84524 18653 84525
rect 16771 84484 16780 84524
rect 16820 84484 17356 84524
rect 17396 84484 17405 84524
rect 17731 84484 17740 84524
rect 17780 84484 18316 84524
rect 18356 84484 18365 84524
rect 18595 84484 18604 84524
rect 18644 84484 18700 84524
rect 18740 84484 18749 84524
rect 16771 84483 16829 84484
rect 17731 84483 17789 84484
rect 18595 84483 18653 84484
rect 5827 84440 5885 84441
rect 6211 84440 6269 84441
rect 6787 84440 6845 84441
rect 10627 84440 10685 84441
rect 12163 84440 12221 84441
rect 13315 84440 13373 84441
rect 13699 84440 13757 84441
rect 13987 84440 14045 84441
rect 14659 84440 14717 84441
rect 15043 84440 15101 84441
rect 15523 84440 15581 84441
rect 17251 84440 17309 84441
rect 17539 84440 17597 84441
rect 3427 84400 3436 84440
rect 3476 84400 4300 84440
rect 4340 84400 4349 84440
rect 5742 84400 5836 84440
rect 5876 84400 5885 84440
rect 6126 84400 6220 84440
rect 6260 84400 6269 84440
rect 6702 84400 6796 84440
rect 6836 84400 6845 84440
rect 8419 84400 8428 84440
rect 8468 84400 10060 84440
rect 10100 84400 10109 84440
rect 10542 84400 10636 84440
rect 10676 84400 10685 84440
rect 12078 84400 12172 84440
rect 12212 84400 12221 84440
rect 13230 84400 13324 84440
rect 13364 84400 13373 84440
rect 13614 84400 13708 84440
rect 13748 84400 13757 84440
rect 13891 84400 13900 84440
rect 13940 84400 13996 84440
rect 14036 84400 14045 84440
rect 14275 84400 14284 84440
rect 14324 84400 14668 84440
rect 14708 84400 14717 84440
rect 14958 84400 15052 84440
rect 15092 84400 15101 84440
rect 15235 84400 15244 84440
rect 15284 84400 15532 84440
rect 15572 84400 15581 84440
rect 17155 84400 17164 84440
rect 17204 84400 17260 84440
rect 17300 84400 17309 84440
rect 17454 84400 17548 84440
rect 17588 84400 17597 84440
rect 5827 84399 5885 84400
rect 6211 84399 6269 84400
rect 6787 84399 6845 84400
rect 10627 84399 10685 84400
rect 12163 84399 12221 84400
rect 13315 84399 13373 84400
rect 13699 84399 13757 84400
rect 13987 84399 14045 84400
rect 14659 84399 14717 84400
rect 15043 84399 15101 84400
rect 15523 84399 15581 84400
rect 17251 84399 17309 84400
rect 17539 84399 17597 84400
rect 17827 84440 17885 84441
rect 18403 84440 18461 84441
rect 19651 84440 19709 84441
rect 21424 84440 21504 84460
rect 17827 84400 17836 84440
rect 17876 84400 18124 84440
rect 18164 84400 18173 84440
rect 18403 84400 18412 84440
rect 18452 84400 18508 84440
rect 18548 84400 18557 84440
rect 19459 84400 19468 84440
rect 19508 84400 19660 84440
rect 19700 84400 19709 84440
rect 20515 84400 20524 84440
rect 20564 84400 21504 84440
rect 17827 84399 17885 84400
rect 18403 84399 18461 84400
rect 19651 84399 19709 84400
rect 21424 84380 21504 84400
rect 8899 84356 8957 84357
rect 4483 84316 4492 84356
rect 4532 84316 8908 84356
rect 8948 84316 8957 84356
rect 8899 84315 8957 84316
rect 21424 84104 21504 84124
rect 4867 84064 4876 84104
rect 4916 84064 5356 84104
rect 5396 84064 5405 84104
rect 20611 84064 20620 84104
rect 20660 84064 21504 84104
rect 21424 84044 21504 84064
rect 7555 83980 7564 84020
rect 7604 83980 8140 84020
rect 8180 83980 8189 84020
rect 4919 83896 4928 83936
rect 4968 83896 5010 83936
rect 5050 83896 5092 83936
rect 5132 83896 5174 83936
rect 5214 83896 5256 83936
rect 5296 83896 5305 83936
rect 7843 83896 7852 83936
rect 7892 83896 8716 83936
rect 8756 83896 8765 83936
rect 9283 83896 9292 83936
rect 9332 83896 9580 83936
rect 9620 83896 9629 83936
rect 20039 83896 20048 83936
rect 20088 83896 20130 83936
rect 20170 83896 20212 83936
rect 20252 83896 20294 83936
rect 20334 83896 20376 83936
rect 20416 83896 20425 83936
rect 3331 83812 3340 83852
rect 3380 83812 4108 83852
rect 4148 83812 4157 83852
rect 6595 83812 6604 83852
rect 6644 83812 11404 83852
rect 11444 83812 11453 83852
rect 21424 83768 21504 83788
rect 6691 83728 6700 83768
rect 6740 83728 7468 83768
rect 7508 83728 7517 83768
rect 7939 83728 7948 83768
rect 7988 83728 14956 83768
rect 14996 83728 15005 83768
rect 19267 83728 19276 83768
rect 19316 83728 21504 83768
rect 21424 83708 21504 83728
rect 5539 83644 5548 83684
rect 5588 83644 10348 83684
rect 10388 83644 10397 83684
rect 10915 83600 10973 83601
rect 2179 83560 2188 83600
rect 2228 83560 2668 83600
rect 2708 83560 2717 83600
rect 4012 83560 10924 83600
rect 10964 83560 10973 83600
rect 1507 83516 1565 83517
rect 2083 83516 2141 83517
rect 1422 83476 1516 83516
rect 1556 83476 1565 83516
rect 1998 83476 2092 83516
rect 2132 83476 2141 83516
rect 1507 83475 1565 83476
rect 2083 83475 2141 83476
rect 2275 83516 2333 83517
rect 4012 83516 4052 83560
rect 10915 83559 10973 83560
rect 7171 83516 7229 83517
rect 7363 83516 7421 83517
rect 8131 83516 8189 83517
rect 13603 83516 13661 83517
rect 15331 83516 15389 83517
rect 16195 83516 16253 83517
rect 2275 83476 2284 83516
rect 2324 83476 2860 83516
rect 2900 83476 2909 83516
rect 4003 83476 4012 83516
rect 4052 83476 4061 83516
rect 6115 83476 6124 83516
rect 6164 83476 6320 83516
rect 6979 83476 6988 83516
rect 7028 83476 7180 83516
rect 7220 83476 7229 83516
rect 7278 83476 7372 83516
rect 7412 83476 7421 83516
rect 8046 83476 8140 83516
rect 8180 83476 8189 83516
rect 8707 83476 8716 83516
rect 8756 83476 9292 83516
rect 9332 83476 9341 83516
rect 13507 83476 13516 83516
rect 13556 83476 13612 83516
rect 13652 83476 13661 83516
rect 15139 83476 15148 83516
rect 15188 83476 15340 83516
rect 15380 83476 15389 83516
rect 15907 83476 15916 83516
rect 15956 83476 16204 83516
rect 16244 83476 16253 83516
rect 2275 83475 2333 83476
rect 6280 83432 6320 83476
rect 7171 83475 7229 83476
rect 7363 83475 7421 83476
rect 8131 83475 8189 83476
rect 13603 83475 13661 83476
rect 15331 83475 15389 83476
rect 16195 83475 16253 83476
rect 21424 83432 21504 83452
rect 6280 83392 10924 83432
rect 10964 83392 10973 83432
rect 19651 83392 19660 83432
rect 19700 83392 21504 83432
rect 21424 83372 21504 83392
rect 2659 83348 2717 83349
rect 2659 83308 2668 83348
rect 2708 83308 3628 83348
rect 3668 83308 3677 83348
rect 4387 83308 4396 83348
rect 4436 83308 8620 83348
rect 8660 83308 8669 83348
rect 18979 83308 18988 83348
rect 19028 83308 19468 83348
rect 19508 83308 19517 83348
rect 2659 83307 2717 83308
rect 5155 83224 5164 83264
rect 5204 83224 8524 83264
rect 8564 83224 8573 83264
rect 9187 83224 9196 83264
rect 9236 83224 11980 83264
rect 12020 83224 12029 83264
rect 6979 83180 7037 83181
rect 8227 83180 8285 83181
rect 3679 83140 3688 83180
rect 3728 83140 3770 83180
rect 3810 83140 3852 83180
rect 3892 83140 3934 83180
rect 3974 83140 4016 83180
rect 4056 83140 4065 83180
rect 4771 83140 4780 83180
rect 4820 83140 5548 83180
rect 5588 83140 5597 83180
rect 6499 83140 6508 83180
rect 6548 83140 6988 83180
rect 7028 83140 7037 83180
rect 7939 83140 7948 83180
rect 7988 83140 8236 83180
rect 8276 83140 8285 83180
rect 9379 83140 9388 83180
rect 9428 83140 10444 83180
rect 10484 83140 10493 83180
rect 18799 83140 18808 83180
rect 18848 83140 18890 83180
rect 18930 83140 18972 83180
rect 19012 83140 19054 83180
rect 19094 83140 19136 83180
rect 19176 83140 19185 83180
rect 6979 83139 7037 83140
rect 8227 83139 8285 83140
rect 21424 83096 21504 83116
rect 15715 83056 15724 83096
rect 15764 83056 21504 83096
rect 21424 83036 21504 83056
rect 2851 82844 2909 82845
rect 3235 82844 3293 82845
rect 2766 82804 2860 82844
rect 2900 82804 2909 82844
rect 3150 82804 3244 82844
rect 3284 82804 3293 82844
rect 2851 82803 2909 82804
rect 3235 82803 3293 82804
rect 3523 82844 3581 82845
rect 3523 82804 3532 82844
rect 3572 82804 3628 82844
rect 3668 82804 3677 82844
rect 4099 82804 4108 82844
rect 4148 82804 4157 82844
rect 4771 82804 4780 82844
rect 4820 82804 7660 82844
rect 7700 82804 7709 82844
rect 13891 82804 13900 82844
rect 13940 82804 18988 82844
rect 19028 82804 19037 82844
rect 3523 82803 3581 82804
rect 4108 82760 4148 82804
rect 19267 82760 19325 82761
rect 21424 82760 21504 82780
rect 4108 82720 19276 82760
rect 19316 82720 19325 82760
rect 21379 82720 21388 82760
rect 21428 82720 21504 82760
rect 19267 82719 19325 82720
rect 21424 82700 21504 82720
rect 21424 82424 21504 82444
rect 4919 82384 4928 82424
rect 4968 82384 5010 82424
rect 5050 82384 5092 82424
rect 5132 82384 5174 82424
rect 5214 82384 5256 82424
rect 5296 82384 5305 82424
rect 20039 82384 20048 82424
rect 20088 82384 20130 82424
rect 20170 82384 20212 82424
rect 20252 82384 20294 82424
rect 20334 82384 20376 82424
rect 20416 82384 20425 82424
rect 20524 82384 21504 82424
rect 20524 82340 20564 82384
rect 21424 82364 21504 82384
rect 10147 82300 10156 82340
rect 10196 82300 11020 82340
rect 11060 82300 11069 82340
rect 19651 82300 19660 82340
rect 19700 82300 20564 82340
rect 14275 82216 14284 82256
rect 14324 82216 21388 82256
rect 21428 82216 21437 82256
rect 21424 82089 21504 82108
rect 21379 82088 21504 82089
rect 21379 82048 21388 82088
rect 21428 82048 21504 82088
rect 21379 82047 21504 82048
rect 21424 82028 21504 82047
rect 6307 81964 6316 82004
rect 6356 81964 12748 82004
rect 12788 81964 12797 82004
rect 15331 81880 15340 81920
rect 15380 81880 15389 81920
rect 15340 81836 15380 81880
rect 11203 81796 11212 81836
rect 11252 81796 15380 81836
rect 21424 81752 21504 81772
rect 19363 81712 19372 81752
rect 19412 81712 19421 81752
rect 19555 81712 19564 81752
rect 19604 81712 21504 81752
rect 3679 81628 3688 81668
rect 3728 81628 3770 81668
rect 3810 81628 3852 81668
rect 3892 81628 3934 81668
rect 3974 81628 4016 81668
rect 4056 81628 4065 81668
rect 18799 81628 18808 81668
rect 18848 81628 18890 81668
rect 18930 81628 18972 81668
rect 19012 81628 19054 81668
rect 19094 81628 19136 81668
rect 19176 81628 19185 81668
rect 19372 81500 19412 81712
rect 21424 81692 21504 81712
rect 19075 81460 19084 81500
rect 19124 81460 19412 81500
rect 21424 81416 21504 81436
rect 19171 81376 19180 81416
rect 19220 81376 19660 81416
rect 19700 81376 19709 81416
rect 19939 81376 19948 81416
rect 19988 81376 21504 81416
rect 21424 81356 21504 81376
rect 13795 81292 13804 81332
rect 13844 81292 19372 81332
rect 19412 81292 19421 81332
rect 5443 81208 5452 81248
rect 5492 81208 12940 81248
rect 12980 81208 12989 81248
rect 2371 81124 2380 81164
rect 2420 81124 18988 81164
rect 19028 81124 19037 81164
rect 21424 81080 21504 81100
rect 18883 81040 18892 81080
rect 18932 81040 21504 81080
rect 21424 81020 21504 81040
rect 4919 80872 4928 80912
rect 4968 80872 5010 80912
rect 5050 80872 5092 80912
rect 5132 80872 5174 80912
rect 5214 80872 5256 80912
rect 5296 80872 5305 80912
rect 20039 80872 20048 80912
rect 20088 80872 20130 80912
rect 20170 80872 20212 80912
rect 20252 80872 20294 80912
rect 20334 80872 20376 80912
rect 20416 80872 20425 80912
rect 21424 80744 21504 80764
rect 19267 80704 19276 80744
rect 19316 80704 21504 80744
rect 21424 80684 21504 80704
rect 13219 80536 13228 80576
rect 13268 80536 19180 80576
rect 19220 80536 19229 80576
rect 19459 80536 19468 80576
rect 19508 80536 20620 80576
rect 20660 80536 20669 80576
rect 8995 80452 9004 80492
rect 9044 80452 19756 80492
rect 19796 80452 19805 80492
rect 21424 80408 21504 80428
rect 16675 80368 16684 80408
rect 16724 80368 21504 80408
rect 21424 80348 21504 80368
rect 16291 80284 16300 80324
rect 16340 80284 19084 80324
rect 19124 80284 19133 80324
rect 13411 80200 13420 80240
rect 13460 80200 19372 80240
rect 19412 80200 19421 80240
rect 3679 80116 3688 80156
rect 3728 80116 3770 80156
rect 3810 80116 3852 80156
rect 3892 80116 3934 80156
rect 3974 80116 4016 80156
rect 4056 80116 4065 80156
rect 18799 80116 18808 80156
rect 18848 80116 18890 80156
rect 18930 80116 18972 80156
rect 19012 80116 19054 80156
rect 19094 80116 19136 80156
rect 19176 80116 19185 80156
rect 21424 80072 21504 80092
rect 19555 80032 19564 80072
rect 19604 80032 21504 80072
rect 21424 80012 21504 80032
rect 11299 79948 11308 79988
rect 11348 79948 19372 79988
rect 19412 79948 19421 79988
rect 11971 79780 11980 79820
rect 12020 79780 12268 79820
rect 12308 79780 14284 79820
rect 14324 79780 15532 79820
rect 15572 79780 15581 79820
rect 15907 79780 15916 79820
rect 15956 79780 18988 79820
rect 19028 79780 19037 79820
rect 21424 79736 21504 79756
rect 11011 79696 11020 79736
rect 11060 79696 12172 79736
rect 12212 79696 14092 79736
rect 14132 79696 14141 79736
rect 19267 79696 19276 79736
rect 19316 79696 19660 79736
rect 19700 79696 19709 79736
rect 19939 79696 19948 79736
rect 19988 79696 21504 79736
rect 21424 79676 21504 79696
rect 9571 79528 9580 79568
rect 9620 79528 13708 79568
rect 13748 79528 13757 79568
rect 15532 79528 19756 79568
rect 19796 79528 19805 79568
rect 15532 79484 15572 79528
rect 3523 79444 3532 79484
rect 3572 79444 15572 79484
rect 16300 79444 16492 79484
rect 16532 79444 16541 79484
rect 19180 79444 20564 79484
rect 4919 79360 4928 79400
rect 4968 79360 5010 79400
rect 5050 79360 5092 79400
rect 5132 79360 5174 79400
rect 5214 79360 5256 79400
rect 5296 79360 5305 79400
rect 10723 79360 10732 79400
rect 10772 79360 11404 79400
rect 11444 79360 11453 79400
rect 12739 79360 12748 79400
rect 12788 79360 13420 79400
rect 13460 79360 13469 79400
rect 14563 79360 14572 79400
rect 14612 79360 16108 79400
rect 16148 79360 16157 79400
rect 11107 79316 11165 79317
rect 16300 79316 16340 79444
rect 19180 79400 19220 79444
rect 20524 79400 20564 79444
rect 21424 79400 21504 79420
rect 16387 79360 16396 79400
rect 16436 79360 16876 79400
rect 16916 79360 16925 79400
rect 19171 79360 19180 79400
rect 19220 79360 19229 79400
rect 20039 79360 20048 79400
rect 20088 79360 20130 79400
rect 20170 79360 20212 79400
rect 20252 79360 20294 79400
rect 20334 79360 20376 79400
rect 20416 79360 20425 79400
rect 20524 79360 21504 79400
rect 21424 79340 21504 79360
rect 10819 79276 10828 79316
rect 10868 79276 11116 79316
rect 11156 79276 11165 79316
rect 13123 79276 13132 79316
rect 13172 79276 14188 79316
rect 14228 79276 14237 79316
rect 15331 79276 15340 79316
rect 15380 79276 16340 79316
rect 11107 79275 11165 79276
rect 9091 79192 9100 79232
rect 9140 79192 9772 79232
rect 9812 79192 9821 79232
rect 9868 79192 19852 79232
rect 19892 79192 19901 79232
rect 9868 79148 9908 79192
rect 6115 79108 6124 79148
rect 6164 79108 9908 79148
rect 10531 79108 10540 79148
rect 10580 79108 10828 79148
rect 10868 79108 10877 79148
rect 11011 79108 11020 79148
rect 11060 79108 11308 79148
rect 11348 79108 11357 79148
rect 11683 79108 11692 79148
rect 11732 79108 19276 79148
rect 19316 79108 19325 79148
rect 11971 79064 12029 79065
rect 21424 79064 21504 79084
rect 10915 79024 10924 79064
rect 10964 79024 11980 79064
rect 12020 79024 12029 79064
rect 16099 79024 16108 79064
rect 16148 79024 16588 79064
rect 16628 79024 16637 79064
rect 18691 79024 18700 79064
rect 18740 79024 21504 79064
rect 11971 79023 12029 79024
rect 21424 79004 21504 79024
rect 11107 78980 11165 78981
rect 11107 78940 11116 78980
rect 11156 78940 11308 78980
rect 11348 78940 11357 78980
rect 11107 78939 11165 78940
rect 9091 78856 9100 78896
rect 9140 78856 15244 78896
rect 15284 78856 15293 78896
rect 20515 78812 20573 78813
rect 5347 78772 5356 78812
rect 5396 78772 18988 78812
rect 19028 78772 19037 78812
rect 19555 78772 19564 78812
rect 19604 78772 20524 78812
rect 20564 78772 20573 78812
rect 20515 78771 20573 78772
rect 21424 78728 21504 78748
rect 19651 78688 19660 78728
rect 19700 78688 21504 78728
rect 21424 78668 21504 78688
rect 3679 78604 3688 78644
rect 3728 78604 3770 78644
rect 3810 78604 3852 78644
rect 3892 78604 3934 78644
rect 3974 78604 4016 78644
rect 4056 78604 4065 78644
rect 18799 78604 18808 78644
rect 18848 78604 18890 78644
rect 18930 78604 18972 78644
rect 19012 78604 19054 78644
rect 19094 78604 19136 78644
rect 19176 78604 19185 78644
rect 0 78560 80 78580
rect 20803 78560 20861 78561
rect 0 78520 172 78560
rect 212 78520 221 78560
rect 19939 78520 19948 78560
rect 19988 78520 20812 78560
rect 20852 78520 20861 78560
rect 0 78500 80 78520
rect 20803 78519 20861 78520
rect 19171 78436 19180 78476
rect 19220 78436 20372 78476
rect 19555 78392 19613 78393
rect 19470 78352 19564 78392
rect 19604 78352 19613 78392
rect 20332 78392 20372 78436
rect 21424 78392 21504 78412
rect 20332 78352 21504 78392
rect 19555 78351 19613 78352
rect 21424 78332 21504 78352
rect 18403 78268 18412 78308
rect 18452 78268 18988 78308
rect 19028 78268 19037 78308
rect 14083 78184 14092 78224
rect 14132 78184 16012 78224
rect 16052 78184 16061 78224
rect 10243 78140 10301 78141
rect 16963 78140 17021 78141
rect 10243 78100 10252 78140
rect 10292 78100 10732 78140
rect 10772 78100 10781 78140
rect 12931 78100 12940 78140
rect 12980 78100 14380 78140
rect 14420 78100 14572 78140
rect 14612 78100 14621 78140
rect 14755 78100 14764 78140
rect 14804 78100 15244 78140
rect 15284 78100 15293 78140
rect 16963 78100 16972 78140
rect 17012 78100 19372 78140
rect 19412 78100 19421 78140
rect 10243 78099 10301 78100
rect 15052 78056 15092 78100
rect 16963 78099 17021 78100
rect 21424 78056 21504 78076
rect 10339 78016 10348 78056
rect 10388 78016 11980 78056
rect 12020 78016 12029 78056
rect 15043 78016 15052 78056
rect 15092 78016 15101 78056
rect 21388 77996 21504 78056
rect 20803 77972 20861 77973
rect 21388 77972 21428 77996
rect 20803 77932 20812 77972
rect 20852 77932 21428 77972
rect 20803 77931 20861 77932
rect 0 77889 80 77908
rect 0 77888 125 77889
rect 0 77848 76 77888
rect 116 77848 125 77888
rect 4919 77848 4928 77888
rect 4968 77848 5010 77888
rect 5050 77848 5092 77888
rect 5132 77848 5174 77888
rect 5214 77848 5256 77888
rect 5296 77848 5305 77888
rect 20039 77848 20048 77888
rect 20088 77848 20130 77888
rect 20170 77848 20212 77888
rect 20252 77848 20294 77888
rect 20334 77848 20376 77888
rect 20416 77848 20425 77888
rect 0 77847 125 77848
rect 0 77828 80 77847
rect 16003 77764 16012 77804
rect 16052 77764 16300 77804
rect 16340 77764 16349 77804
rect 20515 77720 20573 77721
rect 21424 77720 21504 77740
rect 16195 77680 16204 77720
rect 16244 77680 17068 77720
rect 17108 77680 17117 77720
rect 17731 77680 17740 77720
rect 17780 77680 19660 77720
rect 19700 77680 19709 77720
rect 20515 77680 20524 77720
rect 20564 77680 21504 77720
rect 20515 77679 20573 77680
rect 21424 77660 21504 77680
rect 17059 77636 17117 77637
rect 10243 77596 10252 77636
rect 10292 77596 10924 77636
rect 10964 77596 10973 77636
rect 17059 77596 17068 77636
rect 17108 77596 19276 77636
rect 19316 77596 19325 77636
rect 17059 77595 17117 77596
rect 9187 77512 9196 77552
rect 9236 77512 9868 77552
rect 9908 77512 9917 77552
rect 10051 77512 10060 77552
rect 10100 77512 10348 77552
rect 10388 77512 10397 77552
rect 11320 77512 18508 77552
rect 18548 77512 18557 77552
rect 10435 77468 10493 77469
rect 11320 77468 11360 77512
rect 16579 77468 16637 77469
rect 19747 77468 19805 77469
rect 8803 77428 8812 77468
rect 8852 77428 10444 77468
rect 10484 77428 11360 77468
rect 16387 77428 16396 77468
rect 16436 77428 16588 77468
rect 16628 77428 16637 77468
rect 17251 77428 17260 77468
rect 17300 77428 18988 77468
rect 19028 77428 19037 77468
rect 19747 77428 19756 77468
rect 19796 77428 19852 77468
rect 19892 77428 19901 77468
rect 10435 77427 10493 77428
rect 16579 77427 16637 77428
rect 19747 77427 19805 77428
rect 21424 77384 21504 77404
rect 15427 77344 15436 77384
rect 15476 77344 21504 77384
rect 21424 77324 21504 77344
rect 15715 77260 15724 77300
rect 15764 77260 19084 77300
rect 19124 77260 19133 77300
rect 0 77216 80 77236
rect 1507 77216 1565 77217
rect 17059 77216 17117 77217
rect 0 77176 1516 77216
rect 1556 77176 1565 77216
rect 13027 77176 13036 77216
rect 13076 77176 17068 77216
rect 17108 77176 17117 77216
rect 0 77156 80 77176
rect 1507 77175 1565 77176
rect 17059 77175 17117 77176
rect 3679 77092 3688 77132
rect 3728 77092 3770 77132
rect 3810 77092 3852 77132
rect 3892 77092 3934 77132
rect 3974 77092 4016 77132
rect 4056 77092 4065 77132
rect 18799 77092 18808 77132
rect 18848 77092 18890 77132
rect 18930 77092 18972 77132
rect 19012 77092 19054 77132
rect 19094 77092 19136 77132
rect 19176 77092 19185 77132
rect 21424 77048 21504 77068
rect 20035 77008 20044 77048
rect 20084 77008 21504 77048
rect 21424 76988 21504 77008
rect 13411 76964 13469 76965
rect 10339 76924 10348 76964
rect 10388 76924 11020 76964
rect 11060 76924 11069 76964
rect 13315 76924 13324 76964
rect 13364 76924 13420 76964
rect 13460 76924 13469 76964
rect 16195 76924 16204 76964
rect 16244 76924 17740 76964
rect 17780 76924 17789 76964
rect 13411 76923 13469 76924
rect 8419 76840 8428 76880
rect 8468 76840 8908 76880
rect 8948 76840 8957 76880
rect 9187 76840 9196 76880
rect 9236 76840 9964 76880
rect 10004 76840 10013 76880
rect 12835 76840 12844 76880
rect 12884 76840 13708 76880
rect 13748 76840 15628 76880
rect 15668 76840 15677 76880
rect 16675 76840 16684 76880
rect 16724 76840 17548 76880
rect 17588 76840 17597 76880
rect 19939 76796 19997 76797
rect 4291 76756 4300 76796
rect 4340 76756 18604 76796
rect 18644 76756 18653 76796
rect 19843 76756 19852 76796
rect 19892 76756 19948 76796
rect 19988 76756 19997 76796
rect 19939 76755 19997 76756
rect 8515 76712 8573 76713
rect 8995 76712 9053 76713
rect 13507 76712 13565 76713
rect 21424 76712 21504 76732
rect 8430 76672 8524 76712
rect 8564 76672 8573 76712
rect 8910 76672 9004 76712
rect 9044 76672 9053 76712
rect 9475 76672 9484 76712
rect 9524 76672 11404 76712
rect 11444 76672 11453 76712
rect 13123 76672 13132 76712
rect 13172 76672 13181 76712
rect 13422 76672 13516 76712
rect 13556 76672 13565 76712
rect 14083 76672 14092 76712
rect 14132 76672 16108 76712
rect 16148 76672 16157 76712
rect 18787 76672 18796 76712
rect 18836 76672 21504 76712
rect 8515 76671 8573 76672
rect 8995 76671 9053 76672
rect 12931 76628 12989 76629
rect 8707 76588 8716 76628
rect 8756 76588 12748 76628
rect 12788 76588 12940 76628
rect 12980 76588 12989 76628
rect 13132 76628 13172 76672
rect 13507 76671 13565 76672
rect 21424 76652 21504 76672
rect 13132 76588 15148 76628
rect 15188 76588 15197 76628
rect 16684 76588 17452 76628
rect 17492 76588 18700 76628
rect 18740 76588 18749 76628
rect 12931 76587 12989 76588
rect 0 76544 80 76564
rect 643 76544 701 76545
rect 11011 76544 11069 76545
rect 16684 76544 16724 76588
rect 19459 76544 19517 76545
rect 0 76504 652 76544
rect 692 76504 701 76544
rect 10147 76504 10156 76544
rect 10196 76504 10732 76544
rect 10772 76504 10781 76544
rect 10915 76504 10924 76544
rect 10964 76504 11020 76544
rect 11060 76504 11069 76544
rect 12163 76504 12172 76544
rect 12212 76504 16724 76544
rect 16771 76504 16780 76544
rect 16820 76504 18124 76544
rect 18164 76504 18173 76544
rect 19459 76504 19468 76544
rect 19508 76504 19948 76544
rect 19988 76504 19997 76544
rect 20131 76504 20140 76544
rect 20180 76504 20620 76544
rect 20660 76504 20669 76544
rect 0 76484 80 76504
rect 643 76503 701 76504
rect 11011 76503 11069 76504
rect 19459 76503 19517 76504
rect 19555 76460 19613 76461
rect 11203 76420 11212 76460
rect 11252 76420 18988 76460
rect 19028 76420 19037 76460
rect 19363 76420 19372 76460
rect 19412 76420 19421 76460
rect 19555 76420 19564 76460
rect 19604 76420 20564 76460
rect 4919 76336 4928 76376
rect 4968 76336 5010 76376
rect 5050 76336 5092 76376
rect 5132 76336 5174 76376
rect 5214 76336 5256 76376
rect 5296 76336 5305 76376
rect 6691 76336 6700 76376
rect 6740 76336 15340 76376
rect 15380 76336 15389 76376
rect 10435 76292 10493 76293
rect 12931 76292 12989 76293
rect 19372 76292 19412 76420
rect 19555 76419 19613 76420
rect 20524 76376 20564 76420
rect 21424 76376 21504 76396
rect 19459 76336 19468 76376
rect 19508 76336 19948 76376
rect 19988 76336 19997 76376
rect 20039 76336 20048 76376
rect 20088 76336 20130 76376
rect 20170 76336 20212 76376
rect 20252 76336 20294 76376
rect 20334 76336 20376 76376
rect 20416 76336 20425 76376
rect 20524 76336 21504 76376
rect 21424 76316 21504 76336
rect 10350 76252 10444 76292
rect 10484 76252 10493 76292
rect 10435 76251 10493 76252
rect 11320 76252 11884 76292
rect 11924 76252 12172 76292
rect 12212 76252 12748 76292
rect 12788 76252 12797 76292
rect 12931 76252 12940 76292
rect 12980 76252 13420 76292
rect 13460 76252 13469 76292
rect 19372 76252 19756 76292
rect 19796 76252 19805 76292
rect 8419 76168 8428 76208
rect 8468 76168 8908 76208
rect 8948 76168 8957 76208
rect 11320 76040 11360 76252
rect 12931 76251 12989 76252
rect 11971 76168 11980 76208
rect 12020 76168 12268 76208
rect 12308 76168 13324 76208
rect 13364 76168 13373 76208
rect 14755 76168 14764 76208
rect 14804 76168 15052 76208
rect 15092 76168 15101 76208
rect 16963 76168 16972 76208
rect 17012 76168 17644 76208
rect 17684 76168 17693 76208
rect 19171 76168 19180 76208
rect 19220 76168 20372 76208
rect 12643 76084 12652 76124
rect 12692 76084 13612 76124
rect 13652 76084 13661 76124
rect 19363 76084 19372 76124
rect 19412 76084 19660 76124
rect 19700 76084 19709 76124
rect 15139 76040 15197 76041
rect 20332 76040 20372 76168
rect 21424 76040 21504 76060
rect 7939 76000 7948 76040
rect 7988 76000 9964 76040
rect 10004 76000 10156 76040
rect 10196 76000 11360 76040
rect 11491 76000 11500 76040
rect 11540 76000 15148 76040
rect 15188 76000 15244 76040
rect 15284 76000 15293 76040
rect 17539 76000 17548 76040
rect 17588 76000 18220 76040
rect 18260 76000 18269 76040
rect 20332 76000 21504 76040
rect 15139 75999 15197 76000
rect 21424 75980 21504 76000
rect 18883 75956 18941 75957
rect 15715 75916 15724 75956
rect 15764 75916 16108 75956
rect 16148 75916 16157 75956
rect 18883 75916 18892 75956
rect 18932 75916 19948 75956
rect 19988 75916 19997 75956
rect 18883 75915 18941 75916
rect 0 75872 80 75892
rect 259 75872 317 75873
rect 10339 75872 10397 75873
rect 0 75832 268 75872
rect 308 75832 317 75872
rect 10254 75832 10348 75872
rect 10388 75832 11020 75872
rect 11060 75832 11069 75872
rect 11683 75832 11692 75872
rect 11732 75832 19554 75872
rect 19594 75832 19603 75872
rect 0 75812 80 75832
rect 259 75831 317 75832
rect 10339 75831 10397 75832
rect 17059 75748 17068 75788
rect 17108 75748 17548 75788
rect 17588 75748 17597 75788
rect 19747 75748 19756 75788
rect 19796 75748 20716 75788
rect 20756 75748 20765 75788
rect 12067 75704 12125 75705
rect 19747 75704 19805 75705
rect 21424 75704 21504 75724
rect 10627 75664 10636 75704
rect 10676 75664 12076 75704
rect 12116 75664 12125 75704
rect 19555 75664 19564 75704
rect 19604 75664 19756 75704
rect 19796 75664 19805 75704
rect 20035 75664 20044 75704
rect 20084 75664 21504 75704
rect 12067 75663 12125 75664
rect 19747 75663 19805 75664
rect 21424 75644 21504 75664
rect 3679 75580 3688 75620
rect 3728 75580 3770 75620
rect 3810 75580 3852 75620
rect 3892 75580 3934 75620
rect 3974 75580 4016 75620
rect 4056 75580 4065 75620
rect 9571 75580 9580 75620
rect 9620 75580 10252 75620
rect 10292 75580 10301 75620
rect 14083 75580 14092 75620
rect 14132 75580 16148 75620
rect 17059 75580 17068 75620
rect 17108 75580 17260 75620
rect 17300 75580 17740 75620
rect 17780 75580 17789 75620
rect 18799 75580 18808 75620
rect 18848 75580 18890 75620
rect 18930 75580 18972 75620
rect 19012 75580 19054 75620
rect 19094 75580 19136 75620
rect 19176 75580 19185 75620
rect 13411 75536 13469 75537
rect 16108 75536 16148 75580
rect 19459 75536 19517 75537
rect 12931 75496 12940 75536
rect 12980 75496 13420 75536
rect 13460 75496 15340 75536
rect 15380 75496 15389 75536
rect 15619 75496 15628 75536
rect 15668 75496 16012 75536
rect 16052 75496 16061 75536
rect 16108 75496 19468 75536
rect 19508 75496 20044 75536
rect 20084 75496 20093 75536
rect 13411 75495 13469 75496
rect 19459 75495 19517 75496
rect 6787 75412 6796 75452
rect 6836 75412 7756 75452
rect 7796 75412 18508 75452
rect 18548 75412 18557 75452
rect 21424 75368 21504 75388
rect 8899 75328 8908 75368
rect 8948 75328 9196 75368
rect 9236 75328 9245 75368
rect 10915 75328 10924 75368
rect 10964 75328 16012 75368
rect 16052 75328 16061 75368
rect 20611 75328 20620 75368
rect 20660 75328 21504 75368
rect 21424 75308 21504 75328
rect 12076 75244 14284 75284
rect 14324 75244 14572 75284
rect 14612 75244 14621 75284
rect 15619 75244 15628 75284
rect 15668 75244 16204 75284
rect 16244 75244 16253 75284
rect 16867 75244 16876 75284
rect 16916 75244 18220 75284
rect 18260 75244 18796 75284
rect 18836 75244 18845 75284
rect 0 75200 80 75220
rect 1795 75200 1853 75201
rect 12076 75200 12116 75244
rect 17059 75200 17117 75201
rect 0 75160 1804 75200
rect 1844 75160 1853 75200
rect 10147 75160 10156 75200
rect 10196 75160 10444 75200
rect 10484 75160 10493 75200
rect 11587 75160 11596 75200
rect 11636 75160 12076 75200
rect 12116 75160 12125 75200
rect 13027 75160 13036 75200
rect 13076 75160 13900 75200
rect 13940 75160 13949 75200
rect 16963 75160 16972 75200
rect 17012 75160 17068 75200
rect 17108 75160 17117 75200
rect 0 75140 80 75160
rect 1795 75159 1853 75160
rect 17059 75159 17117 75160
rect 19843 75076 19852 75116
rect 19892 75076 20564 75116
rect 20524 75032 20564 75076
rect 21424 75032 21504 75052
rect 8131 74992 8140 75032
rect 8180 74992 10060 75032
rect 10100 74992 10109 75032
rect 10627 74992 10636 75032
rect 10676 74992 11404 75032
rect 11444 74992 11453 75032
rect 18595 74992 18604 75032
rect 18644 74992 19084 75032
rect 19124 74992 19133 75032
rect 20131 74992 20140 75032
rect 20180 74992 20189 75032
rect 20524 74992 21504 75032
rect 20140 74948 20180 74992
rect 21424 74972 21504 74992
rect 7939 74908 7948 74948
rect 7988 74908 8812 74948
rect 8852 74908 8861 74948
rect 9187 74908 9196 74948
rect 9236 74908 14092 74948
rect 14132 74908 14141 74948
rect 20140 74908 20852 74948
rect 4919 74824 4928 74864
rect 4968 74824 5010 74864
rect 5050 74824 5092 74864
rect 5132 74824 5174 74864
rect 5214 74824 5256 74864
rect 5296 74824 5305 74864
rect 20039 74824 20048 74864
rect 20088 74824 20130 74864
rect 20170 74824 20212 74864
rect 20252 74824 20294 74864
rect 20334 74824 20376 74864
rect 20416 74824 20425 74864
rect 10243 74740 10252 74780
rect 10292 74740 18604 74780
rect 18644 74740 18653 74780
rect 20812 74696 20852 74908
rect 21424 74696 21504 74716
rect 5347 74656 5356 74696
rect 5396 74656 5644 74696
rect 5684 74656 5693 74696
rect 6691 74656 6700 74696
rect 6740 74656 10636 74696
rect 10676 74656 11444 74696
rect 11491 74656 11500 74696
rect 11540 74656 12076 74696
rect 12116 74656 12748 74696
rect 12788 74656 12797 74696
rect 12940 74656 15628 74696
rect 15668 74656 15677 74696
rect 20812 74656 21504 74696
rect 11404 74612 11444 74656
rect 12940 74612 12980 74656
rect 21424 74636 21504 74656
rect 11404 74572 12980 74612
rect 14947 74572 14956 74612
rect 14996 74572 18028 74612
rect 18068 74572 18077 74612
rect 0 74528 80 74548
rect 8611 74528 8669 74529
rect 9379 74528 9437 74529
rect 13507 74528 13565 74529
rect 0 74488 1996 74528
rect 2036 74488 2045 74528
rect 4963 74488 4972 74528
rect 5012 74488 6412 74528
rect 6452 74488 6461 74528
rect 7651 74488 7660 74528
rect 7700 74488 8620 74528
rect 8660 74488 8669 74528
rect 8995 74488 9004 74528
rect 9044 74488 9388 74528
rect 9428 74488 9484 74528
rect 9524 74488 9533 74528
rect 12259 74488 12268 74528
rect 12308 74488 12652 74528
rect 12692 74488 12701 74528
rect 12748 74488 13268 74528
rect 0 74468 80 74488
rect 6412 74360 6452 74488
rect 8611 74487 8669 74488
rect 9379 74487 9437 74488
rect 8803 74444 8861 74445
rect 11875 74444 11933 74445
rect 12748 74444 12788 74488
rect 13228 74444 13268 74488
rect 13507 74488 13516 74528
rect 13556 74488 15340 74528
rect 15380 74488 15389 74528
rect 13507 74487 13565 74488
rect 8803 74404 8812 74444
rect 8852 74404 9100 74444
rect 9140 74404 9149 74444
rect 10819 74404 10828 74444
rect 10868 74404 11884 74444
rect 11924 74404 12788 74444
rect 13123 74404 13132 74444
rect 13172 74404 13181 74444
rect 13228 74404 16108 74444
rect 16148 74404 16157 74444
rect 16963 74404 16972 74444
rect 17012 74404 19852 74444
rect 19892 74404 19901 74444
rect 8803 74403 8861 74404
rect 11875 74403 11933 74404
rect 13132 74360 13172 74404
rect 21424 74360 21504 74380
rect 6412 74320 7660 74360
rect 7700 74320 8044 74360
rect 8084 74320 8093 74360
rect 11875 74320 11884 74360
rect 11924 74320 12556 74360
rect 12596 74320 13172 74360
rect 14371 74320 14380 74360
rect 14420 74320 15820 74360
rect 15860 74320 17260 74360
rect 17300 74320 17309 74360
rect 20707 74320 20716 74360
rect 20756 74320 21504 74360
rect 21424 74300 21504 74320
rect 6595 74236 6604 74276
rect 6644 74236 6988 74276
rect 7028 74236 7037 74276
rect 11971 74236 11980 74276
rect 12020 74236 12268 74276
rect 12308 74236 12317 74276
rect 19747 74236 19756 74276
rect 19796 74236 20044 74276
rect 20084 74236 20093 74276
rect 12739 74152 12748 74192
rect 12788 74152 13804 74192
rect 13844 74152 13853 74192
rect 15811 74152 15820 74192
rect 15860 74152 16108 74192
rect 16148 74152 16157 74192
rect 3679 74068 3688 74108
rect 3728 74068 3770 74108
rect 3810 74068 3852 74108
rect 3892 74068 3934 74108
rect 3974 74068 4016 74108
rect 4056 74068 4065 74108
rect 13411 74068 13420 74108
rect 13460 74068 17164 74108
rect 17204 74068 17213 74108
rect 18799 74068 18808 74108
rect 18848 74068 18890 74108
rect 18930 74068 18972 74108
rect 19012 74068 19054 74108
rect 19094 74068 19136 74108
rect 19176 74068 19185 74108
rect 19267 74068 19276 74108
rect 19316 74068 19325 74108
rect 14188 74024 14228 74068
rect 15139 74024 15197 74025
rect 16291 74024 16349 74025
rect 11779 73984 11788 74024
rect 11828 73984 13460 74024
rect 14179 73984 14188 74024
rect 14228 73984 14268 74024
rect 15043 73984 15052 74024
rect 15092 73984 15148 74024
rect 15188 73984 16300 74024
rect 16340 73984 16349 74024
rect 13420 73940 13460 73984
rect 15139 73983 15197 73984
rect 16291 73983 16349 73984
rect 19276 73940 19316 74068
rect 19939 74024 19997 74025
rect 21424 74024 21504 74044
rect 19939 73984 19948 74024
rect 19988 73984 21504 74024
rect 19939 73983 19997 73984
rect 21424 73964 21504 73984
rect 7843 73900 7852 73940
rect 7892 73900 12020 73940
rect 12355 73900 12364 73940
rect 12404 73900 12940 73940
rect 12980 73900 12989 73940
rect 13411 73900 13420 73940
rect 13460 73900 13469 73940
rect 14851 73900 14860 73940
rect 14900 73900 15244 73940
rect 15284 73900 15293 73940
rect 18883 73900 18892 73940
rect 18932 73900 19316 73940
rect 19843 73940 19901 73941
rect 19843 73900 19852 73940
rect 19892 73900 19948 73940
rect 19988 73900 19997 73940
rect 0 73856 80 73876
rect 5347 73856 5405 73857
rect 6403 73856 6461 73857
rect 11980 73856 12020 73900
rect 19843 73899 19901 73900
rect 0 73816 268 73856
rect 308 73816 317 73856
rect 5347 73816 5356 73856
rect 5396 73816 5452 73856
rect 5492 73816 5501 73856
rect 5923 73816 5932 73856
rect 5972 73816 6412 73856
rect 6452 73816 8908 73856
rect 8948 73816 8957 73856
rect 11971 73816 11980 73856
rect 12020 73816 12652 73856
rect 12692 73816 13228 73856
rect 13268 73816 13277 73856
rect 14275 73816 14284 73856
rect 14324 73816 16300 73856
rect 16340 73816 16349 73856
rect 0 73796 80 73816
rect 5347 73815 5405 73816
rect 6403 73815 6461 73816
rect 8995 73732 9004 73772
rect 9044 73732 9676 73772
rect 9716 73732 9725 73772
rect 11320 73732 19756 73772
rect 19796 73732 19805 73772
rect 6019 73688 6077 73689
rect 8707 73688 8765 73689
rect 9091 73688 9149 73689
rect 5934 73648 6028 73688
rect 6068 73648 6077 73688
rect 8622 73648 8716 73688
rect 8756 73648 8765 73688
rect 9006 73648 9100 73688
rect 9140 73648 9149 73688
rect 9571 73648 9580 73688
rect 9620 73648 11116 73688
rect 11156 73648 11165 73688
rect 6019 73647 6077 73648
rect 8707 73647 8765 73648
rect 9091 73647 9149 73648
rect 11320 73604 11360 73732
rect 18691 73688 18749 73689
rect 21424 73688 21504 73708
rect 14659 73648 14668 73688
rect 14708 73648 15340 73688
rect 15380 73648 16588 73688
rect 16628 73648 16637 73688
rect 18595 73648 18604 73688
rect 18644 73648 18700 73688
rect 18740 73648 18749 73688
rect 19171 73648 19180 73688
rect 19220 73648 21504 73688
rect 18691 73647 18749 73648
rect 21424 73628 21504 73648
rect 5155 73564 5164 73604
rect 5204 73564 5452 73604
rect 5492 73564 5501 73604
rect 8227 73564 8236 73604
rect 8276 73564 11360 73604
rect 11875 73604 11933 73605
rect 11875 73564 11884 73604
rect 11924 73564 11980 73604
rect 12020 73564 12029 73604
rect 13123 73564 13132 73604
rect 13172 73564 14284 73604
rect 14324 73564 14333 73604
rect 16195 73564 16204 73604
rect 16244 73564 18412 73604
rect 18452 73564 18700 73604
rect 18740 73564 18749 73604
rect 11875 73563 11933 73564
rect 11491 73396 11500 73436
rect 11540 73396 11788 73436
rect 11828 73396 11837 73436
rect 12451 73396 12460 73436
rect 12500 73396 13036 73436
rect 13076 73396 13708 73436
rect 13748 73396 13757 73436
rect 21424 73352 21504 73372
rect 4919 73312 4928 73352
rect 4968 73312 5010 73352
rect 5050 73312 5092 73352
rect 5132 73312 5174 73352
rect 5214 73312 5256 73352
rect 5296 73312 5305 73352
rect 20039 73312 20048 73352
rect 20088 73312 20130 73352
rect 20170 73312 20212 73352
rect 20252 73312 20294 73352
rect 20334 73312 20376 73352
rect 20416 73312 20425 73352
rect 20524 73312 21504 73352
rect 18115 73268 18173 73269
rect 18030 73228 18124 73268
rect 18164 73228 18173 73268
rect 18115 73227 18173 73228
rect 0 73184 80 73204
rect 12259 73184 12317 73185
rect 0 73144 1900 73184
rect 1940 73144 1949 73184
rect 10339 73144 10348 73184
rect 10388 73144 10580 73184
rect 0 73124 80 73144
rect 7651 73060 7660 73100
rect 7700 73060 7852 73100
rect 7892 73060 7901 73100
rect 10020 73060 10060 73100
rect 10100 73060 10109 73100
rect 10060 73016 10100 73060
rect 10540 73016 10580 73144
rect 12259 73144 12268 73184
rect 12308 73144 19372 73184
rect 19412 73144 19421 73184
rect 12259 73143 12317 73144
rect 17923 73100 17981 73101
rect 20131 73100 20189 73101
rect 20524 73100 20564 73312
rect 21424 73292 21504 73312
rect 13795 73060 13804 73100
rect 13844 73060 16300 73100
rect 16340 73060 17164 73100
rect 17204 73060 17213 73100
rect 17838 73060 17932 73100
rect 17972 73060 17981 73100
rect 18948 73060 18988 73100
rect 19028 73060 19037 73100
rect 20131 73060 20140 73100
rect 20180 73060 20564 73100
rect 17923 73059 17981 73060
rect 12259 73016 12317 73017
rect 18988 73016 19028 73060
rect 20131 73059 20189 73060
rect 21424 73016 21504 73036
rect 8515 72976 8524 73016
rect 8564 72976 10100 73016
rect 10339 72976 10348 73016
rect 10388 72976 10924 73016
rect 10964 72976 10973 73016
rect 11395 72976 11404 73016
rect 11444 72976 12268 73016
rect 12308 72976 12317 73016
rect 12259 72975 12317 72976
rect 15052 72976 15628 73016
rect 15668 72976 15916 73016
rect 15956 72976 15965 73016
rect 18403 72976 18412 73016
rect 18452 72976 19028 73016
rect 19555 72976 19564 73016
rect 19604 72976 21504 73016
rect 11587 72932 11645 72933
rect 15052 72932 15092 72976
rect 21424 72956 21504 72976
rect 20131 72932 20189 72933
rect 7843 72892 7852 72932
rect 7892 72892 8332 72932
rect 8372 72892 8381 72932
rect 8803 72892 8812 72932
rect 8852 72892 11020 72932
rect 11060 72892 11069 72932
rect 11587 72892 11596 72932
rect 11636 72892 15092 72932
rect 15139 72892 15148 72932
rect 15188 72892 18988 72932
rect 19028 72892 19037 72932
rect 19084 72892 20140 72932
rect 20180 72892 20189 72932
rect 11587 72891 11645 72892
rect 17155 72848 17213 72849
rect 18115 72848 18173 72849
rect 19084 72848 19124 72892
rect 20131 72891 20189 72892
rect 21379 72848 21437 72849
rect 10147 72808 10156 72848
rect 10196 72808 12076 72848
rect 12116 72808 12125 72848
rect 17155 72808 17164 72848
rect 17204 72808 17260 72848
rect 17300 72808 17309 72848
rect 18030 72808 18124 72848
rect 18164 72808 18173 72848
rect 18787 72808 18796 72848
rect 18836 72808 19124 72848
rect 19171 72808 19180 72848
rect 19220 72808 21388 72848
rect 21428 72808 21437 72848
rect 17155 72807 17213 72808
rect 18115 72807 18173 72808
rect 21379 72807 21437 72808
rect 1507 72724 1516 72764
rect 1556 72724 3916 72764
rect 3956 72724 4108 72764
rect 4148 72724 4157 72764
rect 7651 72724 7660 72764
rect 7700 72724 11732 72764
rect 11779 72724 11788 72764
rect 11828 72724 13612 72764
rect 13652 72724 13661 72764
rect 13708 72724 19756 72764
rect 19796 72724 19805 72764
rect 3679 72556 3688 72596
rect 3728 72556 3770 72596
rect 3810 72556 3852 72596
rect 3892 72556 3934 72596
rect 3974 72556 4016 72596
rect 4056 72556 4065 72596
rect 0 72512 80 72532
rect 163 72512 221 72513
rect 0 72472 172 72512
rect 212 72472 221 72512
rect 4108 72512 4148 72724
rect 11587 72680 11645 72681
rect 10339 72640 10348 72680
rect 10388 72640 10636 72680
rect 10676 72640 10685 72680
rect 11011 72640 11020 72680
rect 11060 72640 11596 72680
rect 11636 72640 11645 72680
rect 11692 72680 11732 72724
rect 13708 72680 13748 72724
rect 21424 72680 21504 72700
rect 11692 72640 13748 72680
rect 19459 72640 19468 72680
rect 19508 72640 21504 72680
rect 11587 72639 11645 72640
rect 21424 72620 21504 72640
rect 8323 72556 8332 72596
rect 8372 72556 18604 72596
rect 18644 72556 18653 72596
rect 18799 72556 18808 72596
rect 18848 72556 18890 72596
rect 18930 72556 18972 72596
rect 19012 72556 19054 72596
rect 19094 72556 19136 72596
rect 19176 72556 19185 72596
rect 4108 72472 19028 72512
rect 0 72452 80 72472
rect 163 72471 221 72472
rect 18691 72428 18749 72429
rect 18988 72428 19028 72472
rect 2467 72388 2476 72428
rect 2516 72388 3436 72428
rect 3476 72388 9964 72428
rect 10004 72388 11596 72428
rect 11636 72388 11645 72428
rect 18691 72388 18700 72428
rect 18740 72388 18796 72428
rect 18836 72388 18845 72428
rect 18979 72388 18988 72428
rect 19028 72388 19037 72428
rect 18691 72387 18749 72388
rect 21424 72344 21504 72364
rect 1315 72304 1324 72344
rect 1364 72304 2540 72344
rect 2500 72260 2540 72304
rect 11320 72304 15148 72344
rect 15188 72304 15197 72344
rect 16387 72304 16396 72344
rect 16436 72304 16972 72344
rect 17012 72304 17021 72344
rect 19651 72304 19660 72344
rect 19700 72304 21504 72344
rect 4291 72260 4349 72261
rect 11320 72260 11360 72304
rect 21424 72284 21504 72304
rect 19747 72260 19805 72261
rect 2500 72220 4300 72260
rect 4340 72220 11360 72260
rect 13219 72220 13228 72260
rect 13268 72220 15188 72260
rect 15235 72220 15244 72260
rect 15284 72220 19372 72260
rect 19412 72220 19421 72260
rect 19662 72220 19756 72260
rect 19796 72220 19805 72260
rect 4291 72219 4349 72220
rect 15148 72176 15188 72220
rect 19747 72219 19805 72220
rect 19939 72260 19997 72261
rect 19939 72220 19948 72260
rect 19988 72220 20082 72260
rect 19939 72219 19997 72220
rect 16483 72176 16541 72177
rect 5539 72136 5548 72176
rect 5588 72136 7180 72176
rect 7220 72136 7229 72176
rect 7555 72136 7564 72176
rect 7604 72136 12748 72176
rect 12788 72136 13132 72176
rect 13172 72136 13181 72176
rect 13891 72136 13900 72176
rect 13940 72136 14956 72176
rect 14996 72136 15005 72176
rect 15139 72136 15148 72176
rect 15188 72136 15340 72176
rect 15380 72136 15389 72176
rect 16483 72136 16492 72176
rect 16532 72136 20756 72176
rect 16483 72135 16541 72136
rect 13699 72052 13708 72092
rect 13748 72052 17836 72092
rect 17876 72052 17885 72092
rect 20140 72052 20620 72092
rect 20660 72052 20669 72092
rect 17155 72008 17213 72009
rect 17836 72008 17876 72052
rect 20140 72008 20180 72052
rect 5155 71968 5164 72008
rect 5204 71968 5396 72008
rect 7363 71968 7372 72008
rect 7412 71968 8140 72008
rect 8180 71968 8189 72008
rect 11587 71968 11596 72008
rect 11636 71968 13228 72008
rect 13268 71968 13277 72008
rect 13411 71968 13420 72008
rect 13460 71968 13996 72008
rect 14036 71968 14045 72008
rect 15523 71968 15532 72008
rect 15572 71968 16108 72008
rect 16148 71968 16157 72008
rect 17155 71968 17164 72008
rect 17204 71968 17260 72008
rect 17300 71968 17309 72008
rect 17836 71968 18412 72008
rect 18452 71968 18461 72008
rect 19555 71968 19564 72008
rect 19604 71968 20180 72008
rect 20716 72008 20756 72136
rect 21424 72008 21504 72028
rect 20716 71968 21504 72008
rect 0 71840 80 71860
rect 1891 71840 1949 71841
rect 0 71800 1900 71840
rect 1940 71800 1949 71840
rect 4919 71800 4928 71840
rect 4968 71800 5010 71840
rect 5050 71800 5092 71840
rect 5132 71800 5174 71840
rect 5214 71800 5256 71840
rect 5296 71800 5305 71840
rect 0 71780 80 71800
rect 1891 71799 1949 71800
rect 5356 71756 5396 71968
rect 17155 71967 17213 71968
rect 21424 71948 21504 71968
rect 14851 71840 14909 71841
rect 15427 71840 15485 71841
rect 7372 71800 10348 71840
rect 10388 71800 10397 71840
rect 13891 71800 13900 71840
rect 13940 71800 14188 71840
rect 14228 71800 14237 71840
rect 14851 71800 14860 71840
rect 14900 71800 15052 71840
rect 15092 71800 15101 71840
rect 15331 71800 15340 71840
rect 15380 71800 15436 71840
rect 15476 71800 15485 71840
rect 17731 71800 17740 71840
rect 17780 71800 18508 71840
rect 18548 71800 18557 71840
rect 20039 71800 20048 71840
rect 20088 71800 20130 71840
rect 20170 71800 20212 71840
rect 20252 71800 20294 71840
rect 20334 71800 20376 71840
rect 20416 71800 20425 71840
rect 7372 71756 7412 71800
rect 14851 71799 14909 71800
rect 15427 71799 15485 71800
rect 5356 71716 5492 71756
rect 7075 71716 7084 71756
rect 7124 71716 7372 71756
rect 7412 71716 7421 71756
rect 8419 71716 8428 71756
rect 8468 71716 18892 71756
rect 18932 71716 18941 71756
rect 5347 71588 5405 71589
rect 5059 71548 5068 71588
rect 5108 71548 5356 71588
rect 5396 71548 5405 71588
rect 5347 71547 5405 71548
rect 4579 71464 4588 71504
rect 4628 71464 5356 71504
rect 5396 71464 5405 71504
rect 5452 71420 5492 71716
rect 19939 71672 19997 71673
rect 21424 71672 21504 71692
rect 13708 71632 15188 71672
rect 15715 71632 15724 71672
rect 15764 71632 19468 71672
rect 19508 71632 19517 71672
rect 19939 71632 19948 71672
rect 19988 71632 21504 71672
rect 13708 71588 13748 71632
rect 15148 71588 15188 71632
rect 19939 71631 19997 71632
rect 21424 71612 21504 71632
rect 7171 71548 7180 71588
rect 7220 71548 9676 71588
rect 9716 71548 9725 71588
rect 10723 71548 10732 71588
rect 10772 71548 11116 71588
rect 11156 71548 11165 71588
rect 13699 71548 13708 71588
rect 13748 71548 13757 71588
rect 14755 71548 14764 71588
rect 14804 71548 15052 71588
rect 15092 71548 15101 71588
rect 15148 71548 17356 71588
rect 17396 71548 17405 71588
rect 9283 71504 9341 71505
rect 15427 71504 15485 71505
rect 16291 71504 16349 71505
rect 5731 71464 5740 71504
rect 5780 71464 6604 71504
rect 6644 71464 6653 71504
rect 7267 71464 7276 71504
rect 7316 71464 7660 71504
rect 7700 71464 7709 71504
rect 9091 71464 9100 71504
rect 9140 71464 9292 71504
rect 9332 71464 9341 71504
rect 13027 71464 13036 71504
rect 13076 71464 14476 71504
rect 14516 71464 14525 71504
rect 15427 71464 15436 71504
rect 15476 71464 15532 71504
rect 15572 71464 15581 71504
rect 15907 71464 15916 71504
rect 15956 71464 16300 71504
rect 16340 71464 16349 71504
rect 16675 71464 16684 71504
rect 16724 71464 17452 71504
rect 17492 71464 17501 71504
rect 9283 71463 9341 71464
rect 15427 71463 15485 71464
rect 16291 71463 16349 71464
rect 5251 71380 5260 71420
rect 5300 71380 5492 71420
rect 6307 71380 6316 71420
rect 6356 71380 8524 71420
rect 8564 71380 8573 71420
rect 12355 71380 12364 71420
rect 12404 71380 19948 71420
rect 19988 71380 19997 71420
rect 11875 71336 11933 71337
rect 21424 71336 21504 71356
rect 11875 71296 11884 71336
rect 11924 71296 12460 71336
rect 12500 71296 14092 71336
rect 14132 71296 14141 71336
rect 15139 71296 15148 71336
rect 15188 71296 17164 71336
rect 17204 71296 18988 71336
rect 19028 71296 19037 71336
rect 19651 71296 19660 71336
rect 19700 71296 21504 71336
rect 11875 71295 11933 71296
rect 21424 71276 21504 71296
rect 16483 71252 16541 71253
rect 5155 71212 5164 71252
rect 5204 71212 6604 71252
rect 6644 71212 7180 71252
rect 7220 71212 7229 71252
rect 8707 71212 8716 71252
rect 8756 71212 16492 71252
rect 16532 71212 16541 71252
rect 18883 71212 18892 71252
rect 18932 71212 19372 71252
rect 19412 71212 19421 71252
rect 16483 71211 16541 71212
rect 0 71168 80 71188
rect 355 71168 413 71169
rect 17923 71168 17981 71169
rect 0 71128 364 71168
rect 404 71128 413 71168
rect 11971 71128 11980 71168
rect 12020 71128 17932 71168
rect 17972 71128 17981 71168
rect 0 71108 80 71128
rect 355 71127 413 71128
rect 17923 71127 17981 71128
rect 14851 71084 14909 71085
rect 3679 71044 3688 71084
rect 3728 71044 3770 71084
rect 3810 71044 3852 71084
rect 3892 71044 3934 71084
rect 3974 71044 4016 71084
rect 4056 71044 4065 71084
rect 14766 71044 14860 71084
rect 14900 71044 14909 71084
rect 18799 71044 18808 71084
rect 18848 71044 18890 71084
rect 18930 71044 18972 71084
rect 19012 71044 19054 71084
rect 19094 71044 19136 71084
rect 19176 71044 19185 71084
rect 14851 71043 14909 71044
rect 17059 71000 17117 71001
rect 21424 71000 21504 71020
rect 5443 70960 5452 71000
rect 5492 70960 6124 71000
rect 6164 70960 6173 71000
rect 6883 70960 6892 71000
rect 6932 70960 11980 71000
rect 12020 70960 12029 71000
rect 12643 70960 12652 71000
rect 12692 70960 17068 71000
rect 17108 70960 17740 71000
rect 17780 70960 17789 71000
rect 20611 70960 20620 71000
rect 20660 70960 21504 71000
rect 17059 70959 17117 70960
rect 21424 70940 21504 70960
rect 8707 70876 8716 70916
rect 8756 70876 10540 70916
rect 10580 70876 10589 70916
rect 13699 70876 13708 70916
rect 13748 70876 14188 70916
rect 14228 70876 14237 70916
rect 14851 70876 14860 70916
rect 14900 70876 19180 70916
rect 19220 70876 19229 70916
rect 17635 70832 17693 70833
rect 2275 70792 2284 70832
rect 2324 70792 7276 70832
rect 7316 70792 7325 70832
rect 17155 70792 17164 70832
rect 17204 70792 17356 70832
rect 17396 70792 17405 70832
rect 17550 70792 17644 70832
rect 17684 70792 17693 70832
rect 19939 70792 19948 70832
rect 19988 70792 21388 70832
rect 21428 70792 21437 70832
rect 17635 70791 17693 70792
rect 9859 70748 9917 70749
rect 2947 70708 2956 70748
rect 2996 70708 4012 70748
rect 4052 70708 5452 70748
rect 5492 70708 8236 70748
rect 8276 70708 8285 70748
rect 8995 70708 9004 70748
rect 9044 70708 9580 70748
rect 9620 70708 9868 70748
rect 9908 70708 9917 70748
rect 9859 70707 9917 70708
rect 13411 70748 13469 70749
rect 13411 70708 13420 70748
rect 13460 70708 19756 70748
rect 19796 70708 19805 70748
rect 13411 70707 13469 70708
rect 5539 70664 5597 70665
rect 21424 70664 21504 70684
rect 3523 70624 3532 70664
rect 3572 70624 5548 70664
rect 5588 70624 5644 70664
rect 5684 70624 5693 70664
rect 7267 70624 7276 70664
rect 7316 70624 9196 70664
rect 9236 70624 9264 70664
rect 9667 70624 9676 70664
rect 9716 70624 11596 70664
rect 11636 70624 16204 70664
rect 16244 70624 16253 70664
rect 17347 70624 17356 70664
rect 17396 70624 17932 70664
rect 17972 70624 17981 70664
rect 20035 70624 20044 70664
rect 20084 70624 21504 70664
rect 5539 70623 5597 70624
rect 5251 70540 5260 70580
rect 5300 70540 5836 70580
rect 5876 70540 6892 70580
rect 6932 70540 7468 70580
rect 7508 70540 7517 70580
rect 7651 70540 7660 70580
rect 7700 70540 8840 70580
rect 0 70496 80 70516
rect 4483 70496 4541 70497
rect 8800 70496 8840 70540
rect 0 70456 844 70496
rect 884 70456 893 70496
rect 3811 70456 3820 70496
rect 3860 70456 4300 70496
rect 4340 70456 4349 70496
rect 4483 70456 4492 70496
rect 4532 70456 5068 70496
rect 5108 70456 5117 70496
rect 8800 70456 9004 70496
rect 9044 70456 9053 70496
rect 0 70436 80 70456
rect 4483 70455 4541 70456
rect 9100 70412 9140 70624
rect 21424 70604 21504 70624
rect 14083 70580 14141 70581
rect 14851 70580 14909 70581
rect 16099 70580 16157 70581
rect 13998 70540 14092 70580
rect 14132 70540 14141 70580
rect 14766 70540 14860 70580
rect 14900 70540 14909 70580
rect 16014 70540 16108 70580
rect 16148 70540 16157 70580
rect 17155 70540 17164 70580
rect 17204 70540 17740 70580
rect 17780 70540 17789 70580
rect 20131 70540 20140 70580
rect 20180 70540 20189 70580
rect 14083 70539 14141 70540
rect 14851 70539 14909 70540
rect 16099 70539 16157 70540
rect 20140 70496 20180 70540
rect 14755 70456 14764 70496
rect 14804 70456 15148 70496
rect 15188 70456 15197 70496
rect 15331 70456 15340 70496
rect 15380 70456 15628 70496
rect 15668 70456 15677 70496
rect 20140 70456 21332 70496
rect 1315 70372 1324 70412
rect 1364 70372 4396 70412
rect 4436 70372 4445 70412
rect 4579 70372 4588 70412
rect 4628 70372 5548 70412
rect 5588 70372 5597 70412
rect 8899 70372 8908 70412
rect 8948 70372 9140 70412
rect 21292 70328 21332 70456
rect 21424 70328 21504 70348
rect 3619 70288 3628 70328
rect 3668 70288 4204 70328
rect 4244 70288 4253 70328
rect 4919 70288 4928 70328
rect 4968 70288 5010 70328
rect 5050 70288 5092 70328
rect 5132 70288 5174 70328
rect 5214 70288 5256 70328
rect 5296 70288 5305 70328
rect 20039 70288 20048 70328
rect 20088 70288 20130 70328
rect 20170 70288 20212 70328
rect 20252 70288 20294 70328
rect 20334 70288 20376 70328
rect 20416 70288 20425 70328
rect 21292 70288 21504 70328
rect 21424 70268 21504 70288
rect 3532 70204 4492 70244
rect 4532 70204 4541 70244
rect 17347 70204 17356 70244
rect 17396 70204 19372 70244
rect 19412 70204 19421 70244
rect 3532 70076 3572 70204
rect 4387 70120 4396 70160
rect 4436 70120 4972 70160
rect 5012 70120 5021 70160
rect 10531 70120 10540 70160
rect 10580 70120 11212 70160
rect 11252 70120 11261 70160
rect 16963 70076 17021 70077
rect 2467 70036 2476 70076
rect 2516 70036 3572 70076
rect 8227 70036 8236 70076
rect 8276 70036 16972 70076
rect 17012 70036 17021 70076
rect 16963 70035 17021 70036
rect 17836 70036 18124 70076
rect 18164 70036 18173 70076
rect 19651 70036 19660 70076
rect 19700 70036 20044 70076
rect 20084 70036 20093 70076
rect 6595 69992 6653 69993
rect 8323 69992 8381 69993
rect 1507 69952 1516 69992
rect 1556 69952 4492 69992
rect 4532 69952 4541 69992
rect 6019 69952 6028 69992
rect 6068 69952 6220 69992
rect 6260 69952 6604 69992
rect 6644 69952 6653 69992
rect 7747 69952 7756 69992
rect 7796 69952 8332 69992
rect 8372 69952 8428 69992
rect 8468 69952 8477 69992
rect 13507 69952 13516 69992
rect 13556 69952 13900 69992
rect 13940 69952 14380 69992
rect 14420 69952 14429 69992
rect 15427 69952 15436 69992
rect 15476 69952 15724 69992
rect 15764 69952 16588 69992
rect 16628 69952 17740 69992
rect 17780 69952 17789 69992
rect 6595 69951 6653 69952
rect 8323 69951 8381 69952
rect 14947 69908 15005 69909
rect 10723 69868 10732 69908
rect 10772 69868 10924 69908
rect 10964 69868 10973 69908
rect 14862 69868 14956 69908
rect 14996 69868 15005 69908
rect 14947 69867 15005 69868
rect 15139 69908 15197 69909
rect 17836 69908 17876 70036
rect 21424 69992 21504 70012
rect 17923 69952 17932 69992
rect 17972 69952 21504 69992
rect 21424 69932 21504 69952
rect 15139 69868 15148 69908
rect 15188 69868 16108 69908
rect 16148 69868 17876 69908
rect 15139 69867 15197 69868
rect 0 69824 80 69844
rect 2179 69824 2237 69825
rect 0 69784 2188 69824
rect 2228 69784 2237 69824
rect 0 69764 80 69784
rect 2179 69783 2237 69784
rect 15811 69824 15869 69825
rect 16483 69824 16541 69825
rect 15811 69784 15820 69824
rect 15860 69784 16204 69824
rect 16244 69784 16253 69824
rect 16483 69784 16492 69824
rect 16532 69784 17260 69824
rect 17300 69784 18220 69824
rect 18260 69784 18269 69824
rect 15811 69783 15869 69784
rect 16483 69783 16541 69784
rect 17923 69740 17981 69741
rect 6019 69700 6028 69740
rect 6068 69700 6796 69740
rect 6836 69700 6845 69740
rect 14947 69700 14956 69740
rect 14996 69700 15148 69740
rect 15188 69700 15197 69740
rect 17923 69700 17932 69740
rect 17972 69700 18124 69740
rect 18164 69700 18173 69740
rect 20131 69700 20140 69740
rect 20180 69700 20620 69740
rect 20660 69700 20669 69740
rect 17923 69699 17981 69700
rect 21424 69656 21504 69676
rect 20035 69616 20044 69656
rect 20084 69616 21504 69656
rect 21424 69596 21504 69616
rect 3679 69532 3688 69572
rect 3728 69532 3770 69572
rect 3810 69532 3852 69572
rect 3892 69532 3934 69572
rect 3974 69532 4016 69572
rect 4056 69532 4065 69572
rect 18799 69532 18808 69572
rect 18848 69532 18890 69572
rect 18930 69532 18972 69572
rect 19012 69532 19054 69572
rect 19094 69532 19136 69572
rect 19176 69532 19185 69572
rect 19747 69448 19756 69488
rect 19796 69448 20044 69488
rect 20084 69448 20093 69488
rect 13987 69364 13996 69404
rect 14036 69364 14045 69404
rect 19459 69364 19468 69404
rect 19508 69364 20564 69404
rect 4099 69320 4157 69321
rect 8995 69320 9053 69321
rect 13996 69320 14036 69364
rect 4099 69280 4108 69320
rect 4148 69280 4684 69320
rect 4724 69280 4733 69320
rect 5635 69280 5644 69320
rect 5684 69280 5932 69320
rect 5972 69280 5981 69320
rect 7843 69280 7852 69320
rect 7892 69280 9004 69320
rect 9044 69280 11116 69320
rect 11156 69280 11165 69320
rect 12547 69280 12556 69320
rect 12596 69280 14036 69320
rect 17443 69320 17501 69321
rect 20524 69320 20564 69364
rect 21424 69320 21504 69340
rect 17443 69280 17452 69320
rect 17492 69280 17836 69320
rect 17876 69280 17885 69320
rect 19363 69280 19372 69320
rect 19412 69280 19756 69320
rect 19796 69280 19805 69320
rect 20524 69280 21504 69320
rect 4099 69279 4157 69280
rect 8995 69279 9053 69280
rect 17443 69279 17501 69280
rect 21424 69260 21504 69280
rect 15619 69236 15677 69237
rect 18019 69236 18077 69237
rect 7075 69196 7084 69236
rect 7124 69196 8332 69236
rect 8372 69196 8381 69236
rect 10051 69196 10060 69236
rect 10100 69196 10636 69236
rect 10676 69196 10685 69236
rect 15619 69196 15628 69236
rect 15668 69196 16108 69236
rect 16148 69196 16157 69236
rect 17731 69196 17740 69236
rect 17780 69196 18028 69236
rect 18068 69196 18077 69236
rect 15619 69195 15677 69196
rect 18019 69195 18077 69196
rect 0 69152 80 69172
rect 547 69152 605 69153
rect 4483 69152 4541 69153
rect 5635 69152 5693 69153
rect 0 69112 556 69152
rect 596 69112 605 69152
rect 2947 69112 2956 69152
rect 2996 69112 3532 69152
rect 3572 69112 3581 69152
rect 3907 69112 3916 69152
rect 3956 69112 4492 69152
rect 4532 69112 4541 69152
rect 4771 69112 4780 69152
rect 4820 69112 4972 69152
rect 5012 69112 5644 69152
rect 5684 69112 5693 69152
rect 6595 69112 6604 69152
rect 6644 69112 7180 69152
rect 7220 69112 7372 69152
rect 7412 69112 7421 69152
rect 9187 69112 9196 69152
rect 9236 69112 10732 69152
rect 10772 69112 10781 69152
rect 11875 69112 11884 69152
rect 11924 69112 12268 69152
rect 12308 69112 12317 69152
rect 12739 69112 12748 69152
rect 12788 69112 13132 69152
rect 13172 69112 13181 69152
rect 13699 69112 13708 69152
rect 13748 69112 16876 69152
rect 16916 69112 16925 69152
rect 18883 69112 18892 69152
rect 18932 69112 19948 69152
rect 19988 69112 19997 69152
rect 0 69092 80 69112
rect 547 69111 605 69112
rect 4483 69111 4541 69112
rect 5635 69111 5693 69112
rect 3427 69028 3436 69068
rect 3476 69028 4012 69068
rect 4052 69028 9772 69068
rect 9812 69028 9821 69068
rect 14188 69028 14668 69068
rect 14708 69028 18700 69068
rect 18740 69028 18749 69068
rect 14188 68984 14228 69028
rect 17635 68984 17693 68985
rect 21424 68984 21504 69004
rect 4579 68944 4588 68984
rect 4628 68944 10156 68984
rect 10196 68944 10205 68984
rect 10339 68944 10348 68984
rect 10388 68944 10636 68984
rect 10676 68944 10685 68984
rect 14179 68944 14188 68984
rect 14228 68944 14237 68984
rect 15139 68944 15148 68984
rect 15188 68944 16684 68984
rect 16724 68944 16733 68984
rect 16963 68944 16972 68984
rect 17012 68944 17356 68984
rect 17396 68944 17405 68984
rect 17635 68944 17644 68984
rect 17684 68944 17740 68984
rect 17780 68944 17789 68984
rect 20035 68944 20044 68984
rect 20084 68944 20180 68984
rect 21379 68944 21388 68984
rect 21428 68944 21504 68984
rect 17635 68943 17693 68944
rect 20140 68900 20180 68944
rect 21424 68924 21504 68944
rect 20140 68860 20852 68900
rect 4919 68776 4928 68816
rect 4968 68776 5010 68816
rect 5050 68776 5092 68816
rect 5132 68776 5174 68816
rect 5214 68776 5256 68816
rect 5296 68776 5305 68816
rect 20039 68776 20048 68816
rect 20088 68776 20130 68816
rect 20170 68776 20212 68816
rect 20252 68776 20294 68816
rect 20334 68776 20376 68816
rect 20416 68776 20425 68816
rect 10915 68732 10973 68733
rect 20707 68732 20765 68733
rect 3331 68692 3340 68732
rect 3380 68692 3916 68732
rect 3956 68692 3965 68732
rect 5347 68692 5356 68732
rect 5396 68692 5588 68732
rect 5548 68648 5588 68692
rect 10915 68692 10924 68732
rect 10964 68692 20716 68732
rect 20756 68692 20765 68732
rect 10915 68691 10973 68692
rect 20707 68691 20765 68692
rect 15043 68648 15101 68649
rect 15427 68648 15485 68649
rect 5539 68608 5548 68648
rect 5588 68608 5597 68648
rect 15043 68608 15052 68648
rect 15092 68608 15436 68648
rect 15476 68608 15485 68648
rect 15043 68607 15101 68608
rect 15427 68607 15485 68608
rect 17635 68648 17693 68649
rect 20812 68648 20852 68860
rect 21424 68648 21504 68668
rect 17635 68608 17644 68648
rect 17684 68608 18124 68648
rect 18164 68608 18173 68648
rect 20812 68608 21504 68648
rect 17635 68607 17693 68608
rect 21424 68588 21504 68608
rect 6883 68524 6892 68564
rect 6932 68524 6972 68564
rect 8035 68524 8044 68564
rect 8084 68524 18892 68564
rect 18932 68524 18941 68564
rect 0 68480 80 68500
rect 739 68480 797 68481
rect 6892 68480 6932 68524
rect 0 68440 748 68480
rect 788 68440 797 68480
rect 6403 68440 6412 68480
rect 6452 68440 7564 68480
rect 7604 68440 7613 68480
rect 8227 68440 8236 68480
rect 8276 68440 8285 68480
rect 9475 68440 9484 68480
rect 9524 68440 9676 68480
rect 9716 68440 9725 68480
rect 9955 68440 9964 68480
rect 10004 68440 10252 68480
rect 10292 68440 10732 68480
rect 10772 68440 10781 68480
rect 10915 68440 10924 68480
rect 10964 68440 11212 68480
rect 11252 68440 11261 68480
rect 12739 68440 12748 68480
rect 12788 68440 14764 68480
rect 14804 68440 15340 68480
rect 15380 68440 15389 68480
rect 16579 68440 16588 68480
rect 16628 68440 17740 68480
rect 17780 68440 17789 68480
rect 17923 68440 17932 68480
rect 17972 68440 18412 68480
rect 18452 68440 18700 68480
rect 18740 68440 18749 68480
rect 0 68420 80 68440
rect 739 68439 797 68440
rect 4099 68396 4157 68397
rect 6787 68396 6845 68397
rect 8236 68396 8276 68440
rect 3907 68356 3916 68396
rect 3956 68356 4108 68396
rect 4148 68356 4157 68396
rect 6702 68356 6796 68396
rect 6836 68356 7276 68396
rect 7316 68356 7325 68396
rect 7852 68356 8620 68396
rect 8660 68356 8669 68396
rect 9859 68356 9868 68396
rect 9908 68356 19564 68396
rect 19604 68356 19613 68396
rect 4099 68355 4157 68356
rect 6787 68355 6845 68356
rect 7852 68228 7892 68356
rect 11395 68312 11453 68313
rect 14083 68312 14141 68313
rect 21424 68312 21504 68332
rect 8995 68272 9004 68312
rect 9044 68272 11404 68312
rect 11444 68272 11692 68312
rect 11732 68272 11741 68312
rect 13998 68272 14092 68312
rect 14132 68272 14141 68312
rect 15331 68272 15340 68312
rect 15380 68272 16972 68312
rect 17012 68272 19084 68312
rect 19124 68272 19372 68312
rect 19412 68272 19421 68312
rect 20035 68272 20044 68312
rect 20084 68272 21504 68312
rect 11395 68271 11453 68272
rect 14083 68271 14141 68272
rect 21424 68252 21504 68272
rect 14563 68228 14621 68229
rect 3619 68188 3628 68228
rect 3668 68188 3677 68228
rect 7843 68188 7852 68228
rect 7892 68188 7901 68228
rect 11320 68188 14572 68228
rect 14612 68188 14621 68228
rect 15523 68188 15532 68228
rect 15572 68188 16204 68228
rect 16244 68188 16253 68228
rect 3628 68144 3668 68188
rect 11320 68144 11360 68188
rect 14563 68187 14621 68188
rect 17635 68144 17693 68145
rect 3628 68104 11360 68144
rect 11587 68104 11596 68144
rect 11636 68104 12172 68144
rect 12212 68104 12221 68144
rect 17550 68104 17644 68144
rect 17684 68104 17693 68144
rect 17635 68103 17693 68104
rect 18115 68060 18173 68061
rect 3679 68020 3688 68060
rect 3728 68020 3770 68060
rect 3810 68020 3852 68060
rect 3892 68020 3934 68060
rect 3974 68020 4016 68060
rect 4056 68020 4065 68060
rect 6691 68020 6700 68060
rect 6740 68020 7468 68060
rect 7508 68020 7517 68060
rect 14563 68020 14572 68060
rect 14612 68020 16780 68060
rect 16820 68020 16829 68060
rect 18030 68020 18124 68060
rect 18164 68020 18173 68060
rect 18799 68020 18808 68060
rect 18848 68020 18890 68060
rect 18930 68020 18972 68060
rect 19012 68020 19054 68060
rect 19094 68020 19136 68060
rect 19176 68020 19185 68060
rect 18115 68019 18173 68020
rect 21424 67976 21504 67996
rect 7363 67936 7372 67976
rect 7412 67936 8716 67976
rect 8756 67936 10444 67976
rect 10484 67936 10493 67976
rect 10819 67936 10828 67976
rect 10868 67936 17260 67976
rect 17300 67936 17309 67976
rect 17923 67936 17932 67976
rect 17972 67936 19948 67976
rect 19988 67936 19997 67976
rect 20611 67936 20620 67976
rect 20660 67936 21504 67976
rect 21424 67916 21504 67936
rect 16579 67892 16637 67893
rect 6787 67852 6796 67892
rect 6836 67852 7948 67892
rect 7988 67852 7997 67892
rect 9091 67852 9100 67892
rect 9140 67852 9772 67892
rect 9812 67852 11360 67892
rect 15907 67852 15916 67892
rect 15956 67852 16588 67892
rect 16628 67852 16637 67892
rect 0 67808 80 67828
rect 11320 67808 11360 67852
rect 16579 67851 16637 67852
rect 0 67768 2092 67808
rect 2132 67768 2141 67808
rect 2947 67768 2956 67808
rect 2996 67768 3532 67808
rect 3572 67768 3581 67808
rect 6211 67768 6220 67808
rect 6260 67768 10060 67808
rect 10100 67768 10540 67808
rect 10580 67768 10589 67808
rect 11320 67768 11788 67808
rect 11828 67768 12748 67808
rect 12788 67768 12797 67808
rect 0 67748 80 67768
rect 7468 67684 9100 67724
rect 9140 67684 9149 67724
rect 9475 67684 9484 67724
rect 9524 67684 11252 67724
rect 15043 67684 15052 67724
rect 15092 67684 16972 67724
rect 17012 67684 17021 67724
rect 17251 67684 17260 67724
rect 17300 67684 18508 67724
rect 18548 67684 18557 67724
rect 7468 67640 7508 67684
rect 2467 67600 2476 67640
rect 2516 67600 2764 67640
rect 2804 67600 4204 67640
rect 4244 67600 4253 67640
rect 5827 67600 5836 67640
rect 5876 67600 7468 67640
rect 7508 67600 7517 67640
rect 7651 67600 7660 67640
rect 7700 67600 7709 67640
rect 8035 67600 8044 67640
rect 8084 67600 9772 67640
rect 9812 67600 10924 67640
rect 10964 67600 10973 67640
rect 5539 67556 5597 67557
rect 7660 67556 7700 67600
rect 11212 67556 11252 67684
rect 21424 67640 21504 67660
rect 12931 67600 12940 67640
rect 12980 67600 13420 67640
rect 13460 67600 14572 67640
rect 14612 67600 14621 67640
rect 14755 67600 14764 67640
rect 14804 67600 15724 67640
rect 15764 67600 15773 67640
rect 16300 67600 16588 67640
rect 16628 67600 17548 67640
rect 17588 67600 17597 67640
rect 19651 67600 19660 67640
rect 19700 67600 21504 67640
rect 16300 67556 16340 67600
rect 21424 67580 21504 67600
rect 18115 67556 18173 67557
rect 2947 67516 2956 67556
rect 2996 67516 5548 67556
rect 5588 67516 5597 67556
rect 5539 67515 5597 67516
rect 7468 67516 7700 67556
rect 11203 67516 11212 67556
rect 11252 67516 11261 67556
rect 16291 67516 16300 67556
rect 16340 67516 16349 67556
rect 16675 67516 16684 67556
rect 16724 67516 18124 67556
rect 18164 67516 18173 67556
rect 2563 67432 2572 67472
rect 2612 67432 3052 67472
rect 3092 67432 3101 67472
rect 6019 67432 6028 67472
rect 6068 67432 7372 67472
rect 7412 67432 7421 67472
rect 6595 67388 6653 67389
rect 7468 67388 7508 67516
rect 18115 67515 18173 67516
rect 20131 67432 20140 67472
rect 20180 67432 21332 67472
rect 14947 67388 15005 67389
rect 16963 67388 17021 67389
rect 1315 67348 1324 67388
rect 1364 67348 6604 67388
rect 6644 67348 6653 67388
rect 7459 67348 7468 67388
rect 7508 67348 7517 67388
rect 14947 67348 14956 67388
rect 14996 67348 16972 67388
rect 17012 67348 17260 67388
rect 17300 67348 17309 67388
rect 6595 67347 6653 67348
rect 14947 67347 15005 67348
rect 16963 67347 17021 67348
rect 21292 67304 21332 67432
rect 21424 67304 21504 67324
rect 4919 67264 4928 67304
rect 4968 67264 5010 67304
rect 5050 67264 5092 67304
rect 5132 67264 5174 67304
rect 5214 67264 5256 67304
rect 5296 67264 5305 67304
rect 14275 67264 14284 67304
rect 14324 67264 15916 67304
rect 15956 67264 15965 67304
rect 16387 67264 16396 67304
rect 16436 67264 16780 67304
rect 16820 67264 16829 67304
rect 20039 67264 20048 67304
rect 20088 67264 20130 67304
rect 20170 67264 20212 67304
rect 20252 67264 20294 67304
rect 20334 67264 20376 67304
rect 20416 67264 20425 67304
rect 21292 67264 21504 67304
rect 21424 67244 21504 67264
rect 15715 67180 15724 67220
rect 15764 67180 16876 67220
rect 16916 67180 16925 67220
rect 0 67136 80 67156
rect 1027 67136 1085 67137
rect 6307 67136 6365 67137
rect 0 67096 1036 67136
rect 1076 67096 1085 67136
rect 6211 67096 6220 67136
rect 6260 67096 6316 67136
rect 6356 67096 6365 67136
rect 14083 67096 14092 67136
rect 14132 67096 14476 67136
rect 14516 67096 14525 67136
rect 15235 67096 15244 67136
rect 15284 67096 19756 67136
rect 19796 67096 19805 67136
rect 0 67076 80 67096
rect 1027 67095 1085 67096
rect 6307 67095 6365 67096
rect 4387 67052 4445 67053
rect 4291 67012 4300 67052
rect 4340 67012 4396 67052
rect 4436 67012 4972 67052
rect 5012 67012 5021 67052
rect 11320 67012 16684 67052
rect 16724 67012 16733 67052
rect 4387 67011 4445 67012
rect 6115 66968 6173 66969
rect 1219 66928 1228 66968
rect 1268 66928 2284 66968
rect 2324 66928 2333 66968
rect 4579 66928 4588 66968
rect 4628 66928 5836 66968
rect 5876 66928 6124 66968
rect 6164 66928 6173 66968
rect 6115 66927 6173 66928
rect 6316 66928 8524 66968
rect 8564 66928 10156 66968
rect 10196 66928 10205 66968
rect 6316 66884 6356 66928
rect 8419 66884 8477 66885
rect 11320 66884 11360 67012
rect 21424 66968 21504 66988
rect 13027 66928 13036 66968
rect 13076 66928 14764 66968
rect 14804 66928 14813 66968
rect 16867 66928 16876 66968
rect 16916 66928 18508 66968
rect 18548 66928 18557 66968
rect 19939 66928 19948 66968
rect 19988 66928 21504 66968
rect 5347 66844 5356 66884
rect 5396 66844 6356 66884
rect 8334 66844 8428 66884
rect 8468 66844 11360 66884
rect 6316 66800 6356 66844
rect 8419 66843 8477 66844
rect 11779 66800 11837 66801
rect 4771 66760 4780 66800
rect 4820 66760 5836 66800
rect 5876 66760 5885 66800
rect 6316 66760 6452 66800
rect 2659 66676 2668 66716
rect 2708 66676 2956 66716
rect 2996 66676 3005 66716
rect 5731 66592 5740 66632
rect 5780 66592 6220 66632
rect 6260 66592 6269 66632
rect 6412 66548 6452 66760
rect 8140 66760 8716 66800
rect 8756 66760 8765 66800
rect 11779 66760 11788 66800
rect 11828 66760 12076 66800
rect 12116 66760 12125 66800
rect 8140 66632 8180 66760
rect 11779 66759 11837 66760
rect 13612 66632 13652 66928
rect 21424 66908 21504 66928
rect 14563 66844 14572 66884
rect 14612 66844 14956 66884
rect 14996 66844 15148 66884
rect 15188 66844 15197 66884
rect 15619 66844 15628 66884
rect 15668 66844 15820 66884
rect 15860 66844 15869 66884
rect 16579 66676 16588 66716
rect 16628 66676 17068 66716
rect 17108 66676 17117 66716
rect 21424 66632 21504 66652
rect 8131 66592 8140 66632
rect 8180 66592 8189 66632
rect 13603 66592 13612 66632
rect 13652 66592 13661 66632
rect 19459 66592 19468 66632
rect 19508 66592 21504 66632
rect 21424 66572 21504 66592
rect 3679 66508 3688 66548
rect 3728 66508 3770 66548
rect 3810 66508 3852 66548
rect 3892 66508 3934 66548
rect 3974 66508 4016 66548
rect 4056 66508 4065 66548
rect 6403 66508 6412 66548
rect 6452 66508 6461 66548
rect 18799 66508 18808 66548
rect 18848 66508 18890 66548
rect 18930 66508 18972 66548
rect 19012 66508 19054 66548
rect 19094 66508 19136 66548
rect 19176 66508 19185 66548
rect 0 66464 80 66484
rect 0 66424 76 66464
rect 116 66424 125 66464
rect 5635 66424 5644 66464
rect 5684 66424 6892 66464
rect 6932 66424 6941 66464
rect 10723 66424 10732 66464
rect 10772 66424 13036 66464
rect 13076 66424 13085 66464
rect 0 66404 80 66424
rect 3427 66340 3436 66380
rect 3476 66340 3724 66380
rect 3764 66340 3773 66380
rect 8515 66340 8524 66380
rect 8564 66340 10828 66380
rect 10868 66340 10877 66380
rect 13987 66340 13996 66380
rect 14036 66340 14188 66380
rect 14228 66340 14237 66380
rect 21424 66296 21504 66316
rect 2500 66256 3244 66296
rect 3284 66256 5740 66296
rect 5780 66256 19660 66296
rect 19700 66256 19709 66296
rect 19939 66256 19948 66296
rect 19988 66256 21504 66296
rect 2500 66128 2540 66256
rect 21424 66236 21504 66256
rect 4387 66172 4396 66212
rect 4436 66172 5164 66212
rect 5204 66172 5213 66212
rect 11491 66172 11500 66212
rect 11540 66172 19756 66212
rect 19796 66172 19805 66212
rect 17923 66128 17981 66129
rect 1411 66088 1420 66128
rect 1460 66088 2188 66128
rect 2228 66088 2540 66128
rect 2851 66088 2860 66128
rect 2900 66088 4300 66128
rect 4340 66088 4349 66128
rect 4579 66088 4588 66128
rect 4628 66088 6316 66128
rect 6356 66088 6365 66128
rect 9091 66088 9100 66128
rect 9140 66088 9388 66128
rect 9428 66088 9437 66128
rect 10339 66088 10348 66128
rect 10388 66088 11980 66128
rect 12020 66088 13612 66128
rect 13652 66088 13661 66128
rect 16675 66088 16684 66128
rect 16724 66088 17356 66128
rect 17396 66088 17548 66128
rect 17588 66088 17597 66128
rect 17838 66088 17932 66128
rect 17972 66088 17981 66128
rect 17923 66087 17981 66088
rect 4099 66044 4157 66045
rect 3235 66004 3244 66044
rect 3284 66004 4108 66044
rect 4148 66004 4780 66044
rect 4820 66004 4829 66044
rect 4099 66003 4157 66004
rect 16963 65960 17021 65961
rect 16867 65920 16876 65960
rect 16916 65920 16972 65960
rect 17012 65920 17021 65960
rect 16963 65919 17021 65920
rect 18019 65960 18077 65961
rect 21424 65960 21504 65980
rect 18019 65920 18028 65960
rect 18068 65920 19180 65960
rect 19220 65920 19229 65960
rect 19555 65920 19564 65960
rect 19604 65920 21504 65960
rect 18019 65919 18077 65920
rect 21424 65900 21504 65920
rect 0 65792 80 65812
rect 1219 65792 1277 65793
rect 0 65752 1228 65792
rect 1268 65752 1277 65792
rect 4919 65752 4928 65792
rect 4968 65752 5010 65792
rect 5050 65752 5092 65792
rect 5132 65752 5174 65792
rect 5214 65752 5256 65792
rect 5296 65752 5305 65792
rect 20039 65752 20048 65792
rect 20088 65752 20130 65792
rect 20170 65752 20212 65792
rect 20252 65752 20294 65792
rect 20334 65752 20376 65792
rect 20416 65752 20425 65792
rect 0 65732 80 65752
rect 1219 65751 1277 65752
rect 3907 65668 3916 65708
rect 3956 65668 10444 65708
rect 10484 65668 10493 65708
rect 12259 65668 12268 65708
rect 12308 65668 12556 65708
rect 12596 65668 12605 65708
rect 18115 65668 18124 65708
rect 18164 65668 18173 65708
rect 13219 65624 13277 65625
rect 2851 65584 2860 65624
rect 2900 65584 3188 65624
rect 3619 65584 3628 65624
rect 3668 65584 4204 65624
rect 4244 65584 4253 65624
rect 5443 65584 5452 65624
rect 5492 65584 5932 65624
rect 5972 65584 5981 65624
rect 9475 65584 9484 65624
rect 9524 65584 13228 65624
rect 13268 65584 13277 65624
rect 16291 65584 16300 65624
rect 16340 65584 16684 65624
rect 16724 65584 16733 65624
rect 17635 65584 17644 65624
rect 17684 65584 17932 65624
rect 17972 65584 17981 65624
rect 3148 65540 3188 65584
rect 13219 65583 13277 65584
rect 8515 65540 8573 65541
rect 18124 65540 18164 65668
rect 21424 65624 21504 65644
rect 19939 65584 19948 65624
rect 19988 65584 21504 65624
rect 21424 65564 21504 65584
rect 835 65500 844 65540
rect 884 65500 1804 65540
rect 1844 65500 1853 65540
rect 3139 65500 3148 65540
rect 3188 65500 3197 65540
rect 3811 65500 3820 65540
rect 3860 65500 4684 65540
rect 4724 65500 4733 65540
rect 5347 65500 5356 65540
rect 5396 65500 8524 65540
rect 8564 65500 8573 65540
rect 10243 65500 10252 65540
rect 10292 65500 11116 65540
rect 11156 65500 11308 65540
rect 11348 65500 11357 65540
rect 12931 65500 12940 65540
rect 12980 65500 13900 65540
rect 13940 65500 13949 65540
rect 17731 65500 17740 65540
rect 17780 65500 18164 65540
rect 18307 65500 18316 65540
rect 18356 65500 19372 65540
rect 19412 65500 19421 65540
rect 8515 65499 8573 65500
rect 2755 65456 2813 65457
rect 11395 65456 11453 65457
rect 17923 65456 17981 65457
rect 2755 65416 2764 65456
rect 2804 65416 2860 65456
rect 2900 65416 3724 65456
rect 3764 65416 3773 65456
rect 4387 65416 4396 65456
rect 4436 65416 5396 65456
rect 5443 65416 5452 65456
rect 5492 65416 6124 65456
rect 6164 65416 7084 65456
rect 7124 65416 7133 65456
rect 11310 65416 11404 65456
rect 11444 65416 11453 65456
rect 13795 65416 13804 65456
rect 13844 65416 15532 65456
rect 15572 65416 15581 65456
rect 17059 65416 17068 65456
rect 17108 65416 17932 65456
rect 17972 65416 17981 65456
rect 18115 65416 18124 65456
rect 18164 65416 18700 65456
rect 18740 65416 18749 65456
rect 2755 65415 2813 65416
rect 5356 65372 5396 65416
rect 11395 65415 11453 65416
rect 17923 65415 17981 65416
rect 10531 65372 10589 65373
rect 5356 65332 9100 65372
rect 9140 65332 10540 65372
rect 10580 65332 10589 65372
rect 15427 65332 15436 65372
rect 15476 65332 19756 65372
rect 19796 65332 19805 65372
rect 10531 65331 10589 65332
rect 4291 65288 4349 65289
rect 21424 65288 21504 65308
rect 4206 65248 4300 65288
rect 4340 65248 4349 65288
rect 4483 65248 4492 65288
rect 4532 65248 6892 65288
rect 6932 65248 10348 65288
rect 10388 65248 10397 65288
rect 12643 65248 12652 65288
rect 12692 65248 18988 65288
rect 19028 65248 19037 65288
rect 20035 65248 20044 65288
rect 20084 65248 21504 65288
rect 4291 65247 4349 65248
rect 21424 65228 21504 65248
rect 6115 65204 6173 65205
rect 6030 65164 6124 65204
rect 6164 65164 6173 65204
rect 10531 65164 10540 65204
rect 10580 65164 11308 65204
rect 11348 65164 11357 65204
rect 6115 65163 6173 65164
rect 0 65120 80 65140
rect 0 65080 748 65120
rect 788 65080 797 65120
rect 3139 65080 3148 65120
rect 3188 65080 3436 65120
rect 3476 65080 3485 65120
rect 0 65060 80 65080
rect 3679 64996 3688 65036
rect 3728 64996 3770 65036
rect 3810 64996 3852 65036
rect 3892 64996 3934 65036
rect 3974 64996 4016 65036
rect 4056 64996 4065 65036
rect 18799 64996 18808 65036
rect 18848 64996 18890 65036
rect 18930 64996 18972 65036
rect 19012 64996 19054 65036
rect 19094 64996 19136 65036
rect 19176 64996 19185 65036
rect 21424 64952 21504 64972
rect 19267 64912 19276 64952
rect 19316 64912 21504 64952
rect 21424 64892 21504 64912
rect 10531 64868 10589 64869
rect 10531 64828 10540 64868
rect 10580 64828 19852 64868
rect 19892 64828 19901 64868
rect 10531 64827 10589 64828
rect 2659 64744 2668 64784
rect 2708 64744 3148 64784
rect 3188 64744 3820 64784
rect 3860 64744 3869 64784
rect 7075 64660 7084 64700
rect 7124 64660 8524 64700
rect 8564 64660 8716 64700
rect 8756 64660 8765 64700
rect 11011 64660 11020 64700
rect 11060 64660 17740 64700
rect 17780 64660 17789 64700
rect 13795 64616 13853 64617
rect 14851 64616 14909 64617
rect 21424 64616 21504 64636
rect 2563 64576 2572 64616
rect 2612 64576 4396 64616
rect 4436 64576 4445 64616
rect 7267 64576 7276 64616
rect 7316 64576 9772 64616
rect 9812 64576 9821 64616
rect 10819 64576 10828 64616
rect 10868 64576 10877 64616
rect 13795 64576 13804 64616
rect 13844 64576 13996 64616
rect 14036 64576 14860 64616
rect 14900 64576 14909 64616
rect 15715 64576 15724 64616
rect 15764 64576 16300 64616
rect 16340 64576 16349 64616
rect 16675 64576 16684 64616
rect 16724 64576 17068 64616
rect 17108 64576 17117 64616
rect 19555 64576 19564 64616
rect 19604 64576 21504 64616
rect 10828 64532 10868 64576
rect 13795 64575 13853 64576
rect 14851 64575 14909 64576
rect 21424 64556 21504 64576
rect 5635 64492 5644 64532
rect 5684 64492 7564 64532
rect 7604 64492 7613 64532
rect 8611 64492 8620 64532
rect 8660 64492 10868 64532
rect 16963 64492 16972 64532
rect 17012 64492 18988 64532
rect 19028 64492 19660 64532
rect 19700 64492 19709 64532
rect 0 64448 80 64468
rect 0 64408 1132 64448
rect 1172 64408 1181 64448
rect 7267 64408 7276 64448
rect 7316 64408 7948 64448
rect 7988 64408 7997 64448
rect 9283 64408 9292 64448
rect 9332 64408 19756 64448
rect 19796 64408 19805 64448
rect 0 64388 80 64408
rect 2947 64364 3005 64365
rect 2947 64324 2956 64364
rect 2996 64324 4492 64364
rect 4532 64324 4541 64364
rect 6883 64324 6892 64364
rect 6932 64324 8044 64364
rect 8084 64324 8093 64364
rect 9955 64324 9964 64364
rect 10004 64324 11212 64364
rect 11252 64324 11261 64364
rect 14275 64324 14284 64364
rect 14324 64324 18124 64364
rect 18164 64324 18173 64364
rect 19948 64324 20564 64364
rect 2947 64323 3005 64324
rect 3043 64280 3101 64281
rect 7651 64280 7709 64281
rect 19948 64280 19988 64324
rect 20524 64280 20564 64324
rect 21424 64280 21504 64300
rect 3043 64240 3052 64280
rect 3092 64240 3244 64280
rect 3284 64240 3293 64280
rect 4919 64240 4928 64280
rect 4968 64240 5010 64280
rect 5050 64240 5092 64280
rect 5132 64240 5174 64280
rect 5214 64240 5256 64280
rect 5296 64240 5305 64280
rect 7566 64240 7660 64280
rect 7700 64240 7709 64280
rect 3043 64239 3101 64240
rect 7651 64239 7709 64240
rect 14956 64240 15148 64280
rect 15188 64240 15197 64280
rect 19908 64240 19948 64280
rect 19988 64240 19997 64280
rect 20039 64240 20048 64280
rect 20088 64240 20130 64280
rect 20170 64240 20212 64280
rect 20252 64240 20294 64280
rect 20334 64240 20376 64280
rect 20416 64240 20425 64280
rect 20524 64240 21504 64280
rect 14956 64196 14996 64240
rect 21424 64220 21504 64240
rect 4003 64156 4012 64196
rect 4052 64156 6796 64196
rect 6836 64156 6845 64196
rect 13603 64156 13612 64196
rect 13652 64156 14996 64196
rect 18019 64156 18028 64196
rect 18068 64156 18604 64196
rect 18644 64156 18653 64196
rect 1699 64072 1708 64112
rect 1748 64072 2764 64112
rect 2804 64072 3532 64112
rect 3572 64072 3581 64112
rect 4099 64072 4108 64112
rect 4148 64072 4972 64112
rect 5012 64072 5021 64112
rect 7267 64072 7276 64112
rect 7316 64072 7468 64112
rect 7508 64072 7517 64112
rect 8515 64072 8524 64112
rect 8564 64072 19468 64112
rect 19508 64072 19517 64112
rect 8515 64028 8573 64029
rect 5155 63988 5164 64028
rect 5204 63988 5740 64028
rect 5780 63988 5789 64028
rect 8323 63988 8332 64028
rect 8372 63988 8524 64028
rect 8564 63988 8573 64028
rect 11011 63988 11020 64028
rect 11060 63988 12404 64028
rect 12643 63988 12652 64028
rect 12692 63988 19372 64028
rect 19412 63988 19421 64028
rect 8515 63987 8573 63988
rect 4195 63944 4253 63945
rect 8995 63944 9053 63945
rect 12364 63944 12404 63988
rect 21424 63944 21504 63964
rect 2947 63904 2956 63944
rect 2996 63904 3148 63944
rect 3188 63904 4204 63944
rect 4244 63904 4253 63944
rect 7459 63904 7468 63944
rect 7508 63904 9004 63944
rect 9044 63904 11788 63944
rect 11828 63904 11837 63944
rect 12355 63904 12364 63944
rect 12404 63904 12413 63944
rect 13315 63904 13324 63944
rect 13364 63904 13996 63944
rect 14036 63904 14668 63944
rect 14708 63904 14717 63944
rect 14947 63904 14956 63944
rect 14996 63904 18508 63944
rect 18548 63904 18557 63944
rect 19555 63904 19564 63944
rect 19604 63904 21504 63944
rect 4195 63903 4253 63904
rect 8995 63903 9053 63904
rect 21424 63884 21504 63904
rect 11299 63860 11357 63861
rect 15043 63860 15101 63861
rect 3436 63820 4012 63860
rect 4052 63820 4061 63860
rect 6211 63820 6220 63860
rect 6260 63820 6988 63860
rect 7028 63820 7037 63860
rect 8131 63820 8140 63860
rect 8180 63820 8524 63860
rect 8564 63820 8573 63860
rect 10051 63820 10060 63860
rect 10100 63820 10348 63860
rect 10388 63820 10397 63860
rect 11214 63820 11308 63860
rect 11348 63820 11357 63860
rect 14371 63820 14380 63860
rect 14420 63820 14860 63860
rect 14900 63820 15052 63860
rect 15092 63820 15101 63860
rect 15619 63820 15628 63860
rect 15668 63820 19756 63860
rect 19796 63820 19805 63860
rect 0 63776 80 63796
rect 3436 63776 3476 63820
rect 11299 63819 11357 63820
rect 15043 63819 15101 63820
rect 17923 63776 17981 63777
rect 18499 63776 18557 63777
rect 0 63736 2540 63776
rect 3427 63736 3436 63776
rect 3476 63736 3485 63776
rect 3907 63736 3916 63776
rect 3956 63736 4204 63776
rect 4244 63736 6028 63776
rect 6068 63736 6077 63776
rect 10531 63736 10540 63776
rect 10580 63736 11020 63776
rect 11060 63736 11069 63776
rect 17838 63736 17932 63776
rect 17972 63736 18508 63776
rect 18548 63736 18557 63776
rect 0 63716 80 63736
rect 2500 63608 2540 63736
rect 17923 63735 17981 63736
rect 18499 63735 18557 63736
rect 5539 63692 5597 63693
rect 3139 63652 3148 63692
rect 3188 63652 4396 63692
rect 4436 63652 4445 63692
rect 5539 63652 5548 63692
rect 5588 63652 9100 63692
rect 9140 63652 9149 63692
rect 10435 63652 10444 63692
rect 10484 63652 10828 63692
rect 10868 63652 10877 63692
rect 5539 63651 5597 63652
rect 21424 63608 21504 63628
rect 2500 63568 13420 63608
rect 13460 63568 13469 63608
rect 19939 63568 19948 63608
rect 19988 63568 21504 63608
rect 21424 63548 21504 63568
rect 3679 63484 3688 63524
rect 3728 63484 3770 63524
rect 3810 63484 3852 63524
rect 3892 63484 3934 63524
rect 3974 63484 4016 63524
rect 4056 63484 4065 63524
rect 8419 63484 8428 63524
rect 8468 63484 10636 63524
rect 10676 63484 10685 63524
rect 18799 63484 18808 63524
rect 18848 63484 18890 63524
rect 18930 63484 18972 63524
rect 19012 63484 19054 63524
rect 19094 63484 19136 63524
rect 19176 63484 19185 63524
rect 3139 63400 3148 63440
rect 3188 63400 3532 63440
rect 3572 63400 3581 63440
rect 10051 63400 10060 63440
rect 10100 63400 11884 63440
rect 11924 63400 11933 63440
rect 5539 63356 5597 63357
rect 3907 63316 3916 63356
rect 3956 63316 4492 63356
rect 4532 63316 4541 63356
rect 5347 63316 5356 63356
rect 5396 63316 5548 63356
rect 5588 63316 5597 63356
rect 5539 63315 5597 63316
rect 5827 63356 5885 63357
rect 5827 63316 5836 63356
rect 5876 63316 11360 63356
rect 5827 63315 5885 63316
rect 11320 63272 11360 63316
rect 17260 63316 18028 63356
rect 18068 63316 18077 63356
rect 17260 63272 17300 63316
rect 21424 63272 21504 63292
rect 3331 63232 3340 63272
rect 3380 63232 3532 63272
rect 3572 63232 3581 63272
rect 4579 63232 4588 63272
rect 4628 63232 6604 63272
rect 6644 63232 6653 63272
rect 8803 63232 8812 63272
rect 8852 63232 9100 63272
rect 9140 63232 9149 63272
rect 11320 63232 12748 63272
rect 12788 63232 12797 63272
rect 14467 63232 14476 63272
rect 14516 63232 17260 63272
rect 17300 63232 17309 63272
rect 17635 63232 17644 63272
rect 17684 63232 17693 63272
rect 19651 63232 19660 63272
rect 19700 63232 21504 63272
rect 8995 63188 9053 63189
rect 2500 63148 7700 63188
rect 8910 63148 9004 63188
rect 9044 63148 9053 63188
rect 10531 63148 10540 63188
rect 10580 63148 10732 63188
rect 10772 63148 10781 63188
rect 16963 63148 16972 63188
rect 17012 63148 17021 63188
rect 0 63104 80 63124
rect 2500 63104 2540 63148
rect 5539 63104 5597 63105
rect 6595 63104 6653 63105
rect 0 63064 2540 63104
rect 2947 63064 2956 63104
rect 2996 63064 3148 63104
rect 3188 63064 3197 63104
rect 3331 63064 3340 63104
rect 3380 63064 4204 63104
rect 4244 63064 4253 63104
rect 5539 63064 5548 63104
rect 5588 63064 5644 63104
rect 5684 63064 5693 63104
rect 6595 63064 6604 63104
rect 6644 63064 7372 63104
rect 7412 63064 7421 63104
rect 0 63044 80 63064
rect 5539 63063 5597 63064
rect 6595 63063 6653 63064
rect 7660 63020 7700 63148
rect 8995 63147 9053 63148
rect 16099 63104 16157 63105
rect 8611 63064 8620 63104
rect 8660 63064 10060 63104
rect 10100 63064 10252 63104
rect 10292 63064 10301 63104
rect 12739 63064 12748 63104
rect 12788 63064 13804 63104
rect 13844 63064 13853 63104
rect 15139 63064 15148 63104
rect 15188 63064 15532 63104
rect 15572 63064 16108 63104
rect 16148 63064 16157 63104
rect 16099 63063 16157 63064
rect 16972 63020 17012 63148
rect 17155 63064 17164 63104
rect 17204 63064 17548 63104
rect 17588 63064 17597 63104
rect 4675 62980 4684 63020
rect 4724 62980 6220 63020
rect 6260 62980 6269 63020
rect 7075 62980 7084 63020
rect 7124 62980 7564 63020
rect 7604 62980 7613 63020
rect 7660 62980 10732 63020
rect 10772 62980 10781 63020
rect 13699 62980 13708 63020
rect 13748 62980 15052 63020
rect 15092 62980 16780 63020
rect 16820 62980 17012 63020
rect 17644 63020 17684 63232
rect 21424 63212 21504 63232
rect 18115 63104 18173 63105
rect 18019 63064 18028 63104
rect 18068 63064 18124 63104
rect 18164 63064 18173 63104
rect 18115 63063 18173 63064
rect 17644 62980 18508 63020
rect 18548 62980 18557 63020
rect 21424 62936 21504 62956
rect 5443 62896 5452 62936
rect 5492 62896 5932 62936
rect 5972 62896 10924 62936
rect 10964 62896 10973 62936
rect 17155 62896 17164 62936
rect 17204 62896 17644 62936
rect 17684 62896 17693 62936
rect 20515 62896 20524 62936
rect 20564 62896 21504 62936
rect 21424 62876 21504 62896
rect 13795 62852 13853 62853
rect 1699 62812 1708 62852
rect 1748 62812 6356 62852
rect 13603 62812 13612 62852
rect 13652 62812 13804 62852
rect 13844 62812 13853 62852
rect 6316 62769 6356 62812
rect 13795 62811 13853 62812
rect 14083 62852 14141 62853
rect 14083 62812 14092 62852
rect 14132 62812 15052 62852
rect 15092 62812 15101 62852
rect 14083 62811 14141 62812
rect 6307 62768 6365 62769
rect 2563 62728 2572 62768
rect 2612 62728 3052 62768
rect 3092 62728 3101 62768
rect 4919 62728 4928 62768
rect 4968 62728 5010 62768
rect 5050 62728 5092 62768
rect 5132 62728 5174 62768
rect 5214 62728 5256 62768
rect 5296 62728 5305 62768
rect 6307 62728 6316 62768
rect 6356 62728 8812 62768
rect 8852 62728 8861 62768
rect 20039 62728 20048 62768
rect 20088 62728 20130 62768
rect 20170 62728 20212 62768
rect 20252 62728 20294 62768
rect 20334 62728 20376 62768
rect 20416 62728 20425 62768
rect 6307 62727 6365 62728
rect 1987 62644 1996 62684
rect 2036 62644 2540 62684
rect 9283 62644 9292 62684
rect 9332 62644 19660 62684
rect 19700 62644 19709 62684
rect 2500 62600 2540 62644
rect 14467 62600 14525 62601
rect 21424 62600 21504 62620
rect 2500 62560 14476 62600
rect 14516 62560 14525 62600
rect 16483 62560 16492 62600
rect 16532 62560 16780 62600
rect 16820 62560 16829 62600
rect 19843 62560 19852 62600
rect 19892 62560 21504 62600
rect 14467 62559 14525 62560
rect 21424 62540 21504 62560
rect 8323 62516 8381 62517
rect 2956 62476 7948 62516
rect 7988 62476 8332 62516
rect 8372 62476 8381 62516
rect 0 62432 80 62452
rect 1699 62432 1757 62433
rect 2956 62432 2996 62476
rect 8323 62475 8381 62476
rect 4195 62432 4253 62433
rect 7651 62432 7709 62433
rect 0 62392 1708 62432
rect 1748 62392 1757 62432
rect 2947 62392 2956 62432
rect 2996 62392 3005 62432
rect 4110 62392 4204 62432
rect 4244 62392 4253 62432
rect 7566 62392 7660 62432
rect 7700 62392 7709 62432
rect 8227 62392 8236 62432
rect 8276 62392 8620 62432
rect 8660 62392 8669 62432
rect 17731 62392 17740 62432
rect 17780 62392 18028 62432
rect 18068 62392 18077 62432
rect 0 62372 80 62392
rect 1699 62391 1757 62392
rect 4195 62391 4253 62392
rect 7651 62391 7709 62392
rect 4204 62348 4244 62391
rect 1315 62308 1324 62348
rect 1364 62308 1708 62348
rect 1748 62308 1757 62348
rect 2476 62308 4244 62348
rect 6787 62308 6796 62348
rect 6836 62308 7468 62348
rect 7508 62308 8044 62348
rect 8084 62308 8093 62348
rect 15619 62308 15628 62348
rect 15668 62308 20044 62348
rect 20084 62308 20093 62348
rect 2476 62264 2516 62308
rect 21424 62264 21504 62284
rect 2467 62224 2476 62264
rect 2516 62224 2525 62264
rect 14755 62224 14764 62264
rect 14804 62224 14956 62264
rect 14996 62224 18508 62264
rect 18548 62224 18557 62264
rect 18691 62224 18700 62264
rect 18740 62224 21504 62264
rect 21424 62204 21504 62224
rect 11203 62096 11261 62097
rect 7555 62056 7564 62096
rect 7604 62056 11212 62096
rect 11252 62056 11261 62096
rect 11203 62055 11261 62056
rect 3679 61972 3688 62012
rect 3728 61972 3770 62012
rect 3810 61972 3852 62012
rect 3892 61972 3934 62012
rect 3974 61972 4016 62012
rect 4056 61972 4065 62012
rect 6211 61972 6220 62012
rect 6260 61972 6508 62012
rect 6548 61972 6557 62012
rect 18799 61972 18808 62012
rect 18848 61972 18890 62012
rect 18930 61972 18972 62012
rect 19012 61972 19054 62012
rect 19094 61972 19136 62012
rect 19176 61972 19185 62012
rect 16099 61928 16157 61929
rect 21424 61928 21504 61948
rect 1603 61888 1612 61928
rect 1652 61888 8044 61928
rect 8084 61888 8093 61928
rect 16099 61888 16108 61928
rect 16148 61888 16300 61928
rect 16340 61888 16349 61928
rect 19939 61888 19948 61928
rect 19988 61888 21504 61928
rect 16099 61887 16157 61888
rect 21424 61868 21504 61888
rect 11971 61844 12029 61845
rect 17155 61844 17213 61845
rect 2500 61804 10444 61844
rect 10484 61804 10493 61844
rect 11107 61804 11116 61844
rect 11156 61804 11404 61844
rect 11444 61804 11453 61844
rect 11971 61804 11980 61844
rect 12020 61804 17164 61844
rect 17204 61804 17213 61844
rect 18595 61804 18604 61844
rect 18644 61804 18653 61844
rect 0 61760 80 61780
rect 2500 61760 2540 61804
rect 11971 61803 12029 61804
rect 17155 61803 17213 61804
rect 2755 61760 2813 61761
rect 7555 61760 7613 61761
rect 9763 61760 9821 61761
rect 15619 61760 15677 61761
rect 0 61720 2540 61760
rect 2670 61720 2764 61760
rect 2804 61720 2813 61760
rect 4387 61720 4396 61760
rect 4436 61720 4684 61760
rect 4724 61720 4733 61760
rect 6403 61720 6412 61760
rect 6452 61720 6700 61760
rect 6740 61720 6749 61760
rect 7171 61720 7180 61760
rect 7220 61720 7564 61760
rect 7604 61720 7613 61760
rect 8899 61720 8908 61760
rect 8948 61720 9484 61760
rect 9524 61720 9533 61760
rect 9678 61720 9772 61760
rect 9812 61720 9821 61760
rect 10243 61720 10252 61760
rect 10292 61720 10540 61760
rect 10580 61720 10589 61760
rect 11683 61720 11692 61760
rect 11732 61720 13324 61760
rect 13364 61720 13373 61760
rect 14083 61720 14092 61760
rect 14132 61720 14572 61760
rect 14612 61720 14621 61760
rect 15534 61720 15628 61760
rect 15668 61720 15677 61760
rect 18604 61760 18644 61804
rect 18604 61720 19084 61760
rect 19124 61720 19133 61760
rect 0 61700 80 61720
rect 2755 61719 2813 61720
rect 7555 61719 7613 61720
rect 9763 61719 9821 61720
rect 15619 61719 15677 61720
rect 8995 61676 9053 61677
rect 3427 61636 3436 61676
rect 3476 61636 3724 61676
rect 3764 61636 3773 61676
rect 7651 61636 7660 61676
rect 7700 61636 9004 61676
rect 9044 61636 9053 61676
rect 10339 61636 10348 61676
rect 10388 61636 10484 61676
rect 12259 61636 12268 61676
rect 12308 61636 18604 61676
rect 18644 61636 18653 61676
rect 8995 61635 9053 61636
rect 10444 61593 10484 61636
rect 3331 61592 3389 61593
rect 10435 61592 10493 61593
rect 18307 61592 18365 61593
rect 21424 61592 21504 61612
rect 2659 61552 2668 61592
rect 2708 61552 2860 61592
rect 2900 61552 2909 61592
rect 3246 61552 3340 61592
rect 3380 61552 3389 61592
rect 5347 61552 5356 61592
rect 5396 61552 5644 61592
rect 5684 61552 5693 61592
rect 5923 61552 5932 61592
rect 5972 61552 6604 61592
rect 6644 61552 8428 61592
rect 8468 61552 9964 61592
rect 10004 61552 10013 61592
rect 10435 61552 10444 61592
rect 10484 61552 11020 61592
rect 11060 61552 11069 61592
rect 14083 61552 14092 61592
rect 14132 61552 16204 61592
rect 16244 61552 18316 61592
rect 18356 61552 18365 61592
rect 19171 61552 19180 61592
rect 19220 61552 21504 61592
rect 3331 61551 3389 61552
rect 10435 61551 10493 61552
rect 18307 61551 18365 61552
rect 21424 61532 21504 61552
rect 12451 61508 12509 61509
rect 16291 61508 16349 61509
rect 1507 61468 1516 61508
rect 1556 61468 7084 61508
rect 7124 61468 7660 61508
rect 7700 61468 7709 61508
rect 12366 61468 12460 61508
rect 12500 61468 16300 61508
rect 16340 61468 16349 61508
rect 12451 61467 12509 61468
rect 16291 61467 16349 61468
rect 10915 61424 10973 61425
rect 16675 61424 16733 61425
rect 3043 61384 3052 61424
rect 3092 61384 3436 61424
rect 3476 61384 3485 61424
rect 6787 61384 6796 61424
rect 6836 61384 7220 61424
rect 8035 61384 8044 61424
rect 8084 61384 8428 61424
rect 8468 61384 8477 61424
rect 10915 61384 10924 61424
rect 10964 61384 11500 61424
rect 11540 61384 14572 61424
rect 14612 61384 16684 61424
rect 16724 61384 16733 61424
rect 19555 61384 19564 61424
rect 19604 61384 21332 61424
rect 7180 61340 7220 61384
rect 10915 61383 10973 61384
rect 16675 61383 16733 61384
rect 7171 61300 7180 61340
rect 7220 61300 7229 61340
rect 10243 61300 10252 61340
rect 10292 61300 10540 61340
rect 10580 61300 10589 61340
rect 12163 61300 12172 61340
rect 12212 61300 15820 61340
rect 15860 61300 16588 61340
rect 16628 61300 17452 61340
rect 17492 61300 17501 61340
rect 14572 61256 14612 61300
rect 21292 61256 21332 61384
rect 21424 61256 21504 61276
rect 4919 61216 4928 61256
rect 4968 61216 5010 61256
rect 5050 61216 5092 61256
rect 5132 61216 5174 61256
rect 5214 61216 5256 61256
rect 5296 61216 5305 61256
rect 13027 61216 13036 61256
rect 13076 61216 13900 61256
rect 13940 61216 13949 61256
rect 14563 61216 14572 61256
rect 14612 61216 14621 61256
rect 20039 61216 20048 61256
rect 20088 61216 20130 61256
rect 20170 61216 20212 61256
rect 20252 61216 20294 61256
rect 20334 61216 20376 61256
rect 20416 61216 20425 61256
rect 21292 61216 21504 61256
rect 21424 61196 21504 61216
rect 1891 61132 1900 61172
rect 1940 61132 9772 61172
rect 9812 61132 9821 61172
rect 12451 61132 12460 61172
rect 12500 61132 19372 61172
rect 19412 61132 19421 61172
rect 0 61088 80 61108
rect 1123 61088 1181 61089
rect 11683 61088 11741 61089
rect 0 61048 1132 61088
rect 1172 61048 1181 61088
rect 2851 61048 2860 61088
rect 2900 61048 4396 61088
rect 4436 61048 4445 61088
rect 5443 61048 5452 61088
rect 5492 61048 7276 61088
rect 7316 61048 7325 61088
rect 10531 61048 10540 61088
rect 10580 61048 10828 61088
rect 10868 61048 10877 61088
rect 11683 61048 11692 61088
rect 11732 61048 15148 61088
rect 15188 61048 15197 61088
rect 17827 61048 17836 61088
rect 17876 61048 18988 61088
rect 19028 61048 19037 61088
rect 0 61028 80 61048
rect 1123 61047 1181 61048
rect 11683 61047 11741 61048
rect 13795 61004 13853 61005
rect 259 60964 268 61004
rect 308 60964 13804 61004
rect 13844 60964 13853 61004
rect 13795 60963 13853 60964
rect 2467 60920 2525 60921
rect 15619 60920 15677 60921
rect 21424 60920 21504 60940
rect 2467 60880 2476 60920
rect 2516 60880 2572 60920
rect 2612 60880 2621 60920
rect 2668 60880 3148 60920
rect 3188 60880 3197 60920
rect 6211 60880 6220 60920
rect 6260 60880 7276 60920
rect 7316 60880 10004 60920
rect 10051 60880 10060 60920
rect 10100 60880 15628 60920
rect 15668 60880 15677 60920
rect 19459 60880 19468 60920
rect 19508 60880 21504 60920
rect 2467 60879 2525 60880
rect 1603 60796 1612 60836
rect 1652 60796 2284 60836
rect 2324 60796 2540 60836
rect 2500 60668 2540 60796
rect 2668 60752 2708 60880
rect 9187 60836 9245 60837
rect 2956 60796 5452 60836
rect 5492 60796 5501 60836
rect 6499 60796 6508 60836
rect 6548 60796 6988 60836
rect 7028 60796 7660 60836
rect 7700 60796 7709 60836
rect 8995 60796 9004 60836
rect 9044 60796 9196 60836
rect 9236 60796 9245 60836
rect 9964 60836 10004 60880
rect 15619 60879 15677 60880
rect 21424 60860 21504 60880
rect 11203 60836 11261 60837
rect 9964 60796 10540 60836
rect 10580 60796 10589 60836
rect 11118 60796 11212 60836
rect 11252 60796 11261 60836
rect 14947 60796 14956 60836
rect 14996 60796 20044 60836
rect 20084 60796 20093 60836
rect 2659 60712 2668 60752
rect 2708 60712 2717 60752
rect 2956 60668 2996 60796
rect 9187 60795 9245 60796
rect 3331 60752 3389 60753
rect 3331 60712 3340 60752
rect 3380 60712 3628 60752
rect 3668 60712 3677 60752
rect 5827 60712 5836 60752
rect 5876 60712 6700 60752
rect 6740 60712 9044 60752
rect 3331 60711 3389 60712
rect 9004 60668 9044 60712
rect 10540 60668 10580 60796
rect 11203 60795 11261 60796
rect 14371 60752 14429 60753
rect 18499 60752 18557 60753
rect 10819 60712 10828 60752
rect 10868 60712 11308 60752
rect 11348 60712 11357 60752
rect 14371 60712 14380 60752
rect 14420 60712 14860 60752
rect 14900 60712 16588 60752
rect 16628 60712 16637 60752
rect 18499 60712 18508 60752
rect 18548 60712 18604 60752
rect 18644 60712 18653 60752
rect 14371 60711 14429 60712
rect 18499 60711 18557 60712
rect 19363 60668 19421 60669
rect 2500 60628 2996 60668
rect 3715 60628 3724 60668
rect 3764 60628 4108 60668
rect 4148 60628 4157 60668
rect 6883 60628 6892 60668
rect 6932 60628 7660 60668
rect 7700 60628 7709 60668
rect 8995 60628 9004 60668
rect 9044 60628 9053 60668
rect 10540 60628 12172 60668
rect 12212 60628 12221 60668
rect 17155 60628 17164 60668
rect 17204 60628 19180 60668
rect 19220 60628 19372 60668
rect 19412 60628 19421 60668
rect 19363 60627 19421 60628
rect 21424 60584 21504 60604
rect 1411 60544 1420 60584
rect 1460 60544 1996 60584
rect 2036 60544 8524 60584
rect 8564 60544 8573 60584
rect 10339 60544 10348 60584
rect 10388 60544 14668 60584
rect 14708 60544 16204 60584
rect 16244 60544 16253 60584
rect 16675 60544 16684 60584
rect 16724 60544 17260 60584
rect 17300 60544 18604 60584
rect 18644 60544 18653 60584
rect 20995 60544 21004 60584
rect 21044 60544 21504 60584
rect 21424 60524 21504 60544
rect 6787 60500 6845 60501
rect 3679 60460 3688 60500
rect 3728 60460 3770 60500
rect 3810 60460 3852 60500
rect 3892 60460 3934 60500
rect 3974 60460 4016 60500
rect 4056 60460 4065 60500
rect 4771 60460 4780 60500
rect 4820 60460 6796 60500
rect 6836 60460 6845 60500
rect 10627 60460 10636 60500
rect 10676 60460 11360 60500
rect 12451 60460 12460 60500
rect 12500 60460 13324 60500
rect 13364 60460 13373 60500
rect 14275 60460 14284 60500
rect 14324 60460 17356 60500
rect 17396 60460 18220 60500
rect 18260 60460 18269 60500
rect 18799 60460 18808 60500
rect 18848 60460 18890 60500
rect 18930 60460 18972 60500
rect 19012 60460 19054 60500
rect 19094 60460 19136 60500
rect 19176 60460 19185 60500
rect 6787 60459 6845 60460
rect 0 60416 80 60436
rect 11320 60416 11360 60460
rect 0 60376 940 60416
rect 980 60376 989 60416
rect 11320 60376 12652 60416
rect 12692 60376 12701 60416
rect 14659 60376 14668 60416
rect 14708 60376 15052 60416
rect 15092 60376 15101 60416
rect 0 60356 80 60376
rect 12835 60292 12844 60332
rect 12884 60292 13804 60332
rect 13844 60292 17164 60332
rect 17204 60292 17213 60332
rect 17443 60292 17452 60332
rect 17492 60292 18124 60332
rect 18164 60292 18173 60332
rect 4387 60248 4445 60249
rect 21424 60248 21504 60268
rect 4387 60208 4396 60248
rect 4436 60208 9196 60248
rect 9236 60208 9245 60248
rect 20227 60208 20236 60248
rect 20276 60208 21504 60248
rect 4387 60207 4445 60208
rect 21424 60188 21504 60208
rect 15235 60164 15293 60165
rect 4867 60124 4876 60164
rect 4916 60124 6700 60164
rect 6740 60124 7756 60164
rect 7796 60124 7805 60164
rect 12931 60124 12940 60164
rect 12980 60124 12989 60164
rect 15235 60124 15244 60164
rect 15284 60124 15628 60164
rect 15668 60124 15677 60164
rect 3139 60080 3197 60081
rect 6115 60080 6173 60081
rect 6691 60080 6749 60081
rect 8515 60080 8573 60081
rect 3043 60040 3052 60080
rect 3092 60040 3148 60080
rect 3188 60040 4204 60080
rect 4244 60040 4253 60080
rect 6115 60040 6124 60080
rect 6164 60040 6220 60080
rect 6260 60040 6269 60080
rect 6595 60040 6604 60080
rect 6644 60040 6700 60080
rect 6740 60040 7468 60080
rect 7508 60040 7517 60080
rect 7843 60040 7852 60080
rect 7892 60040 8524 60080
rect 8564 60040 8573 60080
rect 10435 60040 10444 60080
rect 10484 60040 12076 60080
rect 12116 60040 12748 60080
rect 12788 60040 12797 60080
rect 3139 60039 3197 60040
rect 6115 60039 6173 60040
rect 6691 60039 6749 60040
rect 8515 60039 8573 60040
rect 12940 59996 12980 60124
rect 15235 60123 15293 60124
rect 13315 60040 13324 60080
rect 13364 60040 15052 60080
rect 15092 60040 15101 60080
rect 15427 60040 15436 60080
rect 15476 60040 16108 60080
rect 16148 60040 16157 60080
rect 16579 60040 16588 60080
rect 16628 60040 17260 60080
rect 17300 60040 19372 60080
rect 19412 60040 19421 60080
rect 11491 59956 11500 59996
rect 11540 59956 12844 59996
rect 12884 59956 12980 59996
rect 14092 59956 14668 59996
rect 14708 59956 16012 59996
rect 16052 59956 16061 59996
rect 16867 59956 16876 59996
rect 16916 59956 17644 59996
rect 17684 59956 17693 59996
rect 6691 59872 6700 59912
rect 6740 59872 7180 59912
rect 7220 59872 7229 59912
rect 7555 59872 7564 59912
rect 7604 59872 7852 59912
rect 7892 59872 7901 59912
rect 9859 59872 9868 59912
rect 9908 59872 13708 59912
rect 13748 59872 13757 59912
rect 11971 59828 12029 59829
rect 14092 59828 14132 59956
rect 21424 59912 21504 59932
rect 163 59788 172 59828
rect 212 59788 11980 59828
rect 12020 59788 12029 59828
rect 12931 59788 12940 59828
rect 12980 59788 14132 59828
rect 14572 59872 18220 59912
rect 18260 59872 18269 59912
rect 19939 59872 19948 59912
rect 19988 59872 21504 59912
rect 11971 59787 12029 59788
rect 0 59744 80 59764
rect 9475 59744 9533 59745
rect 14083 59744 14141 59745
rect 0 59704 364 59744
rect 404 59704 413 59744
rect 4919 59704 4928 59744
rect 4968 59704 5010 59744
rect 5050 59704 5092 59744
rect 5132 59704 5174 59744
rect 5214 59704 5256 59744
rect 5296 59704 5305 59744
rect 9379 59704 9388 59744
rect 9428 59704 9484 59744
rect 9524 59704 9533 59744
rect 9955 59704 9964 59744
rect 10004 59704 13804 59744
rect 13844 59704 13853 59744
rect 14083 59704 14092 59744
rect 14132 59704 14284 59744
rect 14324 59704 14333 59744
rect 0 59684 80 59704
rect 9475 59703 9533 59704
rect 14083 59703 14141 59704
rect 13411 59660 13469 59661
rect 4195 59620 4204 59660
rect 4244 59620 9676 59660
rect 9716 59620 10252 59660
rect 10292 59620 10301 59660
rect 11395 59620 11404 59660
rect 11444 59620 13420 59660
rect 13460 59620 13469 59660
rect 13699 59620 13708 59660
rect 13748 59620 13996 59660
rect 14036 59620 14045 59660
rect 13411 59619 13469 59620
rect 3235 59576 3293 59577
rect 14572 59576 14612 59872
rect 21424 59852 21504 59872
rect 3150 59536 3244 59576
rect 3284 59536 3293 59576
rect 7843 59536 7852 59576
rect 7892 59536 14612 59576
rect 14668 59788 19756 59828
rect 19796 59788 19805 59828
rect 3235 59535 3293 59536
rect 14668 59492 14708 59788
rect 15235 59744 15293 59745
rect 15235 59704 15244 59744
rect 15284 59704 18124 59744
rect 18164 59704 18173 59744
rect 20039 59704 20048 59744
rect 20088 59704 20130 59744
rect 20170 59704 20212 59744
rect 20252 59704 20294 59744
rect 20334 59704 20376 59744
rect 20416 59704 20425 59744
rect 15235 59703 15293 59704
rect 15907 59660 15965 59661
rect 15822 59620 15916 59660
rect 15956 59620 15965 59660
rect 16104 59620 16113 59660
rect 16153 59620 16972 59660
rect 17012 59620 17021 59660
rect 15907 59619 15965 59620
rect 16867 59576 16925 59577
rect 21424 59576 21504 59596
rect 16782 59536 16876 59576
rect 16916 59536 16925 59576
rect 19171 59536 19180 59576
rect 19220 59536 19892 59576
rect 19939 59536 19948 59576
rect 19988 59536 21504 59576
rect 16867 59535 16925 59536
rect 4867 59452 4876 59492
rect 4916 59452 14708 59492
rect 15340 59452 19796 59492
rect 15340 59408 15380 59452
rect 1315 59368 1324 59408
rect 1364 59368 2284 59408
rect 2324 59368 2540 59408
rect 2755 59368 2764 59408
rect 2804 59368 3244 59408
rect 3284 59368 3293 59408
rect 3715 59368 3724 59408
rect 3764 59368 5452 59408
rect 5492 59368 5501 59408
rect 6019 59368 6028 59408
rect 6068 59368 6077 59408
rect 6979 59368 6988 59408
rect 7028 59368 15380 59408
rect 15427 59368 15436 59408
rect 15476 59368 15916 59408
rect 15956 59368 15965 59408
rect 16012 59368 19412 59408
rect 2500 59324 2540 59368
rect 6028 59324 6068 59368
rect 16012 59324 16052 59368
rect 18691 59324 18749 59325
rect 19372 59324 19412 59368
rect 19756 59324 19796 59452
rect 19852 59408 19892 59536
rect 21424 59516 21504 59536
rect 19843 59368 19852 59408
rect 19892 59368 19901 59408
rect 2500 59284 6412 59324
rect 6452 59284 7852 59324
rect 7892 59284 7901 59324
rect 14380 59284 16052 59324
rect 18499 59284 18508 59324
rect 18548 59284 18700 59324
rect 18740 59284 18749 59324
rect 19363 59284 19372 59324
rect 19412 59284 19421 59324
rect 19747 59284 19756 59324
rect 19796 59284 19805 59324
rect 4195 59240 4253 59241
rect 10051 59240 10109 59241
rect 11299 59240 11357 59241
rect 14380 59240 14420 59284
rect 18691 59283 18749 59284
rect 21424 59240 21504 59260
rect 4110 59200 4204 59240
rect 4244 59200 4253 59240
rect 6787 59200 6796 59240
rect 6836 59200 7180 59240
rect 7220 59200 8812 59240
rect 8852 59200 8861 59240
rect 9966 59200 10060 59240
rect 10100 59200 10109 59240
rect 10915 59200 10924 59240
rect 10964 59200 11308 59240
rect 11348 59200 11357 59240
rect 13795 59200 13804 59240
rect 13844 59200 14420 59240
rect 20140 59200 21504 59240
rect 4195 59199 4253 59200
rect 10051 59199 10109 59200
rect 11299 59199 11357 59200
rect 2947 59156 3005 59157
rect 20140 59156 20180 59200
rect 21424 59180 21504 59200
rect 2755 59116 2764 59156
rect 2804 59116 2956 59156
rect 2996 59116 3148 59156
rect 3188 59116 3628 59156
rect 3668 59116 3677 59156
rect 8227 59116 8236 59156
rect 8276 59116 8620 59156
rect 8660 59116 10636 59156
rect 10676 59116 10685 59156
rect 15715 59116 15724 59156
rect 15764 59116 17260 59156
rect 17300 59116 17309 59156
rect 19939 59116 19948 59156
rect 19988 59116 20180 59156
rect 2947 59115 3005 59116
rect 0 59072 80 59092
rect 3628 59072 3668 59116
rect 0 59032 172 59072
rect 212 59032 221 59072
rect 3628 59032 17068 59072
rect 17108 59032 17548 59072
rect 17588 59032 17597 59072
rect 0 59012 80 59032
rect 15907 58988 15965 58989
rect 3679 58948 3688 58988
rect 3728 58948 3770 58988
rect 3810 58948 3852 58988
rect 3892 58948 3934 58988
rect 3974 58948 4016 58988
rect 4056 58948 4065 58988
rect 5347 58948 5356 58988
rect 5396 58948 5932 58988
rect 5972 58948 5981 58988
rect 9091 58948 9100 58988
rect 9140 58948 11020 58988
rect 11060 58948 11069 58988
rect 15907 58948 15916 58988
rect 15956 58948 16204 58988
rect 16244 58948 16253 58988
rect 18799 58948 18808 58988
rect 18848 58948 18890 58988
rect 18930 58948 18972 58988
rect 19012 58948 19054 58988
rect 19094 58948 19136 58988
rect 19176 58948 19185 58988
rect 15907 58947 15965 58948
rect 21424 58904 21504 58924
rect 9283 58864 9292 58904
rect 9332 58864 9964 58904
rect 10004 58864 10013 58904
rect 20707 58864 20716 58904
rect 20756 58864 21504 58904
rect 21424 58844 21504 58864
rect 5635 58820 5693 58821
rect 13027 58820 13085 58821
rect 2659 58780 2668 58820
rect 2708 58780 4300 58820
rect 4340 58780 4780 58820
rect 4820 58780 4829 58820
rect 5616 58780 5644 58820
rect 5684 58780 5740 58820
rect 5780 58780 10348 58820
rect 10388 58780 10397 58820
rect 13027 58780 13036 58820
rect 13076 58780 13420 58820
rect 13460 58780 13469 58820
rect 15331 58780 15340 58820
rect 15380 58780 16972 58820
rect 17012 58780 17021 58820
rect 5635 58779 5693 58780
rect 13027 58779 13085 58780
rect 7843 58736 7901 58737
rect 4099 58696 4108 58736
rect 4148 58696 4492 58736
rect 4532 58696 5836 58736
rect 5876 58696 5885 58736
rect 7651 58696 7660 58736
rect 7700 58696 7852 58736
rect 7892 58696 9388 58736
rect 9428 58696 9868 58736
rect 9908 58696 9917 58736
rect 13324 58696 13708 58736
rect 13748 58696 13757 58736
rect 18403 58696 18412 58736
rect 18452 58696 18796 58736
rect 18836 58696 18845 58736
rect 7843 58695 7901 58696
rect 2083 58612 2092 58652
rect 2132 58612 12596 58652
rect 2563 58568 2621 58569
rect 6307 58568 6365 58569
rect 7651 58568 7709 58569
rect 2563 58528 2572 58568
rect 2612 58528 3532 58568
rect 3572 58528 3581 58568
rect 6222 58528 6316 58568
rect 6356 58528 7660 58568
rect 7700 58528 7709 58568
rect 2563 58527 2621 58528
rect 6307 58527 6365 58528
rect 7651 58527 7709 58528
rect 7939 58568 7997 58569
rect 11395 58568 11453 58569
rect 11779 58568 11837 58569
rect 7939 58528 7948 58568
rect 7988 58528 8044 58568
rect 8084 58528 8093 58568
rect 9955 58528 9964 58568
rect 10004 58528 11404 58568
rect 11444 58528 11453 58568
rect 11694 58528 11788 58568
rect 11828 58528 11837 58568
rect 7939 58527 7997 58528
rect 11395 58527 11453 58528
rect 11779 58527 11837 58528
rect 3235 58484 3293 58485
rect 12556 58484 12596 58612
rect 12739 58568 12797 58569
rect 13324 58568 13364 58696
rect 13411 58612 13420 58652
rect 13460 58612 19756 58652
rect 19796 58612 19805 58652
rect 12739 58528 12748 58568
rect 12788 58528 13364 58568
rect 16675 58568 16733 58569
rect 18019 58568 18077 58569
rect 21424 58568 21504 58588
rect 16675 58528 16684 58568
rect 16724 58528 16780 58568
rect 16820 58528 16829 58568
rect 17635 58528 17644 58568
rect 17684 58528 18028 58568
rect 18068 58528 18077 58568
rect 12739 58527 12797 58528
rect 16675 58527 16733 58528
rect 18019 58527 18077 58528
rect 21292 58528 21504 58568
rect 3235 58444 3244 58484
rect 3284 58444 5356 58484
rect 5396 58444 5405 58484
rect 6691 58444 6700 58484
rect 6740 58444 7180 58484
rect 7220 58444 8140 58484
rect 8180 58444 10156 58484
rect 10196 58444 10205 58484
rect 10435 58444 10444 58484
rect 10484 58444 10924 58484
rect 10964 58444 11212 58484
rect 11252 58444 11261 58484
rect 12556 58444 13804 58484
rect 13844 58444 13853 58484
rect 3235 58443 3293 58444
rect 0 58400 80 58420
rect 21292 58400 21332 58528
rect 21424 58508 21504 58528
rect 0 58360 6220 58400
rect 6260 58360 6269 58400
rect 7363 58360 7372 58400
rect 7412 58360 21332 58400
rect 0 58340 80 58360
rect 2851 58316 2909 58317
rect 2851 58276 2860 58316
rect 2900 58276 4780 58316
rect 4820 58276 4829 58316
rect 2851 58275 2909 58276
rect 21424 58232 21504 58252
rect 4919 58192 4928 58232
rect 4968 58192 5010 58232
rect 5050 58192 5092 58232
rect 5132 58192 5174 58232
rect 5214 58192 5256 58232
rect 5296 58192 5305 58232
rect 14755 58192 14764 58232
rect 14804 58192 15628 58232
rect 15668 58192 15677 58232
rect 20039 58192 20048 58232
rect 20088 58192 20130 58232
rect 20170 58192 20212 58232
rect 20252 58192 20294 58232
rect 20334 58192 20376 58232
rect 20416 58192 20425 58232
rect 21187 58192 21196 58232
rect 21236 58192 21504 58232
rect 21424 58172 21504 58192
rect 17539 58108 17548 58148
rect 17588 58108 20716 58148
rect 20756 58108 20765 58148
rect 18211 58064 18269 58065
rect 3235 58024 3244 58064
rect 3284 58024 3436 58064
rect 3476 58024 12748 58064
rect 12788 58024 12797 58064
rect 15619 58024 15628 58064
rect 15668 58024 16012 58064
rect 16052 58024 16061 58064
rect 17155 58024 17164 58064
rect 17204 58024 18164 58064
rect 16099 57980 16157 57981
rect 18124 57980 18164 58024
rect 18211 58024 18220 58064
rect 18260 58024 18316 58064
rect 18356 58024 18365 58064
rect 18211 58023 18269 58024
rect 4675 57940 4684 57980
rect 4724 57940 6604 57980
rect 6644 57940 6653 57980
rect 7555 57940 7564 57980
rect 7604 57940 7948 57980
rect 7988 57940 9868 57980
rect 9908 57940 9917 57980
rect 11875 57940 11884 57980
rect 11924 57940 12172 57980
rect 12212 57940 16108 57980
rect 16148 57940 16157 57980
rect 16291 57940 16300 57980
rect 16340 57940 18028 57980
rect 18068 57940 18077 57980
rect 18124 57940 18892 57980
rect 18932 57940 18941 57980
rect 6604 57896 6644 57940
rect 16099 57939 16157 57940
rect 21424 57896 21504 57916
rect 3715 57856 3724 57896
rect 3764 57856 5260 57896
rect 5300 57856 5309 57896
rect 6604 57856 9100 57896
rect 9140 57856 9149 57896
rect 10915 57856 10924 57896
rect 10964 57856 13132 57896
rect 13172 57856 13181 57896
rect 14659 57856 14668 57896
rect 14708 57856 15244 57896
rect 15284 57856 15293 57896
rect 16771 57856 16780 57896
rect 16820 57856 17548 57896
rect 17588 57856 17597 57896
rect 17827 57856 17836 57896
rect 17876 57856 19084 57896
rect 19124 57856 19133 57896
rect 20611 57856 20620 57896
rect 20660 57856 21504 57896
rect 21424 57836 21504 57856
rect 5347 57812 5405 57813
rect 3331 57772 3340 57812
rect 3380 57772 3916 57812
rect 3956 57772 3965 57812
rect 5262 57772 5356 57812
rect 5396 57772 8840 57812
rect 17635 57772 17644 57812
rect 17684 57772 18124 57812
rect 18164 57772 18173 57812
rect 18979 57772 18988 57812
rect 19028 57772 19948 57812
rect 19988 57772 19997 57812
rect 5347 57771 5405 57772
rect 0 57728 80 57748
rect 8800 57728 8840 57772
rect 9475 57728 9533 57729
rect 18988 57728 19028 57772
rect 0 57688 2540 57728
rect 3235 57688 3244 57728
rect 3284 57688 4113 57728
rect 4153 57688 4972 57728
rect 5012 57688 5021 57728
rect 8800 57688 9484 57728
rect 9524 57688 11884 57728
rect 11924 57688 11933 57728
rect 17155 57688 17164 57728
rect 17204 57688 17740 57728
rect 17780 57688 17789 57728
rect 17836 57688 19028 57728
rect 20035 57688 20044 57728
rect 20084 57688 21004 57728
rect 21044 57688 21053 57728
rect 0 57668 80 57688
rect 1507 57604 1516 57644
rect 1556 57604 1708 57644
rect 1748 57604 1757 57644
rect 2500 57560 2540 57688
rect 9475 57687 9533 57688
rect 3434 57604 3443 57644
rect 3483 57604 3628 57644
rect 3668 57604 3677 57644
rect 4003 57604 4012 57644
rect 4052 57604 5356 57644
rect 5396 57604 5405 57644
rect 9955 57560 10013 57561
rect 17836 57560 17876 57688
rect 18691 57604 18700 57644
rect 18740 57604 20236 57644
rect 20276 57604 20285 57644
rect 21424 57560 21504 57580
rect 2500 57520 9964 57560
rect 10004 57520 10013 57560
rect 17731 57520 17740 57560
rect 17780 57520 17876 57560
rect 17932 57520 21504 57560
rect 9955 57519 10013 57520
rect 12259 57476 12317 57477
rect 17932 57476 17972 57520
rect 21424 57500 21504 57520
rect 3679 57436 3688 57476
rect 3728 57436 3770 57476
rect 3810 57436 3852 57476
rect 3892 57436 3934 57476
rect 3974 57436 4016 57476
rect 4056 57436 4065 57476
rect 6211 57436 6220 57476
rect 6260 57436 12268 57476
rect 12308 57436 12317 57476
rect 15619 57436 15628 57476
rect 15668 57436 17972 57476
rect 18799 57436 18808 57476
rect 18848 57436 18890 57476
rect 18930 57436 18972 57476
rect 19012 57436 19054 57476
rect 19094 57436 19136 57476
rect 19176 57436 19185 57476
rect 12259 57435 12317 57436
rect 4483 57392 4541 57393
rect 4483 57352 4492 57392
rect 4532 57352 7564 57392
rect 7604 57352 7613 57392
rect 11395 57352 11404 57392
rect 11444 57352 19564 57392
rect 19604 57352 19613 57392
rect 4483 57351 4541 57352
rect 8131 57308 8189 57309
rect 2755 57268 2764 57308
rect 2804 57268 3340 57308
rect 3380 57268 3389 57308
rect 7171 57268 7180 57308
rect 7220 57268 8140 57308
rect 8180 57268 8189 57308
rect 8131 57267 8189 57268
rect 13123 57308 13181 57309
rect 13123 57268 13132 57308
rect 13172 57268 13516 57308
rect 13556 57268 13565 57308
rect 18115 57268 18124 57308
rect 18164 57268 19660 57308
rect 19700 57268 19709 57308
rect 13123 57267 13181 57268
rect 20803 57224 20861 57225
rect 21424 57224 21504 57244
rect 17923 57184 17932 57224
rect 17972 57184 19948 57224
rect 19988 57184 19997 57224
rect 20803 57184 20812 57224
rect 20852 57184 21504 57224
rect 20803 57183 20861 57184
rect 21424 57164 21504 57184
rect 8131 57140 8189 57141
rect 10051 57140 10109 57141
rect 14179 57140 14237 57141
rect 17443 57140 17501 57141
rect 8131 57100 8140 57140
rect 8180 57100 8620 57140
rect 8660 57100 8669 57140
rect 9966 57100 10060 57140
rect 10100 57100 10109 57140
rect 13219 57100 13228 57140
rect 13268 57100 14188 57140
rect 14228 57100 14956 57140
rect 14996 57100 15005 57140
rect 17443 57100 17452 57140
rect 17492 57100 18028 57140
rect 18068 57100 18077 57140
rect 19180 57100 19372 57140
rect 19412 57100 19564 57140
rect 19604 57100 19613 57140
rect 8131 57099 8189 57100
rect 10051 57099 10109 57100
rect 14179 57099 14237 57100
rect 17443 57099 17501 57100
rect 0 57056 80 57076
rect 2467 57056 2525 57057
rect 16291 57056 16349 57057
rect 19180 57056 19220 57100
rect 0 57016 1900 57056
rect 1940 57016 1949 57056
rect 2467 57016 2476 57056
rect 2516 57016 2572 57056
rect 2612 57016 2860 57056
rect 2900 57016 2909 57056
rect 7171 57016 7180 57056
rect 7220 57016 8812 57056
rect 8852 57016 8861 57056
rect 11971 57016 11980 57056
rect 12020 57016 12364 57056
rect 12404 57016 12413 57056
rect 14179 57016 14188 57056
rect 14228 57016 15628 57056
rect 15668 57016 15677 57056
rect 16206 57016 16300 57056
rect 16340 57016 16349 57056
rect 0 56996 80 57016
rect 2467 57015 2525 57016
rect 16291 57015 16349 57016
rect 17548 57016 19220 57056
rect 19267 57016 19276 57056
rect 19316 57016 19948 57056
rect 19988 57016 19997 57056
rect 17548 56972 17588 57016
rect 13411 56932 13420 56972
rect 13460 56932 13708 56972
rect 13748 56932 13757 56972
rect 14659 56932 14668 56972
rect 14708 56932 16684 56972
rect 16724 56932 17548 56972
rect 17588 56932 17597 56972
rect 19459 56932 19468 56972
rect 19508 56932 19756 56972
rect 19796 56932 19805 56972
rect 19363 56888 19421 56889
rect 3043 56848 3052 56888
rect 3092 56848 3244 56888
rect 3284 56848 3293 56888
rect 7651 56848 7660 56888
rect 7700 56848 8140 56888
rect 8180 56848 8189 56888
rect 8419 56848 8428 56888
rect 8468 56848 15436 56888
rect 15476 56848 15485 56888
rect 17731 56848 17740 56888
rect 17780 56848 17932 56888
rect 17972 56848 17981 56888
rect 19267 56848 19276 56888
rect 19316 56848 19372 56888
rect 19412 56848 19421 56888
rect 19363 56847 19421 56848
rect 19555 56888 19613 56889
rect 21424 56888 21504 56908
rect 19555 56848 19564 56888
rect 19604 56848 21504 56888
rect 19555 56847 19613 56848
rect 21424 56828 21504 56848
rect 7939 56764 7948 56804
rect 7988 56764 8468 56804
rect 9091 56764 9100 56804
rect 9140 56764 9484 56804
rect 9524 56764 9533 56804
rect 14371 56764 14380 56804
rect 14420 56764 16876 56804
rect 16916 56764 16925 56804
rect 8323 56720 8381 56721
rect 2659 56680 2668 56720
rect 2708 56680 4588 56720
rect 4628 56680 4637 56720
rect 4919 56680 4928 56720
rect 4968 56680 5010 56720
rect 5050 56680 5092 56720
rect 5132 56680 5174 56720
rect 5214 56680 5256 56720
rect 5296 56680 5305 56720
rect 6979 56680 6988 56720
rect 7028 56680 8332 56720
rect 8372 56680 8381 56720
rect 8428 56720 8468 56764
rect 13411 56720 13469 56721
rect 17635 56720 17693 56721
rect 8428 56680 10636 56720
rect 10676 56680 10828 56720
rect 10868 56680 10877 56720
rect 13411 56680 13420 56720
rect 13460 56680 13612 56720
rect 13652 56680 13661 56720
rect 13891 56680 13900 56720
rect 13940 56680 17644 56720
rect 17684 56680 18028 56720
rect 18068 56680 18077 56720
rect 20039 56680 20048 56720
rect 20088 56680 20130 56720
rect 20170 56680 20212 56720
rect 20252 56680 20294 56720
rect 20334 56680 20376 56720
rect 20416 56680 20425 56720
rect 8323 56679 8381 56680
rect 13411 56679 13469 56680
rect 17635 56679 17693 56680
rect 17443 56636 17501 56637
rect 1315 56596 1324 56636
rect 1364 56596 5932 56636
rect 5972 56596 5981 56636
rect 7075 56596 7084 56636
rect 7124 56596 7276 56636
rect 7316 56596 7325 56636
rect 7468 56596 7988 56636
rect 11011 56596 11020 56636
rect 11060 56596 15764 56636
rect 16387 56596 16396 56636
rect 16436 56596 17452 56636
rect 17492 56596 17660 56636
rect 4387 56552 4445 56553
rect 1603 56512 1612 56552
rect 1652 56512 4396 56552
rect 4436 56512 4445 56552
rect 6979 56512 6988 56552
rect 7028 56512 7372 56552
rect 7412 56512 7421 56552
rect 4387 56511 4445 56512
rect 7468 56468 7508 56596
rect 2500 56428 7508 56468
rect 7756 56512 7852 56552
rect 7892 56512 7901 56552
rect 0 56384 80 56404
rect 2500 56384 2540 56428
rect 0 56344 2540 56384
rect 2755 56384 2813 56385
rect 5827 56384 5885 56385
rect 2755 56344 2764 56384
rect 2804 56344 3436 56384
rect 3476 56344 5644 56384
rect 5684 56344 5693 56384
rect 5827 56344 5836 56384
rect 5876 56344 5970 56384
rect 0 56324 80 56344
rect 2755 56343 2813 56344
rect 5827 56343 5885 56344
rect 7756 56301 7796 56512
rect 7948 56468 7988 56596
rect 13228 56512 14668 56552
rect 14708 56512 14717 56552
rect 10915 56468 10973 56469
rect 7948 56428 10924 56468
rect 10964 56428 10973 56468
rect 10915 56427 10973 56428
rect 10531 56384 10589 56385
rect 13228 56384 13268 56512
rect 15724 56468 15764 56596
rect 17443 56595 17501 56596
rect 17251 56552 17309 56553
rect 16675 56512 16684 56552
rect 16724 56512 17260 56552
rect 17300 56512 17309 56552
rect 17620 56552 17660 56596
rect 19363 56552 19421 56553
rect 21424 56552 21504 56572
rect 17620 56512 18988 56552
rect 19028 56512 19037 56552
rect 19363 56512 19372 56552
rect 19412 56512 21504 56552
rect 17251 56511 17309 56512
rect 19363 56511 19421 56512
rect 21424 56492 21504 56512
rect 15724 56428 20180 56468
rect 20140 56384 20180 56428
rect 7843 56344 7852 56384
rect 7892 56344 8236 56384
rect 8276 56344 8285 56384
rect 8899 56344 8908 56384
rect 8948 56344 8957 56384
rect 9667 56344 9676 56384
rect 9716 56344 10540 56384
rect 10580 56344 10589 56384
rect 12451 56344 12460 56384
rect 12500 56344 13228 56384
rect 13268 56344 13277 56384
rect 14275 56344 14284 56384
rect 14324 56344 14668 56384
rect 14708 56344 16780 56384
rect 16820 56344 16829 56384
rect 16963 56344 16972 56384
rect 17012 56344 17740 56384
rect 17780 56344 19468 56384
rect 19508 56344 19517 56384
rect 20140 56344 21388 56384
rect 21428 56344 21437 56384
rect 7747 56300 7805 56301
rect 2500 56260 7756 56300
rect 7796 56260 7805 56300
rect 2500 56048 2540 56260
rect 7747 56259 7805 56260
rect 3523 56216 3581 56217
rect 7852 56216 7892 56344
rect 3523 56176 3532 56216
rect 3572 56176 3628 56216
rect 3668 56176 3677 56216
rect 6787 56176 6796 56216
rect 6836 56176 7276 56216
rect 7316 56176 7325 56216
rect 7555 56176 7564 56216
rect 7604 56176 7892 56216
rect 8323 56216 8381 56217
rect 8323 56176 8332 56216
rect 8372 56176 8428 56216
rect 8468 56176 8477 56216
rect 3523 56175 3581 56176
rect 8323 56175 8381 56176
rect 2659 56132 2717 56133
rect 7651 56132 7709 56133
rect 8908 56132 8948 56344
rect 10531 56343 10589 56344
rect 14179 56300 14237 56301
rect 17347 56300 17405 56301
rect 9475 56260 9484 56300
rect 9524 56260 10924 56300
rect 10964 56260 10973 56300
rect 14179 56260 14188 56300
rect 14228 56260 16492 56300
rect 16532 56260 16541 56300
rect 16867 56260 16876 56300
rect 16916 56260 17356 56300
rect 17396 56260 17405 56300
rect 14179 56259 14237 56260
rect 17347 56259 17405 56260
rect 21424 56216 21504 56236
rect 20803 56176 20812 56216
rect 20852 56176 21504 56216
rect 21424 56156 21504 56176
rect 2659 56092 2668 56132
rect 2708 56092 7660 56132
rect 7700 56092 7709 56132
rect 7939 56092 7948 56132
rect 7988 56092 8948 56132
rect 9283 56092 9292 56132
rect 9332 56092 9868 56132
rect 9908 56092 12596 56132
rect 13699 56092 13708 56132
rect 13748 56092 14668 56132
rect 14708 56092 14717 56132
rect 2659 56091 2717 56092
rect 7651 56091 7709 56092
rect 11587 56048 11645 56049
rect 12451 56048 12509 56049
rect 1411 56008 1420 56048
rect 1460 56008 2188 56048
rect 2228 56008 2540 56048
rect 4483 56008 4492 56048
rect 4532 56008 11596 56048
rect 11636 56008 12460 56048
rect 12500 56008 12509 56048
rect 11587 56007 11645 56008
rect 12451 56007 12509 56008
rect 3043 55964 3101 55965
rect 12556 55964 12596 56092
rect 13987 56008 13996 56048
rect 14036 56008 18220 56048
rect 18260 56008 18269 56048
rect 3043 55924 3052 55964
rect 3092 55924 3532 55964
rect 3572 55924 3581 55964
rect 3679 55924 3688 55964
rect 3728 55924 3770 55964
rect 3810 55924 3852 55964
rect 3892 55924 3934 55964
rect 3974 55924 4016 55964
rect 4056 55924 4065 55964
rect 5155 55924 5164 55964
rect 5204 55924 5356 55964
rect 5396 55924 11020 55964
rect 11060 55924 11069 55964
rect 12556 55924 18412 55964
rect 18452 55924 18461 55964
rect 18799 55924 18808 55964
rect 18848 55924 18890 55964
rect 18930 55924 18972 55964
rect 19012 55924 19054 55964
rect 19094 55924 19136 55964
rect 19176 55924 19185 55964
rect 3043 55923 3101 55924
rect 21424 55880 21504 55900
rect 4108 55840 13268 55880
rect 15715 55840 15724 55880
rect 15764 55840 20812 55880
rect 20852 55840 20861 55880
rect 21379 55840 21388 55880
rect 21428 55840 21504 55880
rect 4108 55797 4148 55840
rect 4099 55796 4157 55797
rect 4099 55756 4108 55796
rect 4148 55756 4157 55796
rect 5923 55756 5932 55796
rect 5972 55756 6220 55796
rect 6260 55756 8140 55796
rect 8180 55756 8620 55796
rect 8660 55756 8669 55796
rect 4099 55755 4157 55756
rect 0 55712 80 55732
rect 13228 55712 13268 55840
rect 21424 55820 21504 55840
rect 16675 55796 16733 55797
rect 16483 55756 16492 55796
rect 16532 55756 16684 55796
rect 16724 55756 16733 55796
rect 17155 55756 17164 55796
rect 17204 55756 17452 55796
rect 17492 55756 17501 55796
rect 19459 55756 19468 55796
rect 19508 55756 19852 55796
rect 19892 55756 19901 55796
rect 16675 55755 16733 55756
rect 0 55672 1324 55712
rect 1364 55672 1373 55712
rect 4003 55672 4012 55712
rect 4052 55672 4588 55712
rect 4628 55672 4637 55712
rect 6787 55672 6796 55712
rect 6836 55672 8332 55712
rect 8372 55672 9100 55712
rect 9140 55672 9149 55712
rect 10051 55672 10060 55712
rect 10100 55672 10348 55712
rect 10388 55672 10397 55712
rect 13228 55672 21332 55712
rect 0 55652 80 55672
rect 7747 55628 7805 55629
rect 14851 55628 14909 55629
rect 3244 55588 4204 55628
rect 4244 55588 4253 55628
rect 6595 55588 6604 55628
rect 6644 55588 7316 55628
rect 3244 55544 3284 55588
rect 7276 55544 7316 55588
rect 7747 55588 7756 55628
rect 7796 55588 8620 55628
rect 8660 55588 11212 55628
rect 11252 55588 11261 55628
rect 11320 55588 12076 55628
rect 12116 55588 12125 55628
rect 12451 55588 12460 55628
rect 12500 55588 14860 55628
rect 14900 55588 14909 55628
rect 15811 55588 15820 55628
rect 15860 55588 17548 55628
rect 17588 55588 17597 55628
rect 7747 55587 7805 55588
rect 10147 55544 10205 55545
rect 11320 55544 11360 55588
rect 14851 55587 14909 55588
rect 3235 55504 3244 55544
rect 3284 55504 3293 55544
rect 3907 55504 3916 55544
rect 3956 55504 3965 55544
rect 6691 55504 6700 55544
rect 6740 55504 6749 55544
rect 7267 55504 7276 55544
rect 7316 55504 7325 55544
rect 7459 55504 7468 55544
rect 7508 55504 7756 55544
rect 7796 55504 7805 55544
rect 7852 55504 10100 55544
rect 3916 55376 3956 55504
rect 2755 55336 2764 55376
rect 2804 55336 3628 55376
rect 3668 55336 3956 55376
rect 6700 55376 6740 55504
rect 7651 55460 7709 55461
rect 7852 55460 7892 55504
rect 7651 55420 7660 55460
rect 7700 55420 7892 55460
rect 10060 55460 10100 55504
rect 10147 55504 10156 55544
rect 10196 55504 10252 55544
rect 10292 55504 10301 55544
rect 10348 55504 11360 55544
rect 13411 55544 13469 55545
rect 21292 55544 21332 55672
rect 21424 55544 21504 55564
rect 13411 55504 13420 55544
rect 13460 55504 15724 55544
rect 15764 55504 15773 55544
rect 16099 55504 16108 55544
rect 16148 55504 16972 55544
rect 17012 55504 17021 55544
rect 17635 55504 17644 55544
rect 17684 55504 17693 55544
rect 19363 55504 19372 55544
rect 19412 55504 19660 55544
rect 19700 55504 19709 55544
rect 21292 55504 21504 55544
rect 10147 55503 10205 55504
rect 10348 55460 10388 55504
rect 13411 55503 13469 55504
rect 14851 55460 14909 55461
rect 10060 55420 10388 55460
rect 14820 55420 14860 55460
rect 14900 55420 14909 55460
rect 17644 55460 17684 55504
rect 21424 55484 21504 55504
rect 18691 55460 18749 55461
rect 19459 55460 19517 55461
rect 17644 55420 18700 55460
rect 18740 55420 19468 55460
rect 19508 55420 19517 55460
rect 7651 55419 7709 55420
rect 14851 55419 14909 55420
rect 18691 55419 18749 55420
rect 19459 55419 19517 55420
rect 14860 55376 14900 55419
rect 6700 55336 7756 55376
rect 7796 55336 7805 55376
rect 14467 55336 14476 55376
rect 14516 55336 14900 55376
rect 19843 55336 19852 55376
rect 19892 55336 20140 55376
rect 20180 55336 20189 55376
rect 4492 55252 9676 55292
rect 9716 55252 9725 55292
rect 2851 55084 2860 55124
rect 2900 55084 3340 55124
rect 3380 55084 3389 55124
rect 0 55040 80 55060
rect 0 55000 1612 55040
rect 1652 55000 1661 55040
rect 0 54980 80 55000
rect 4492 54956 4532 55252
rect 15907 55208 15965 55209
rect 21424 55208 21504 55228
rect 4919 55168 4928 55208
rect 4968 55168 5010 55208
rect 5050 55168 5092 55208
rect 5132 55168 5174 55208
rect 5214 55168 5256 55208
rect 5296 55168 5305 55208
rect 6499 55168 6508 55208
rect 6548 55168 6988 55208
rect 7028 55168 7037 55208
rect 7171 55168 7180 55208
rect 7220 55168 7229 55208
rect 10627 55168 10636 55208
rect 10676 55168 10828 55208
rect 10868 55168 10877 55208
rect 15822 55168 15916 55208
rect 15956 55168 15965 55208
rect 20039 55168 20048 55208
rect 20088 55168 20130 55208
rect 20170 55168 20212 55208
rect 20252 55168 20294 55208
rect 20334 55168 20376 55208
rect 20416 55168 20425 55208
rect 20524 55168 21504 55208
rect 6595 55124 6653 55125
rect 7180 55124 7220 55168
rect 15907 55167 15965 55168
rect 6595 55084 6604 55124
rect 6644 55084 7220 55124
rect 19651 55124 19709 55125
rect 20524 55124 20564 55168
rect 21424 55148 21504 55168
rect 19651 55084 19660 55124
rect 19700 55084 20564 55124
rect 6595 55083 6653 55084
rect 19651 55083 19709 55084
rect 15811 55040 15869 55041
rect 6403 55000 6412 55040
rect 6452 55000 6796 55040
rect 6836 55000 6845 55040
rect 6979 55000 6988 55040
rect 7028 55000 7468 55040
rect 7508 55000 7517 55040
rect 9859 55000 9868 55040
rect 9908 55000 11828 55040
rect 11788 54956 11828 55000
rect 15811 55000 15820 55040
rect 15860 55000 15916 55040
rect 15956 55000 15965 55040
rect 16291 55000 16300 55040
rect 16340 55000 17836 55040
rect 17876 55000 17885 55040
rect 18115 55000 18124 55040
rect 18164 55000 18173 55040
rect 18499 55000 18508 55040
rect 18548 55000 19564 55040
rect 19604 55000 19613 55040
rect 15811 54999 15869 55000
rect 14179 54956 14237 54957
rect 18124 54956 18164 55000
rect 1411 54916 1420 54956
rect 1460 54916 4532 54956
rect 7555 54916 7564 54956
rect 7604 54916 10156 54956
rect 10196 54916 10205 54956
rect 11779 54916 11788 54956
rect 11828 54916 14188 54956
rect 14228 54916 14237 54956
rect 17443 54916 17452 54956
rect 17492 54916 18164 54956
rect 14179 54915 14237 54916
rect 21424 54872 21504 54892
rect 2500 54832 3340 54872
rect 3380 54832 9004 54872
rect 9044 54832 9053 54872
rect 10243 54832 10252 54872
rect 10292 54832 11404 54872
rect 11444 54832 11453 54872
rect 13219 54832 13228 54872
rect 13268 54832 19948 54872
rect 19988 54832 19997 54872
rect 20140 54832 21504 54872
rect 1987 54788 2045 54789
rect 2500 54788 2540 54832
rect 4099 54788 4157 54789
rect 8995 54788 9053 54789
rect 1987 54748 1996 54788
rect 2036 54748 2540 54788
rect 3139 54748 3148 54788
rect 3188 54748 4108 54788
rect 4148 54748 4157 54788
rect 8323 54748 8332 54788
rect 8372 54748 9004 54788
rect 9044 54748 9053 54788
rect 9667 54748 9676 54788
rect 9716 54748 10540 54788
rect 10580 54748 11360 54788
rect 1987 54747 2045 54748
rect 4099 54747 4157 54748
rect 8995 54747 9053 54748
rect 10051 54704 10109 54705
rect 11320 54704 11360 54748
rect 13228 54704 13268 54832
rect 18211 54788 18269 54789
rect 17539 54748 17548 54788
rect 17588 54748 18220 54788
rect 18260 54748 19372 54788
rect 19412 54748 19421 54788
rect 18211 54747 18269 54748
rect 2659 54664 2668 54704
rect 2708 54664 4588 54704
rect 4628 54664 5740 54704
rect 5780 54664 6796 54704
rect 6836 54664 7084 54704
rect 7124 54664 8140 54704
rect 8180 54664 8189 54704
rect 10051 54664 10060 54704
rect 10100 54664 10156 54704
rect 10196 54664 10205 54704
rect 11320 54664 13268 54704
rect 10051 54663 10109 54664
rect 10819 54620 10877 54621
rect 11683 54620 11741 54621
rect 16675 54620 16733 54621
rect 20140 54620 20180 54832
rect 21424 54812 21504 54832
rect 5539 54580 5548 54620
rect 5588 54580 10828 54620
rect 10868 54580 11692 54620
rect 11732 54580 11741 54620
rect 16590 54580 16684 54620
rect 16724 54580 16733 54620
rect 17155 54580 17164 54620
rect 17204 54580 20180 54620
rect 10819 54579 10877 54580
rect 11683 54579 11741 54580
rect 16675 54579 16733 54580
rect 2755 54536 2813 54537
rect 21424 54536 21504 54556
rect 2755 54496 2764 54536
rect 2804 54496 8084 54536
rect 9475 54496 9484 54536
rect 9524 54496 21504 54536
rect 2755 54495 2813 54496
rect 3679 54412 3688 54452
rect 3728 54412 3770 54452
rect 3810 54412 3852 54452
rect 3892 54412 3934 54452
rect 3974 54412 4016 54452
rect 4056 54412 4065 54452
rect 5644 54412 7372 54452
rect 7412 54412 7421 54452
rect 0 54368 80 54388
rect 3523 54368 3581 54369
rect 5644 54368 5684 54412
rect 8044 54368 8084 54496
rect 21424 54476 21504 54496
rect 11395 54452 11453 54453
rect 15235 54452 15293 54453
rect 8995 54412 9004 54452
rect 9044 54412 11404 54452
rect 11444 54412 11453 54452
rect 14371 54412 14380 54452
rect 14420 54412 15244 54452
rect 15284 54412 15293 54452
rect 18799 54412 18808 54452
rect 18848 54412 18890 54452
rect 18930 54412 18972 54452
rect 19012 54412 19054 54452
rect 19094 54412 19136 54452
rect 19176 54412 19185 54452
rect 11395 54411 11453 54412
rect 15235 54411 15293 54412
rect 0 54328 1420 54368
rect 1460 54328 1469 54368
rect 3523 54328 3532 54368
rect 3572 54328 5684 54368
rect 5731 54328 5740 54368
rect 5780 54328 6124 54368
rect 6164 54328 6173 54368
rect 6307 54328 6316 54368
rect 6356 54328 7988 54368
rect 8044 54328 14860 54368
rect 14900 54328 14909 54368
rect 0 54308 80 54328
rect 3523 54327 3581 54328
rect 3724 54284 3764 54328
rect 3715 54244 3724 54284
rect 3764 54244 3773 54284
rect 5827 54244 5836 54284
rect 5876 54244 7852 54284
rect 7892 54244 7901 54284
rect 1027 54200 1085 54201
rect 942 54160 1036 54200
rect 1076 54160 1085 54200
rect 1027 54159 1085 54160
rect 3523 54200 3581 54201
rect 5731 54200 5789 54201
rect 3523 54160 3532 54200
rect 3572 54160 5452 54200
rect 5492 54160 5501 54200
rect 5731 54160 5740 54200
rect 5780 54160 6796 54200
rect 6836 54160 6845 54200
rect 7171 54160 7180 54200
rect 7220 54160 7564 54200
rect 7604 54160 7613 54200
rect 3523 54159 3581 54160
rect 5731 54159 5789 54160
rect 7948 54116 7988 54328
rect 8995 54284 9053 54285
rect 9475 54284 9533 54285
rect 8995 54244 9004 54284
rect 9044 54244 9484 54284
rect 9524 54244 9533 54284
rect 10051 54244 10060 54284
rect 10100 54244 10109 54284
rect 8995 54243 9053 54244
rect 9475 54243 9533 54244
rect 10060 54200 10100 54244
rect 21424 54201 21504 54220
rect 10915 54200 10973 54201
rect 12931 54200 12989 54201
rect 21379 54200 21504 54201
rect 8611 54160 8620 54200
rect 8660 54160 9676 54200
rect 9716 54160 10540 54200
rect 10580 54160 10589 54200
rect 10830 54160 10924 54200
rect 10964 54160 10973 54200
rect 12846 54160 12940 54200
rect 12980 54160 12989 54200
rect 15139 54160 15148 54200
rect 15188 54160 15197 54200
rect 15331 54160 15340 54200
rect 15380 54160 16588 54200
rect 16628 54160 16637 54200
rect 17251 54160 17260 54200
rect 17300 54160 17548 54200
rect 17588 54160 17597 54200
rect 18211 54160 18220 54200
rect 18260 54160 19852 54200
rect 19892 54160 19901 54200
rect 21379 54160 21388 54200
rect 21428 54160 21504 54200
rect 10915 54159 10973 54160
rect 12931 54159 12989 54160
rect 10147 54116 10205 54117
rect 7948 54076 9100 54116
rect 9140 54076 9149 54116
rect 9571 54076 9580 54116
rect 9620 54076 10156 54116
rect 10196 54076 10205 54116
rect 9100 54032 9140 54076
rect 10147 54075 10205 54076
rect 2500 53992 7276 54032
rect 7316 53992 7325 54032
rect 7939 53992 7948 54032
rect 7988 53992 8524 54032
rect 8564 53992 8573 54032
rect 8707 53992 8716 54032
rect 8756 53992 9004 54032
rect 9044 53992 9053 54032
rect 9100 53992 9676 54032
rect 9716 53992 9725 54032
rect 10051 53992 10060 54032
rect 10100 53992 10109 54032
rect 11491 53992 11500 54032
rect 11540 53992 12076 54032
rect 12116 53992 12125 54032
rect 12643 53992 12652 54032
rect 12692 53992 13804 54032
rect 13844 53992 13853 54032
rect 13987 53992 13996 54032
rect 14036 53992 14188 54032
rect 14228 53992 14237 54032
rect 2500 53948 2540 53992
rect 10060 53948 10100 53992
rect 14179 53948 14237 53949
rect 2275 53908 2284 53948
rect 2324 53908 2540 53948
rect 3619 53908 3628 53948
rect 3668 53908 6604 53948
rect 6644 53908 6653 53948
rect 6700 53908 10100 53948
rect 11203 53908 11212 53948
rect 11252 53908 14188 53948
rect 14228 53908 14237 53948
rect 6700 53864 6740 53908
rect 14179 53907 14237 53908
rect 14563 53948 14621 53949
rect 14563 53908 14572 53948
rect 14612 53908 14668 53948
rect 14708 53908 14717 53948
rect 14563 53907 14621 53908
rect 8515 53864 8573 53865
rect 15148 53864 15188 54160
rect 21379 54159 21504 54160
rect 21424 54140 21504 54159
rect 17443 54116 17501 54117
rect 16675 54076 16684 54116
rect 16724 54076 17452 54116
rect 17492 54076 18932 54116
rect 17443 54075 17501 54076
rect 17635 54032 17693 54033
rect 18892 54032 18932 54076
rect 19939 54032 19997 54033
rect 17635 53992 17644 54032
rect 17684 53992 17932 54032
rect 17972 53992 17981 54032
rect 18883 53992 18892 54032
rect 18932 53992 18941 54032
rect 19854 53992 19948 54032
rect 19988 53992 19997 54032
rect 17635 53991 17693 53992
rect 19939 53991 19997 53992
rect 16867 53948 16925 53949
rect 15331 53908 15340 53948
rect 15380 53908 16012 53948
rect 16052 53908 16061 53948
rect 16867 53908 16876 53948
rect 16916 53908 17164 53948
rect 17204 53908 18316 53948
rect 18356 53908 18365 53948
rect 16867 53907 16925 53908
rect 21424 53864 21504 53884
rect 4291 53824 4300 53864
rect 4340 53824 4876 53864
rect 4916 53824 4925 53864
rect 5059 53824 5068 53864
rect 5108 53824 5117 53864
rect 5251 53824 5260 53864
rect 5300 53824 6316 53864
rect 6356 53824 6365 53864
rect 6691 53824 6700 53864
rect 6740 53824 6749 53864
rect 8419 53824 8428 53864
rect 8468 53824 8524 53864
rect 8564 53824 8573 53864
rect 10723 53824 10732 53864
rect 10772 53824 11596 53864
rect 11636 53824 11645 53864
rect 13507 53824 13516 53864
rect 13556 53824 13565 53864
rect 15139 53824 15148 53864
rect 15188 53824 15197 53864
rect 15619 53824 15628 53864
rect 15668 53824 16204 53864
rect 16244 53824 17452 53864
rect 17492 53824 17501 53864
rect 20140 53824 21504 53864
rect 5068 53780 5108 53824
rect 8515 53823 8573 53824
rect 9763 53780 9821 53781
rect 13219 53780 13277 53781
rect 13516 53780 13556 53824
rect 17251 53780 17309 53781
rect 20140 53780 20180 53824
rect 21424 53804 21504 53824
rect 4099 53740 4108 53780
rect 4148 53740 4396 53780
rect 4436 53740 4445 53780
rect 5068 53740 5876 53780
rect 6403 53740 6412 53780
rect 6452 53740 9580 53780
rect 9620 53740 9629 53780
rect 9763 53740 9772 53780
rect 9812 53740 9964 53780
rect 10004 53740 10013 53780
rect 13219 53740 13228 53780
rect 13268 53740 16244 53780
rect 0 53696 80 53716
rect 5347 53696 5405 53697
rect 5836 53696 5876 53740
rect 9763 53739 9821 53740
rect 13219 53739 13277 53740
rect 15907 53696 15965 53697
rect 0 53656 1228 53696
rect 1268 53656 1277 53696
rect 3235 53656 3244 53696
rect 3284 53656 4724 53696
rect 4919 53656 4928 53696
rect 4968 53656 5010 53696
rect 5050 53656 5092 53696
rect 5132 53656 5174 53696
rect 5214 53656 5256 53696
rect 5296 53656 5305 53696
rect 5347 53656 5356 53696
rect 5396 53656 5452 53696
rect 5492 53656 5501 53696
rect 5827 53656 5836 53696
rect 5876 53656 6508 53696
rect 6548 53656 6557 53696
rect 11491 53656 11500 53696
rect 11540 53656 12460 53696
rect 12500 53656 12509 53696
rect 15619 53656 15628 53696
rect 15668 53656 15916 53696
rect 15956 53656 15965 53696
rect 0 53636 80 53656
rect 4684 53612 4724 53656
rect 5347 53655 5405 53656
rect 15907 53655 15965 53656
rect 9187 53612 9245 53613
rect 4675 53572 4684 53612
rect 4724 53572 6220 53612
rect 6260 53572 6269 53612
rect 7555 53572 7564 53612
rect 7604 53572 7756 53612
rect 7796 53572 7805 53612
rect 8899 53572 8908 53612
rect 8948 53572 9196 53612
rect 9236 53572 9245 53612
rect 9187 53571 9245 53572
rect 10531 53612 10589 53613
rect 16204 53612 16244 53740
rect 17251 53740 17260 53780
rect 17300 53740 20180 53780
rect 17251 53739 17309 53740
rect 17347 53696 17405 53697
rect 16387 53656 16396 53696
rect 16436 53656 16780 53696
rect 16820 53656 16829 53696
rect 17251 53656 17260 53696
rect 17300 53656 17356 53696
rect 17396 53656 17405 53696
rect 20039 53656 20048 53696
rect 20088 53656 20130 53696
rect 20170 53656 20212 53696
rect 20252 53656 20294 53696
rect 20334 53656 20376 53696
rect 20416 53656 20425 53696
rect 17347 53655 17405 53656
rect 19363 53612 19421 53613
rect 19843 53612 19901 53613
rect 10531 53572 10540 53612
rect 10580 53572 15436 53612
rect 15476 53572 16108 53612
rect 16148 53572 16157 53612
rect 16204 53572 19372 53612
rect 19412 53572 19421 53612
rect 19758 53572 19852 53612
rect 19892 53572 19901 53612
rect 10531 53571 10589 53572
rect 19363 53571 19421 53572
rect 19843 53571 19901 53572
rect 12931 53528 12989 53529
rect 21424 53528 21504 53548
rect 5539 53488 5548 53528
rect 5588 53488 6260 53528
rect 7459 53488 7468 53528
rect 7508 53488 8524 53528
rect 8564 53488 8573 53528
rect 8995 53488 9004 53528
rect 9044 53488 9292 53528
rect 9332 53488 9341 53528
rect 12739 53488 12748 53528
rect 12788 53488 12940 53528
rect 12980 53488 12989 53528
rect 13219 53488 13228 53528
rect 13268 53488 13420 53528
rect 13460 53488 13469 53528
rect 15235 53488 15244 53528
rect 15284 53488 16972 53528
rect 17012 53488 17021 53528
rect 17155 53488 17164 53528
rect 17204 53488 17740 53528
rect 17780 53488 17789 53528
rect 19459 53488 19468 53528
rect 19508 53488 21504 53528
rect 6220 53444 6260 53488
rect 12931 53487 12989 53488
rect 21424 53468 21504 53488
rect 21283 53444 21341 53445
rect 6211 53404 6220 53444
rect 6260 53404 6269 53444
rect 7651 53404 7660 53444
rect 7700 53404 13556 53444
rect 13603 53404 13612 53444
rect 13652 53404 21292 53444
rect 21332 53404 21341 53444
rect 3235 53360 3293 53361
rect 13516 53360 13556 53404
rect 21283 53403 21341 53404
rect 18019 53360 18077 53361
rect 1315 53320 1324 53360
rect 1364 53320 2188 53360
rect 2228 53320 2237 53360
rect 3150 53320 3244 53360
rect 3284 53320 3293 53360
rect 6499 53320 6508 53360
rect 6548 53320 7756 53360
rect 7796 53320 7805 53360
rect 8227 53320 8236 53360
rect 8276 53320 8620 53360
rect 8660 53320 8669 53360
rect 9379 53320 9388 53360
rect 9428 53320 9468 53360
rect 10147 53320 10156 53360
rect 10196 53320 10828 53360
rect 10868 53320 10877 53360
rect 11107 53320 11116 53360
rect 11156 53320 11692 53360
rect 11732 53320 11741 53360
rect 12643 53320 12652 53360
rect 12692 53320 13132 53360
rect 13172 53320 13181 53360
rect 13516 53320 14476 53360
rect 14516 53320 14525 53360
rect 15811 53320 15820 53360
rect 15860 53320 17068 53360
rect 17108 53320 17117 53360
rect 17934 53320 18028 53360
rect 18068 53320 18077 53360
rect 18403 53320 18412 53360
rect 18452 53320 18700 53360
rect 18740 53320 19276 53360
rect 19316 53320 19325 53360
rect 19372 53320 19660 53360
rect 19700 53320 19709 53360
rect 20227 53320 20236 53360
rect 20276 53320 20716 53360
rect 20756 53320 20765 53360
rect 3235 53319 3293 53320
rect 7267 53276 7325 53277
rect 9388 53276 9428 53320
rect 18019 53319 18077 53320
rect 10531 53276 10589 53277
rect 17443 53276 17501 53277
rect 7182 53236 7276 53276
rect 7316 53236 7325 53276
rect 7939 53236 7948 53276
rect 7988 53236 10252 53276
rect 10292 53236 10540 53276
rect 10580 53236 10589 53276
rect 11299 53236 11308 53276
rect 11348 53236 12460 53276
rect 12500 53236 12509 53276
rect 13219 53236 13228 53276
rect 13268 53236 17452 53276
rect 17492 53236 17501 53276
rect 7267 53235 7325 53236
rect 10531 53235 10589 53236
rect 11320 53192 11360 53236
rect 13228 53192 13268 53236
rect 17443 53235 17501 53236
rect 16291 53192 16349 53193
rect 2563 53152 2572 53192
rect 2612 53152 2956 53192
rect 2996 53152 3005 53192
rect 4387 53152 4396 53192
rect 4436 53152 11360 53192
rect 12931 53152 12940 53192
rect 12980 53152 13268 53192
rect 15715 53152 15724 53192
rect 15764 53152 16300 53192
rect 16340 53152 16349 53192
rect 16291 53151 16349 53152
rect 8131 53108 8189 53109
rect 11683 53108 11741 53109
rect 19372 53108 19412 53320
rect 19939 53192 19997 53193
rect 20131 53192 20189 53193
rect 21424 53192 21504 53212
rect 19459 53152 19468 53192
rect 19508 53152 19948 53192
rect 19988 53152 20084 53192
rect 19939 53151 19997 53152
rect 20044 53108 20084 53152
rect 20131 53152 20140 53192
rect 20180 53152 21504 53192
rect 20131 53151 20189 53152
rect 21424 53132 21504 53152
rect 8131 53068 8140 53108
rect 8180 53068 8332 53108
rect 8372 53068 8620 53108
rect 8660 53068 8669 53108
rect 8995 53068 9004 53108
rect 9044 53068 9676 53108
rect 9716 53068 9725 53108
rect 10531 53068 10540 53108
rect 10580 53068 10828 53108
rect 10868 53068 10877 53108
rect 11107 53068 11116 53108
rect 11156 53068 11692 53108
rect 11732 53068 11741 53108
rect 12355 53068 12364 53108
rect 12404 53068 16684 53108
rect 16724 53068 16733 53108
rect 17059 53068 17068 53108
rect 17108 53068 19412 53108
rect 19747 53068 19756 53108
rect 19796 53068 19805 53108
rect 20035 53068 20044 53108
rect 20084 53068 20093 53108
rect 8131 53067 8189 53068
rect 11683 53067 11741 53068
rect 0 53024 80 53044
rect 13027 53024 13085 53025
rect 18019 53024 18077 53025
rect 0 52984 9868 53024
rect 9908 52984 9917 53024
rect 13027 52984 13036 53024
rect 13076 52984 13132 53024
rect 13172 52984 13181 53024
rect 16579 52984 16588 53024
rect 16628 52984 16637 53024
rect 17731 52984 17740 53024
rect 17780 52984 18028 53024
rect 18068 52984 18077 53024
rect 0 52964 80 52984
rect 13027 52983 13085 52984
rect 10147 52940 10205 52941
rect 3679 52900 3688 52940
rect 3728 52900 3770 52940
rect 3810 52900 3852 52940
rect 3892 52900 3934 52940
rect 3974 52900 4016 52940
rect 4056 52900 4065 52940
rect 4396 52900 8140 52940
rect 8180 52900 8189 52940
rect 10062 52900 10156 52940
rect 10196 52900 10205 52940
rect 2563 52856 2621 52857
rect 4396 52856 4436 52900
rect 10147 52899 10205 52900
rect 10531 52940 10589 52941
rect 16588 52940 16628 52984
rect 18019 52983 18077 52984
rect 18691 53024 18749 53025
rect 18691 52984 18700 53024
rect 18740 52984 19564 53024
rect 19604 52984 19613 53024
rect 18691 52983 18749 52984
rect 10531 52900 10540 52940
rect 10580 52900 10732 52940
rect 10772 52900 10781 52940
rect 11971 52900 11980 52940
rect 12020 52900 12364 52940
rect 12404 52900 12413 52940
rect 12931 52900 12940 52940
rect 12980 52900 13228 52940
rect 13268 52900 13277 52940
rect 15811 52900 15820 52940
rect 15860 52900 16628 52940
rect 16675 52900 16684 52940
rect 16724 52900 18220 52940
rect 18260 52900 18269 52940
rect 18799 52900 18808 52940
rect 18848 52900 18890 52940
rect 18930 52900 18972 52940
rect 19012 52900 19054 52940
rect 19094 52900 19136 52940
rect 19176 52900 19185 52940
rect 10531 52899 10589 52900
rect 5923 52856 5981 52857
rect 16099 52856 16157 52857
rect 1507 52816 1516 52856
rect 1556 52816 2572 52856
rect 2612 52816 4436 52856
rect 4579 52816 4588 52856
rect 4628 52816 5452 52856
rect 5492 52816 5501 52856
rect 5838 52816 5932 52856
rect 5972 52816 5981 52856
rect 8035 52816 8044 52856
rect 8084 52816 11116 52856
rect 11156 52816 11165 52856
rect 11212 52816 13036 52856
rect 13076 52816 13085 52856
rect 16014 52816 16108 52856
rect 16148 52816 16876 52856
rect 16916 52816 17548 52856
rect 17588 52816 17597 52856
rect 18019 52816 18028 52856
rect 18068 52816 18700 52856
rect 18740 52816 18749 52856
rect 2563 52815 2621 52816
rect 5923 52815 5981 52816
rect 11212 52772 11252 52816
rect 16099 52815 16157 52816
rect 20 52732 2540 52772
rect 4195 52732 4204 52772
rect 4244 52732 8332 52772
rect 8372 52732 11252 52772
rect 11395 52772 11453 52773
rect 11395 52732 11404 52772
rect 11444 52732 14764 52772
rect 14804 52732 14813 52772
rect 18211 52732 18220 52772
rect 18260 52732 19660 52772
rect 19700 52732 19709 52772
rect 20 52520 60 52732
rect 2500 52688 2540 52732
rect 11395 52731 11453 52732
rect 19756 52688 19796 53068
rect 19852 52900 19948 52940
rect 19988 52900 19997 52940
rect 19852 52772 19892 52900
rect 19939 52856 19997 52857
rect 21424 52856 21504 52876
rect 19939 52816 19948 52856
rect 19988 52816 21504 52856
rect 19939 52815 19997 52816
rect 21424 52796 21504 52816
rect 19843 52732 19852 52772
rect 19892 52732 19901 52772
rect 2500 52648 4244 52688
rect 4291 52648 4300 52688
rect 4340 52648 6412 52688
rect 6452 52648 6461 52688
rect 6595 52648 6604 52688
rect 6644 52648 7180 52688
rect 7220 52648 7229 52688
rect 7747 52648 7756 52688
rect 7796 52648 10924 52688
rect 10964 52648 10973 52688
rect 11779 52648 11788 52688
rect 11828 52648 12556 52688
rect 12596 52648 12605 52688
rect 16483 52648 16492 52688
rect 16532 52648 16972 52688
rect 17012 52648 17021 52688
rect 17155 52648 17164 52688
rect 17204 52648 17548 52688
rect 17588 52648 17597 52688
rect 19756 52648 19948 52688
rect 19988 52648 19997 52688
rect 4204 52604 4244 52648
rect 14179 52604 14237 52605
rect 1411 52564 1420 52604
rect 1460 52564 2540 52604
rect 4204 52564 7084 52604
rect 7124 52564 8044 52604
rect 8084 52564 8093 52604
rect 10339 52564 10348 52604
rect 10388 52564 11828 52604
rect 12739 52564 12748 52604
rect 12788 52564 13713 52604
rect 13753 52564 13762 52604
rect 14179 52564 14188 52604
rect 14228 52564 19700 52604
rect 20131 52564 20140 52604
rect 20180 52564 20812 52604
rect 20852 52564 20861 52604
rect 2500 52520 2540 52564
rect 5539 52520 5597 52521
rect 11788 52520 11828 52564
rect 14179 52563 14237 52564
rect 19660 52520 19700 52564
rect 21424 52520 21504 52540
rect 20 52480 212 52520
rect 2500 52480 5548 52520
rect 5588 52480 5597 52520
rect 6883 52480 6892 52520
rect 6932 52480 6941 52520
rect 8707 52480 8716 52520
rect 8756 52480 10732 52520
rect 10772 52480 10781 52520
rect 10915 52480 10924 52520
rect 10964 52480 11252 52520
rect 11779 52480 11788 52520
rect 11828 52480 11837 52520
rect 13603 52480 13612 52520
rect 13652 52480 14188 52520
rect 14228 52480 14237 52520
rect 16579 52480 16588 52520
rect 16628 52480 17068 52520
rect 17108 52480 17117 52520
rect 18019 52480 18028 52520
rect 18068 52480 18796 52520
rect 18836 52480 18845 52520
rect 19651 52480 19660 52520
rect 19700 52480 19709 52520
rect 20428 52480 21504 52520
rect 0 52352 80 52372
rect 172 52352 212 52480
rect 5539 52479 5597 52480
rect 2275 52436 2333 52437
rect 6892 52436 6932 52480
rect 2275 52396 2284 52436
rect 2324 52396 6604 52436
rect 6644 52396 6653 52436
rect 6892 52396 7084 52436
rect 7124 52396 7133 52436
rect 9091 52396 9100 52436
rect 9140 52396 10156 52436
rect 10196 52396 11156 52436
rect 2275 52395 2333 52396
rect 8995 52352 9053 52353
rect 10915 52352 10973 52353
rect 11116 52352 11156 52396
rect 0 52312 212 52352
rect 2851 52312 2860 52352
rect 2900 52312 3532 52352
rect 3572 52312 3581 52352
rect 8227 52312 8236 52352
rect 8276 52312 9004 52352
rect 9044 52312 9580 52352
rect 9620 52312 9629 52352
rect 10243 52312 10252 52352
rect 10292 52312 10636 52352
rect 10676 52312 10685 52352
rect 10830 52312 10924 52352
rect 10964 52312 10973 52352
rect 11107 52312 11116 52352
rect 11156 52312 11165 52352
rect 0 52292 80 52312
rect 8995 52311 9053 52312
rect 10915 52311 10973 52312
rect 11212 52268 11252 52480
rect 11779 52436 11837 52437
rect 14563 52436 14621 52437
rect 19363 52436 19421 52437
rect 20428 52436 20468 52480
rect 21424 52460 21504 52480
rect 11779 52396 11788 52436
rect 11828 52396 13036 52436
rect 13076 52396 14572 52436
rect 14612 52396 14621 52436
rect 16483 52396 16492 52436
rect 16532 52396 18220 52436
rect 18260 52396 18269 52436
rect 19363 52396 19372 52436
rect 19412 52396 20468 52436
rect 11779 52395 11837 52396
rect 14563 52395 14621 52396
rect 19363 52395 19421 52396
rect 20803 52352 20861 52353
rect 12259 52312 12268 52352
rect 12308 52312 13324 52352
rect 13364 52312 13373 52352
rect 17923 52312 17932 52352
rect 17972 52312 18508 52352
rect 18548 52312 18557 52352
rect 20140 52312 20812 52352
rect 20852 52312 20861 52352
rect 20140 52268 20180 52312
rect 20803 52311 20861 52312
rect 10435 52228 10444 52268
rect 10484 52228 11020 52268
rect 11060 52228 11069 52268
rect 11212 52228 20180 52268
rect 16867 52184 16925 52185
rect 20 52144 4204 52184
rect 4244 52144 4253 52184
rect 4919 52144 4928 52184
rect 4968 52144 5010 52184
rect 5050 52144 5092 52184
rect 5132 52144 5174 52184
rect 5214 52144 5256 52184
rect 5296 52144 5305 52184
rect 5347 52144 5356 52184
rect 5396 52144 5644 52184
rect 5684 52144 5693 52184
rect 12931 52144 12940 52184
rect 12980 52144 13516 52184
rect 13556 52144 13565 52184
rect 14275 52144 14284 52184
rect 14324 52144 16532 52184
rect 16782 52144 16876 52184
rect 16916 52144 16925 52184
rect 20 51848 60 52144
rect 3043 52100 3101 52101
rect 10531 52100 10589 52101
rect 16291 52100 16349 52101
rect 3043 52060 3052 52100
rect 3092 52060 7756 52100
rect 7796 52060 7805 52100
rect 10531 52060 10540 52100
rect 10580 52060 10636 52100
rect 10676 52060 10685 52100
rect 11875 52060 11884 52100
rect 11924 52060 12460 52100
rect 12500 52060 13556 52100
rect 15907 52060 15916 52100
rect 15956 52060 15965 52100
rect 16206 52060 16300 52100
rect 16340 52060 16349 52100
rect 3043 52059 3101 52060
rect 10531 52059 10589 52060
rect 13123 52016 13181 52017
rect 13516 52016 13556 52060
rect 15916 52016 15956 52060
rect 16291 52059 16349 52060
rect 16492 52016 16532 52144
rect 16867 52143 16925 52144
rect 17923 52184 17981 52185
rect 19939 52184 19997 52185
rect 21424 52184 21504 52204
rect 17923 52144 17932 52184
rect 17972 52144 19948 52184
rect 19988 52144 19997 52184
rect 20039 52144 20048 52184
rect 20088 52144 20130 52184
rect 20170 52144 20212 52184
rect 20252 52144 20294 52184
rect 20334 52144 20376 52184
rect 20416 52144 20425 52184
rect 20524 52144 21504 52184
rect 17923 52143 17981 52144
rect 19939 52143 19997 52144
rect 20524 52100 20564 52144
rect 21424 52124 21504 52144
rect 16675 52060 16684 52100
rect 16724 52060 20564 52100
rect 19651 52016 19709 52017
rect 5443 51976 5452 52016
rect 5492 51976 6412 52016
rect 6452 51976 6461 52016
rect 7171 51976 7180 52016
rect 7220 51976 7260 52016
rect 13027 51976 13036 52016
rect 13076 51976 13132 52016
rect 13172 51976 13181 52016
rect 13507 51976 13516 52016
rect 13556 51976 13565 52016
rect 15916 51976 16396 52016
rect 16436 51976 16445 52016
rect 16492 51976 19660 52016
rect 19700 51976 19709 52016
rect 7180 51932 7220 51976
rect 13123 51975 13181 51976
rect 19651 51975 19709 51976
rect 5347 51892 5356 51932
rect 5396 51892 10444 51932
rect 10484 51892 10493 51932
rect 11500 51892 15572 51932
rect 15907 51892 15916 51932
rect 15956 51892 16780 51932
rect 16820 51892 16829 51932
rect 17548 51892 18700 51932
rect 18740 51892 18749 51932
rect 3427 51848 3485 51849
rect 4291 51848 4349 51849
rect 11500 51848 11540 51892
rect 15532 51848 15572 51892
rect 17548 51848 17588 51892
rect 20 51808 212 51848
rect 1411 51808 1420 51848
rect 1460 51808 1996 51848
rect 2036 51808 2045 51848
rect 2851 51808 2860 51848
rect 2900 51808 3244 51848
rect 3284 51808 3293 51848
rect 3427 51808 3436 51848
rect 3476 51808 3724 51848
rect 3764 51808 3773 51848
rect 4206 51808 4300 51848
rect 4340 51808 4349 51848
rect 6115 51808 6124 51848
rect 6164 51808 7180 51848
rect 7220 51808 7229 51848
rect 8323 51808 8332 51848
rect 8372 51808 8381 51848
rect 9859 51808 9868 51848
rect 9908 51808 11500 51848
rect 11540 51808 11549 51848
rect 12547 51808 12556 51848
rect 12596 51808 12748 51848
rect 12788 51808 15148 51848
rect 15188 51808 15197 51848
rect 15532 51808 17588 51848
rect 17635 51848 17693 51849
rect 21424 51848 21504 51868
rect 17635 51808 17644 51848
rect 17684 51808 21504 51848
rect 0 51680 80 51700
rect 172 51680 212 51808
rect 3427 51807 3485 51808
rect 4291 51807 4349 51808
rect 8332 51764 8372 51808
rect 17635 51807 17693 51808
rect 21424 51788 21504 51808
rect 3043 51724 3052 51764
rect 3092 51724 3916 51764
rect 3956 51724 3965 51764
rect 6220 51724 8372 51764
rect 12835 51764 12893 51765
rect 14851 51764 14909 51765
rect 12835 51724 12844 51764
rect 12884 51724 14668 51764
rect 14708 51724 14717 51764
rect 14851 51724 14860 51764
rect 14900 51724 14994 51764
rect 16291 51724 16300 51764
rect 16340 51724 16916 51764
rect 17059 51724 17068 51764
rect 17108 51724 17356 51764
rect 17396 51724 17740 51764
rect 17780 51724 17789 51764
rect 18307 51724 18316 51764
rect 18356 51724 18604 51764
rect 18644 51724 18653 51764
rect 5443 51680 5501 51681
rect 6220 51680 6260 51724
rect 12835 51723 12893 51724
rect 14851 51723 14909 51724
rect 16099 51680 16157 51681
rect 16876 51680 16916 51724
rect 18019 51680 18077 51681
rect 19267 51680 19325 51681
rect 0 51640 212 51680
rect 2851 51640 2860 51680
rect 2900 51640 3340 51680
rect 3380 51640 3389 51680
rect 5443 51640 5452 51680
rect 5492 51640 5932 51680
rect 5972 51640 5981 51680
rect 6211 51640 6220 51680
rect 6260 51640 6269 51680
rect 7363 51640 7372 51680
rect 7412 51640 9196 51680
rect 9236 51640 9245 51680
rect 14179 51640 14188 51680
rect 14228 51640 15532 51680
rect 15572 51640 15581 51680
rect 16099 51640 16108 51680
rect 16148 51640 16204 51680
rect 16244 51640 16253 51680
rect 16387 51640 16396 51680
rect 16436 51640 16820 51680
rect 16876 51640 17548 51680
rect 17588 51640 17597 51680
rect 18019 51640 18028 51680
rect 18068 51640 18220 51680
rect 18260 51640 18269 51680
rect 18403 51640 18412 51680
rect 18452 51640 19276 51680
rect 19316 51640 19325 51680
rect 0 51620 80 51640
rect 5443 51639 5501 51640
rect 5539 51596 5597 51597
rect 10723 51596 10781 51597
rect 5539 51556 5548 51596
rect 5588 51556 5644 51596
rect 5684 51556 5693 51596
rect 7843 51556 7852 51596
rect 7892 51556 8524 51596
rect 8564 51556 8573 51596
rect 10723 51556 10732 51596
rect 10772 51556 13036 51596
rect 13076 51556 13085 51596
rect 5539 51555 5597 51556
rect 10723 51555 10781 51556
rect 13027 51512 13085 51513
rect 15532 51512 15572 51640
rect 16099 51639 16157 51640
rect 16291 51596 16349 51597
rect 16780 51596 16820 51640
rect 18019 51639 18077 51640
rect 19267 51639 19325 51640
rect 17251 51596 17309 51597
rect 16206 51556 16300 51596
rect 16340 51556 16349 51596
rect 16771 51556 16780 51596
rect 16820 51556 16829 51596
rect 17166 51556 17260 51596
rect 17300 51556 17309 51596
rect 18595 51556 18604 51596
rect 18644 51556 20140 51596
rect 20180 51556 20189 51596
rect 16291 51555 16349 51556
rect 17251 51555 17309 51556
rect 21424 51512 21504 51532
rect 13027 51472 13036 51512
rect 13076 51472 13804 51512
rect 13844 51472 13853 51512
rect 15532 51472 17164 51512
rect 17204 51472 17213 51512
rect 20899 51472 20908 51512
rect 20948 51472 21504 51512
rect 13027 51471 13085 51472
rect 21424 51452 21504 51472
rect 11587 51428 11645 51429
rect 3679 51388 3688 51428
rect 3728 51388 3770 51428
rect 3810 51388 3852 51428
rect 3892 51388 3934 51428
rect 3974 51388 4016 51428
rect 4056 51388 4065 51428
rect 11587 51388 11596 51428
rect 11636 51388 15532 51428
rect 15572 51388 15581 51428
rect 18799 51388 18808 51428
rect 18848 51388 18890 51428
rect 18930 51388 18972 51428
rect 19012 51388 19054 51428
rect 19094 51388 19136 51428
rect 19176 51388 19185 51428
rect 11587 51387 11645 51388
rect 7267 51344 7325 51345
rect 2467 51304 2476 51344
rect 2516 51304 4876 51344
rect 4916 51304 5932 51344
rect 5972 51304 7084 51344
rect 7124 51304 7133 51344
rect 7267 51304 7276 51344
rect 7316 51304 7948 51344
rect 7988 51304 7997 51344
rect 8611 51304 8620 51344
rect 8660 51304 21196 51344
rect 21236 51304 21245 51344
rect 7267 51303 7325 51304
rect 3139 51260 3197 51261
rect 7651 51260 7709 51261
rect 8035 51260 8093 51261
rect 3139 51220 3148 51260
rect 3188 51220 3628 51260
rect 3668 51220 3677 51260
rect 7555 51220 7564 51260
rect 7604 51220 7660 51260
rect 7700 51220 7709 51260
rect 7950 51220 8044 51260
rect 8084 51220 8093 51260
rect 3139 51219 3197 51220
rect 7651 51219 7709 51220
rect 8035 51219 8093 51220
rect 8323 51260 8381 51261
rect 8323 51220 8332 51260
rect 8372 51220 16396 51260
rect 16436 51220 16445 51260
rect 18883 51220 18892 51260
rect 18932 51220 19948 51260
rect 19988 51220 19997 51260
rect 8323 51219 8381 51220
rect 7843 51176 7901 51177
rect 7651 51136 7660 51176
rect 7700 51136 7852 51176
rect 7892 51136 7901 51176
rect 7843 51135 7901 51136
rect 8515 51176 8573 51177
rect 21424 51176 21504 51196
rect 8515 51136 8524 51176
rect 8564 51136 8620 51176
rect 8660 51136 8669 51176
rect 12259 51136 12268 51176
rect 12308 51136 14092 51176
rect 14132 51136 14141 51176
rect 17443 51136 17452 51176
rect 17492 51136 18028 51176
rect 18068 51136 18077 51176
rect 18124 51136 21504 51176
rect 8515 51135 8573 51136
rect 16099 51092 16157 51093
rect 18124 51092 18164 51136
rect 21424 51116 21504 51136
rect 2755 51052 2764 51092
rect 2804 51052 3340 51092
rect 3380 51052 4012 51092
rect 4052 51052 4780 51092
rect 4820 51052 4829 51092
rect 7372 51052 9292 51092
rect 9332 51052 9341 51092
rect 13411 51052 13420 51092
rect 13460 51052 13469 51092
rect 16099 51052 16108 51092
rect 16148 51052 18164 51092
rect 19555 51052 19564 51092
rect 19604 51052 20812 51092
rect 20852 51052 20861 51092
rect 0 51008 80 51028
rect 7372 51008 7412 51052
rect 0 50968 2540 51008
rect 2851 50968 2860 51008
rect 2900 50968 3916 51008
rect 3956 50968 3965 51008
rect 4099 50968 4108 51008
rect 4148 50968 7412 51008
rect 7459 50968 7468 51008
rect 7508 50968 9100 51008
rect 9140 50968 9149 51008
rect 0 50948 80 50968
rect 2500 50924 2540 50968
rect 1315 50884 1324 50924
rect 1364 50884 2092 50924
rect 2132 50884 2141 50924
rect 2500 50884 4300 50924
rect 4340 50884 6316 50924
rect 6356 50884 6365 50924
rect 7747 50884 7756 50924
rect 7796 50884 8044 50924
rect 8084 50884 8093 50924
rect 8323 50884 8332 50924
rect 8372 50884 13268 50924
rect 8035 50840 8093 50841
rect 9763 50840 9821 50841
rect 2659 50800 2668 50840
rect 2708 50800 4396 50840
rect 4436 50800 4445 50840
rect 8035 50800 8044 50840
rect 8084 50800 8236 50840
rect 8276 50800 8285 50840
rect 9678 50800 9772 50840
rect 9812 50800 9821 50840
rect 8035 50799 8093 50800
rect 9763 50799 9821 50800
rect 8323 50756 8381 50757
rect 12163 50756 12221 50757
rect 2275 50716 2284 50756
rect 2324 50716 4684 50756
rect 4724 50716 8332 50756
rect 8372 50716 8381 50756
rect 9187 50716 9196 50756
rect 9236 50716 12172 50756
rect 12212 50716 12221 50756
rect 8323 50715 8381 50716
rect 12163 50715 12221 50716
rect 13228 50672 13268 50884
rect 13420 50840 13460 51052
rect 16099 51051 16157 51052
rect 19267 51008 19325 51009
rect 13699 50968 13708 51008
rect 13748 50968 14092 51008
rect 14132 50968 14572 51008
rect 14612 50968 14621 51008
rect 16675 50968 16684 51008
rect 16724 50968 17644 51008
rect 17684 50968 17693 51008
rect 19075 50968 19084 51008
rect 19124 50968 19276 51008
rect 19316 50968 19372 51008
rect 19412 50968 19440 51008
rect 19267 50967 19325 50968
rect 19843 50924 19901 50925
rect 19843 50884 19852 50924
rect 19892 50884 20276 50924
rect 19843 50883 19901 50884
rect 17059 50840 17117 50841
rect 19939 50840 19997 50841
rect 20236 50840 20276 50884
rect 21424 50840 21504 50860
rect 13420 50800 13708 50840
rect 13748 50800 13757 50840
rect 13891 50800 13900 50840
rect 13940 50800 14572 50840
rect 14612 50800 14621 50840
rect 17059 50800 17068 50840
rect 17108 50800 17836 50840
rect 17876 50800 17885 50840
rect 19939 50800 19948 50840
rect 19988 50800 20140 50840
rect 20180 50800 20189 50840
rect 20236 50800 21504 50840
rect 17059 50799 17117 50800
rect 19939 50799 19997 50800
rect 21424 50780 21504 50800
rect 15619 50716 15628 50756
rect 15668 50716 17644 50756
rect 17684 50716 17693 50756
rect 15715 50672 15773 50673
rect 19843 50672 19901 50673
rect 4919 50632 4928 50672
rect 4968 50632 5010 50672
rect 5050 50632 5092 50672
rect 5132 50632 5174 50672
rect 5214 50632 5256 50672
rect 5296 50632 5305 50672
rect 6883 50632 6892 50672
rect 6932 50632 7660 50672
rect 7700 50632 7709 50672
rect 13228 50632 15148 50672
rect 15188 50632 15197 50672
rect 15630 50632 15724 50672
rect 15764 50632 15773 50672
rect 16963 50632 16972 50672
rect 17012 50632 18220 50672
rect 18260 50632 18269 50672
rect 19843 50632 19852 50672
rect 19892 50632 19948 50672
rect 19988 50632 19997 50672
rect 20039 50632 20048 50672
rect 20088 50632 20130 50672
rect 20170 50632 20212 50672
rect 20252 50632 20294 50672
rect 20334 50632 20376 50672
rect 20416 50632 20425 50672
rect 7075 50548 7084 50588
rect 7124 50548 7468 50588
rect 7508 50548 7517 50588
rect 7660 50504 7700 50632
rect 15715 50631 15773 50632
rect 19843 50631 19901 50632
rect 13219 50588 13277 50589
rect 13134 50548 13228 50588
rect 13268 50548 13277 50588
rect 14467 50548 14476 50588
rect 14516 50548 20180 50588
rect 13219 50547 13277 50548
rect 20140 50504 20180 50548
rect 21424 50504 21504 50524
rect 7660 50464 8084 50504
rect 8227 50464 8236 50504
rect 8276 50464 11404 50504
rect 11444 50464 15532 50504
rect 15572 50464 15581 50504
rect 15715 50464 15724 50504
rect 15764 50464 17356 50504
rect 17396 50464 17405 50504
rect 17539 50464 17548 50504
rect 17588 50464 17597 50504
rect 20140 50464 21504 50504
rect 8044 50420 8084 50464
rect 8995 50420 9053 50421
rect 17548 50420 17588 50464
rect 21424 50444 21504 50464
rect 19939 50420 19997 50421
rect 6499 50380 6508 50420
rect 6548 50380 7948 50420
rect 7988 50380 7997 50420
rect 8044 50380 9004 50420
rect 9044 50380 9484 50420
rect 9524 50380 9533 50420
rect 12643 50380 12652 50420
rect 12692 50380 14764 50420
rect 14804 50380 14813 50420
rect 15427 50380 15436 50420
rect 15476 50380 17588 50420
rect 18979 50380 18988 50420
rect 19028 50380 19948 50420
rect 19988 50380 19997 50420
rect 8995 50379 9053 50380
rect 19939 50379 19997 50380
rect 0 50336 80 50356
rect 4291 50336 4349 50337
rect 4483 50336 4541 50337
rect 0 50296 1708 50336
rect 1748 50296 1757 50336
rect 3811 50296 3820 50336
rect 3860 50296 4300 50336
rect 4340 50296 4492 50336
rect 4532 50296 4541 50336
rect 6019 50296 6028 50336
rect 6068 50296 7700 50336
rect 0 50276 80 50296
rect 4291 50295 4349 50296
rect 4483 50295 4541 50296
rect 3139 50252 3197 50253
rect 7660 50252 7700 50296
rect 8332 50296 11212 50336
rect 11252 50296 12172 50336
rect 12212 50296 12364 50336
rect 12404 50296 12413 50336
rect 15619 50296 15628 50336
rect 15668 50296 16204 50336
rect 16244 50296 17356 50336
rect 17396 50296 17405 50336
rect 18403 50296 18412 50336
rect 18452 50296 19180 50336
rect 19220 50296 19229 50336
rect 19363 50296 19372 50336
rect 19412 50296 20140 50336
rect 20180 50296 20189 50336
rect 1411 50212 1420 50252
rect 1460 50212 3148 50252
rect 3188 50212 3197 50252
rect 7651 50212 7660 50252
rect 7700 50212 7709 50252
rect 3139 50211 3197 50212
rect 8332 50168 8372 50296
rect 9475 50212 9484 50252
rect 9524 50212 11116 50252
rect 11156 50212 13036 50252
rect 13076 50212 13085 50252
rect 16387 50212 16396 50252
rect 16436 50212 16972 50252
rect 17012 50212 17021 50252
rect 17644 50212 20236 50252
rect 20276 50212 20620 50252
rect 20660 50212 20669 50252
rect 17644 50168 17684 50212
rect 20803 50168 20861 50169
rect 21424 50168 21504 50188
rect 1603 50128 1612 50168
rect 1652 50128 8372 50168
rect 8428 50128 15532 50168
rect 15572 50128 15581 50168
rect 17635 50128 17644 50168
rect 17684 50128 17693 50168
rect 18115 50128 18124 50168
rect 18164 50128 18796 50168
rect 18836 50128 18845 50168
rect 19363 50128 19372 50168
rect 19412 50128 19756 50168
rect 19796 50128 19805 50168
rect 20803 50128 20812 50168
rect 20852 50128 21504 50168
rect 2371 50044 2380 50084
rect 2420 50044 2860 50084
rect 2900 50044 2909 50084
rect 3235 50044 3244 50084
rect 3284 50044 4012 50084
rect 4052 50044 4061 50084
rect 5731 50044 5740 50084
rect 5780 50044 6028 50084
rect 6068 50044 6077 50084
rect 3139 50000 3197 50001
rect 5827 50000 5885 50001
rect 8428 50000 8468 50128
rect 20803 50127 20861 50128
rect 21424 50108 21504 50128
rect 12163 50084 12221 50085
rect 19651 50084 19709 50085
rect 12163 50044 12172 50084
rect 12212 50044 14956 50084
rect 14996 50044 15005 50084
rect 19566 50044 19660 50084
rect 19700 50044 19709 50084
rect 12163 50043 12221 50044
rect 19651 50043 19709 50044
rect 3139 49960 3148 50000
rect 3188 49960 4588 50000
rect 4628 49960 4637 50000
rect 5827 49960 5836 50000
rect 5876 49960 8468 50000
rect 8611 49960 8620 50000
rect 8660 49960 20524 50000
rect 20564 49960 20573 50000
rect 3139 49959 3197 49960
rect 5827 49959 5885 49960
rect 3679 49876 3688 49916
rect 3728 49876 3770 49916
rect 3810 49876 3852 49916
rect 3892 49876 3934 49916
rect 3974 49876 4016 49916
rect 4056 49876 4065 49916
rect 5827 49876 5836 49916
rect 5876 49876 6124 49916
rect 6164 49876 6173 49916
rect 13411 49876 13420 49916
rect 13460 49876 14092 49916
rect 14132 49876 16396 49916
rect 16436 49876 16445 49916
rect 18799 49876 18808 49916
rect 18848 49876 18890 49916
rect 18930 49876 18972 49916
rect 19012 49876 19054 49916
rect 19094 49876 19136 49916
rect 19176 49876 19185 49916
rect 19363 49876 19372 49916
rect 19412 49876 19660 49916
rect 19700 49876 19709 49916
rect 7363 49832 7421 49833
rect 19555 49832 19613 49833
rect 21424 49832 21504 49852
rect 7363 49792 7372 49832
rect 7412 49792 8236 49832
rect 8276 49792 8285 49832
rect 10147 49792 10156 49832
rect 10196 49792 19564 49832
rect 19604 49792 19613 49832
rect 20611 49792 20620 49832
rect 20660 49792 21504 49832
rect 7363 49791 7421 49792
rect 19555 49791 19613 49792
rect 21424 49772 21504 49792
rect 5347 49748 5405 49749
rect 5827 49748 5885 49749
rect 15331 49748 15389 49749
rect 5347 49708 5356 49748
rect 5396 49708 5836 49748
rect 5876 49708 5885 49748
rect 7075 49708 7084 49748
rect 7124 49708 7852 49748
rect 7892 49708 7901 49748
rect 14371 49708 14380 49748
rect 14420 49708 14764 49748
rect 14804 49708 14813 49748
rect 15235 49708 15244 49748
rect 15284 49708 15340 49748
rect 15380 49708 15389 49748
rect 5347 49707 5405 49708
rect 5827 49707 5885 49708
rect 15331 49707 15389 49708
rect 0 49664 80 49684
rect 7651 49664 7709 49665
rect 0 49624 1420 49664
rect 1460 49624 1469 49664
rect 3811 49624 3820 49664
rect 3860 49624 4204 49664
rect 4244 49624 4253 49664
rect 5443 49624 5452 49664
rect 5492 49624 7660 49664
rect 7700 49624 7709 49664
rect 0 49604 80 49624
rect 7651 49623 7709 49624
rect 8323 49664 8381 49665
rect 8323 49624 8332 49664
rect 8372 49624 8428 49664
rect 8468 49624 8477 49664
rect 11779 49624 11788 49664
rect 11828 49624 12940 49664
rect 12980 49624 12989 49664
rect 13891 49624 13900 49664
rect 13940 49624 17644 49664
rect 17684 49624 17693 49664
rect 8323 49623 8381 49624
rect 4579 49580 4637 49581
rect 3907 49540 3916 49580
rect 3956 49540 4588 49580
rect 4628 49540 10156 49580
rect 10196 49540 10205 49580
rect 12835 49540 12844 49580
rect 12884 49540 12980 49580
rect 14371 49540 14380 49580
rect 14420 49540 14668 49580
rect 14708 49540 14717 49580
rect 15043 49540 15052 49580
rect 15092 49540 17452 49580
rect 17492 49540 17501 49580
rect 18115 49540 18124 49580
rect 18164 49540 19892 49580
rect 4579 49539 4637 49540
rect 12940 49496 12980 49540
rect 18307 49496 18365 49497
rect 19852 49496 19892 49540
rect 21424 49496 21504 49516
rect 4291 49456 4300 49496
rect 4340 49456 5836 49496
rect 5876 49456 5885 49496
rect 6307 49456 6316 49496
rect 6356 49456 8428 49496
rect 8468 49456 8477 49496
rect 12931 49456 12940 49496
rect 12980 49456 12989 49496
rect 13123 49456 13132 49496
rect 13172 49456 14476 49496
rect 14516 49456 14525 49496
rect 15235 49456 15244 49496
rect 15284 49456 17164 49496
rect 17204 49456 17213 49496
rect 18307 49456 18316 49496
rect 18356 49456 18604 49496
rect 18644 49456 18653 49496
rect 19843 49456 19852 49496
rect 19892 49456 19901 49496
rect 20140 49456 21504 49496
rect 18307 49455 18365 49456
rect 2083 49412 2141 49413
rect 4099 49412 4157 49413
rect 4771 49412 4829 49413
rect 11491 49412 11549 49413
rect 20140 49412 20180 49456
rect 21424 49436 21504 49456
rect 2083 49372 2092 49412
rect 2132 49372 2668 49412
rect 2708 49372 2717 49412
rect 4099 49372 4108 49412
rect 4148 49372 4780 49412
rect 4820 49372 4972 49412
rect 5012 49372 5021 49412
rect 6115 49372 6124 49412
rect 6164 49372 6892 49412
rect 6932 49372 6941 49412
rect 11299 49372 11308 49412
rect 11348 49372 11500 49412
rect 11540 49372 11549 49412
rect 13987 49372 13996 49412
rect 14036 49372 14188 49412
rect 14228 49372 20180 49412
rect 2083 49371 2141 49372
rect 4099 49371 4157 49372
rect 4771 49371 4829 49372
rect 11491 49371 11549 49372
rect 10147 49328 10205 49329
rect 19939 49328 19997 49329
rect 2851 49288 2860 49328
rect 2900 49288 4684 49328
rect 4724 49288 4733 49328
rect 7459 49288 7468 49328
rect 7508 49288 9292 49328
rect 9332 49288 9341 49328
rect 10147 49288 10156 49328
rect 10196 49288 10636 49328
rect 10676 49288 10685 49328
rect 18019 49288 18028 49328
rect 18068 49288 18412 49328
rect 18452 49288 18461 49328
rect 19939 49288 19948 49328
rect 19988 49288 20044 49328
rect 20084 49288 20093 49328
rect 10147 49287 10205 49288
rect 19939 49287 19997 49288
rect 5923 49244 5981 49245
rect 4291 49204 4300 49244
rect 4340 49204 5932 49244
rect 5972 49204 6508 49244
rect 6548 49204 6557 49244
rect 15331 49204 15340 49244
rect 15380 49204 15628 49244
rect 15668 49204 15677 49244
rect 16003 49204 16012 49244
rect 16052 49204 16396 49244
rect 16436 49204 16972 49244
rect 17012 49204 17548 49244
rect 17588 49204 17597 49244
rect 5923 49203 5981 49204
rect 21424 49160 21504 49180
rect 3436 49120 4780 49160
rect 4820 49120 4829 49160
rect 4919 49120 4928 49160
rect 4968 49120 5010 49160
rect 5050 49120 5092 49160
rect 5132 49120 5174 49160
rect 5214 49120 5256 49160
rect 5296 49120 5305 49160
rect 11107 49120 11116 49160
rect 11156 49120 11596 49160
rect 11636 49120 11645 49160
rect 15523 49120 15532 49160
rect 15572 49120 17356 49160
rect 17396 49120 17405 49160
rect 20039 49120 20048 49160
rect 20088 49120 20130 49160
rect 20170 49120 20212 49160
rect 20252 49120 20294 49160
rect 20334 49120 20376 49160
rect 20416 49120 20425 49160
rect 20515 49120 20524 49160
rect 20564 49120 21504 49160
rect 0 48992 80 49012
rect 0 48952 1324 48992
rect 1364 48952 1516 48992
rect 1556 48952 1565 48992
rect 3043 48952 3052 48992
rect 3092 48952 3340 48992
rect 3380 48952 3389 48992
rect 0 48932 80 48952
rect 2563 48740 2621 48741
rect 2563 48700 2572 48740
rect 2612 48700 2764 48740
rect 2804 48700 2813 48740
rect 2563 48699 2621 48700
rect 3436 48656 3476 49120
rect 21424 49100 21504 49120
rect 6211 49036 6220 49076
rect 6260 49036 20180 49076
rect 17923 48992 17981 48993
rect 4867 48952 4876 48992
rect 4916 48952 17932 48992
rect 17972 48952 17981 48992
rect 18499 48952 18508 48992
rect 18548 48952 19852 48992
rect 19892 48952 19901 48992
rect 17923 48951 17981 48952
rect 11491 48908 11549 48909
rect 19363 48908 19421 48909
rect 4771 48868 4780 48908
rect 4820 48868 5452 48908
rect 5492 48868 5501 48908
rect 6307 48868 6316 48908
rect 6356 48868 6988 48908
rect 7028 48868 7037 48908
rect 11406 48868 11500 48908
rect 11540 48868 11549 48908
rect 16291 48868 16300 48908
rect 16340 48868 18892 48908
rect 18932 48868 18941 48908
rect 19075 48868 19084 48908
rect 19124 48868 19372 48908
rect 19412 48868 19421 48908
rect 20140 48908 20180 49036
rect 20803 48908 20861 48909
rect 20140 48868 20812 48908
rect 20852 48868 20861 48908
rect 11491 48867 11549 48868
rect 19363 48867 19421 48868
rect 20803 48867 20861 48868
rect 21424 48824 21504 48844
rect 5251 48784 5260 48824
rect 5300 48784 6220 48824
rect 6260 48784 6269 48824
rect 6499 48784 6508 48824
rect 6548 48784 6796 48824
rect 6836 48784 6845 48824
rect 7267 48784 7276 48824
rect 7316 48784 7948 48824
rect 7988 48784 7997 48824
rect 10051 48784 10060 48824
rect 10100 48784 10252 48824
rect 10292 48784 21504 48824
rect 7564 48740 7604 48784
rect 21424 48764 21504 48784
rect 4099 48700 4108 48740
rect 4148 48700 4157 48740
rect 7555 48700 7564 48740
rect 7604 48700 7644 48740
rect 13411 48700 13420 48740
rect 13460 48700 13900 48740
rect 13940 48700 13949 48740
rect 13996 48700 14956 48740
rect 14996 48700 15005 48740
rect 19459 48700 19468 48740
rect 19508 48700 20180 48740
rect 4108 48656 4148 48700
rect 13996 48656 14036 48700
rect 16483 48656 16541 48657
rect 20140 48656 20180 48700
rect 3427 48616 3436 48656
rect 3476 48616 3485 48656
rect 3619 48616 3628 48656
rect 3668 48616 7468 48656
rect 7508 48616 7517 48656
rect 7651 48616 7660 48656
rect 7700 48616 8236 48656
rect 8276 48616 8285 48656
rect 12931 48616 12940 48656
rect 12980 48616 14036 48656
rect 14179 48616 14188 48656
rect 14228 48616 16492 48656
rect 16532 48616 16541 48656
rect 16771 48616 16780 48656
rect 16820 48616 17548 48656
rect 17588 48616 17597 48656
rect 18691 48616 18700 48656
rect 18740 48616 20044 48656
rect 20084 48616 20093 48656
rect 20140 48616 20620 48656
rect 20660 48616 20669 48656
rect 16483 48615 16541 48616
rect 12547 48572 12605 48573
rect 2755 48532 2764 48572
rect 2804 48532 3148 48572
rect 3188 48532 4588 48572
rect 4628 48532 5356 48572
rect 5396 48532 5405 48572
rect 6508 48532 8044 48572
rect 8084 48532 8620 48572
rect 8660 48532 11692 48572
rect 11732 48532 11741 48572
rect 12547 48532 12556 48572
rect 12596 48532 19852 48572
rect 19892 48532 19901 48572
rect 2851 48488 2909 48489
rect 6508 48488 6548 48532
rect 12547 48531 12605 48532
rect 2851 48448 2860 48488
rect 2900 48448 6548 48488
rect 6595 48488 6653 48489
rect 12835 48488 12893 48489
rect 16483 48488 16541 48489
rect 21283 48488 21341 48489
rect 21424 48488 21504 48508
rect 6595 48448 6604 48488
rect 6644 48448 11884 48488
rect 11924 48448 12844 48488
rect 12884 48448 12893 48488
rect 15043 48448 15052 48488
rect 15092 48448 16300 48488
rect 16340 48448 16349 48488
rect 16483 48448 16492 48488
rect 16532 48448 18508 48488
rect 18548 48448 18557 48488
rect 21283 48448 21292 48488
rect 21332 48448 21504 48488
rect 2851 48447 2909 48448
rect 6595 48447 6653 48448
rect 12835 48447 12893 48448
rect 16483 48447 16541 48448
rect 21283 48447 21341 48448
rect 5923 48404 5981 48405
rect 6604 48404 6644 48447
rect 21424 48428 21504 48448
rect 8515 48404 8573 48405
rect 2947 48364 2956 48404
rect 2996 48364 3148 48404
rect 3188 48364 3197 48404
rect 3679 48364 3688 48404
rect 3728 48364 3770 48404
rect 3810 48364 3852 48404
rect 3892 48364 3934 48404
rect 3974 48364 4016 48404
rect 4056 48364 4065 48404
rect 5347 48364 5356 48404
rect 5396 48364 5932 48404
rect 5972 48364 6644 48404
rect 7459 48364 7468 48404
rect 7508 48364 8524 48404
rect 8564 48364 8573 48404
rect 5923 48363 5981 48364
rect 8515 48363 8573 48364
rect 14851 48404 14909 48405
rect 14851 48364 14860 48404
rect 14900 48364 18604 48404
rect 18644 48364 18653 48404
rect 18799 48364 18808 48404
rect 18848 48364 18890 48404
rect 18930 48364 18972 48404
rect 19012 48364 19054 48404
rect 19094 48364 19136 48404
rect 19176 48364 19185 48404
rect 14851 48363 14909 48364
rect 0 48320 80 48340
rect 0 48280 2284 48320
rect 2324 48280 2333 48320
rect 11491 48280 11500 48320
rect 11540 48280 12172 48320
rect 12212 48280 12460 48320
rect 12500 48280 12509 48320
rect 16675 48280 16684 48320
rect 16724 48280 17452 48320
rect 17492 48280 17501 48320
rect 18316 48280 19468 48320
rect 19508 48280 19517 48320
rect 0 48260 80 48280
rect 2851 48236 2909 48237
rect 18316 48236 18356 48280
rect 1315 48196 1324 48236
rect 1364 48196 2860 48236
rect 2900 48196 2909 48236
rect 3811 48196 3820 48236
rect 3860 48196 4204 48236
rect 4244 48196 6988 48236
rect 7028 48196 7037 48236
rect 10243 48196 10252 48236
rect 10292 48196 14284 48236
rect 14324 48196 14333 48236
rect 15907 48196 15916 48236
rect 15956 48196 18356 48236
rect 18403 48196 18412 48236
rect 18452 48196 19564 48236
rect 19604 48196 19613 48236
rect 2851 48195 2909 48196
rect 21424 48152 21504 48172
rect 9187 48112 9196 48152
rect 9236 48112 9676 48152
rect 9716 48112 9725 48152
rect 13027 48112 13036 48152
rect 13076 48112 13324 48152
rect 13364 48112 14092 48152
rect 14132 48112 16396 48152
rect 16436 48112 16445 48152
rect 21292 48112 21504 48152
rect 19459 48068 19517 48069
rect 2467 48028 2476 48068
rect 2516 48028 3340 48068
rect 3380 48028 5548 48068
rect 5588 48028 5597 48068
rect 6787 48028 6796 48068
rect 6836 48028 7084 48068
rect 7124 48028 7564 48068
rect 7604 48028 7613 48068
rect 8131 48028 8140 48068
rect 8180 48028 9868 48068
rect 9908 48028 11360 48068
rect 12355 48028 12364 48068
rect 12404 48028 17012 48068
rect 11320 47984 11360 48028
rect 16972 47984 17012 48028
rect 19459 48028 19468 48068
rect 19508 48028 19564 48068
rect 19604 48028 19613 48068
rect 19459 48027 19517 48028
rect 21292 47984 21332 48112
rect 21424 48092 21504 48112
rect 1699 47944 1708 47984
rect 1748 47944 4684 47984
rect 4724 47944 6892 47984
rect 6932 47944 6941 47984
rect 7267 47944 7276 47984
rect 7316 47944 7660 47984
rect 7700 47944 7709 47984
rect 7756 47944 10252 47984
rect 10292 47944 10301 47984
rect 11320 47944 12460 47984
rect 12500 47944 12509 47984
rect 13603 47944 13612 47984
rect 13652 47944 13900 47984
rect 13940 47944 13949 47984
rect 14947 47944 14956 47984
rect 14996 47944 16012 47984
rect 16052 47944 16204 47984
rect 16244 47944 16253 47984
rect 16963 47944 16972 47984
rect 17012 47944 17021 47984
rect 17731 47944 17740 47984
rect 17780 47944 18220 47984
rect 18260 47944 18269 47984
rect 19267 47944 19276 47984
rect 19316 47944 19948 47984
rect 19988 47944 21332 47984
rect 6892 47900 6932 47944
rect 7756 47900 7796 47944
rect 2371 47860 2380 47900
rect 2420 47860 4204 47900
rect 4244 47860 5588 47900
rect 6595 47860 6604 47900
rect 6644 47860 6653 47900
rect 6892 47860 7796 47900
rect 8227 47900 8285 47901
rect 8515 47900 8573 47901
rect 14275 47900 14333 47901
rect 8227 47860 8236 47900
rect 8276 47860 8524 47900
rect 8564 47860 8573 47900
rect 5548 47816 5588 47860
rect 6604 47816 6644 47860
rect 8227 47859 8285 47860
rect 8515 47859 8573 47860
rect 9868 47860 11404 47900
rect 11444 47860 11453 47900
rect 14190 47860 14284 47900
rect 14324 47860 14333 47900
rect 18220 47900 18260 47944
rect 18220 47860 19852 47900
rect 19892 47860 19901 47900
rect 9868 47816 9908 47860
rect 14275 47859 14333 47860
rect 21424 47816 21504 47836
rect 2467 47776 2476 47816
rect 2516 47776 2956 47816
rect 2996 47776 3005 47816
rect 5548 47776 6124 47816
rect 6164 47776 6644 47816
rect 9283 47776 9292 47816
rect 9332 47776 9908 47816
rect 10723 47776 10732 47816
rect 10772 47776 10924 47816
rect 10964 47776 21504 47816
rect 21424 47756 21504 47776
rect 2563 47692 2572 47732
rect 2612 47692 3244 47732
rect 3284 47692 3293 47732
rect 3340 47692 18124 47732
rect 18164 47692 18173 47732
rect 0 47648 80 47668
rect 1987 47648 2045 47649
rect 0 47608 1996 47648
rect 2036 47608 2045 47648
rect 0 47588 80 47608
rect 1987 47607 2045 47608
rect 3139 47648 3197 47649
rect 3340 47648 3380 47692
rect 3139 47608 3148 47648
rect 3188 47608 3380 47648
rect 4919 47608 4928 47648
rect 4968 47608 5010 47648
rect 5050 47608 5092 47648
rect 5132 47608 5174 47648
rect 5214 47608 5256 47648
rect 5296 47608 5305 47648
rect 5644 47608 6412 47648
rect 6452 47608 6461 47648
rect 20039 47608 20048 47648
rect 20088 47608 20130 47648
rect 20170 47608 20212 47648
rect 20252 47608 20294 47648
rect 20334 47608 20376 47648
rect 20416 47608 20425 47648
rect 3139 47607 3197 47608
rect 5644 47564 5684 47608
rect 9571 47564 9629 47565
rect 18307 47564 18365 47565
rect 5635 47524 5644 47564
rect 5684 47524 5693 47564
rect 9571 47524 9580 47564
rect 9620 47524 18316 47564
rect 18356 47524 18365 47564
rect 9571 47523 9629 47524
rect 18307 47523 18365 47524
rect 9187 47480 9245 47481
rect 10819 47480 10877 47481
rect 21424 47480 21504 47500
rect 9187 47440 9196 47480
rect 9236 47440 9292 47480
rect 9332 47440 9341 47480
rect 10819 47440 10828 47480
rect 10868 47440 10908 47480
rect 16291 47440 16300 47480
rect 16340 47440 21504 47480
rect 9187 47439 9245 47440
rect 10819 47439 10877 47440
rect 10828 47396 10868 47439
rect 21424 47420 21504 47440
rect 15715 47396 15773 47397
rect 5731 47356 5740 47396
rect 5780 47356 10868 47396
rect 10915 47356 10924 47396
rect 10964 47356 15724 47396
rect 15764 47356 15773 47396
rect 16579 47356 16588 47396
rect 16628 47356 16876 47396
rect 16916 47356 16925 47396
rect 4579 47312 4637 47313
rect 8515 47312 8573 47313
rect 10828 47312 10868 47356
rect 15715 47355 15773 47356
rect 4494 47272 4588 47312
rect 4628 47272 6124 47312
rect 6164 47272 6173 47312
rect 6691 47272 6700 47312
rect 6740 47272 6988 47312
rect 7028 47272 7037 47312
rect 8515 47272 8524 47312
rect 8564 47272 8716 47312
rect 8756 47272 8765 47312
rect 10819 47272 10828 47312
rect 10868 47272 10877 47312
rect 12163 47272 12172 47312
rect 12212 47272 13804 47312
rect 13844 47272 18028 47312
rect 18068 47272 18077 47312
rect 4579 47271 4637 47272
rect 8515 47271 8573 47272
rect 5539 47188 5548 47228
rect 5588 47188 10924 47228
rect 10964 47188 10973 47228
rect 10627 47144 10685 47145
rect 21424 47144 21504 47164
rect 9091 47104 9100 47144
rect 9140 47104 10348 47144
rect 10388 47104 10636 47144
rect 10676 47104 10685 47144
rect 19267 47104 19276 47144
rect 19316 47104 21504 47144
rect 10627 47103 10685 47104
rect 21424 47084 21504 47104
rect 2179 47020 2188 47060
rect 2228 47020 14956 47060
rect 14996 47020 16684 47060
rect 16724 47020 16733 47060
rect 17635 47020 17644 47060
rect 17684 47020 18604 47060
rect 18644 47020 18653 47060
rect 0 46976 80 46996
rect 13411 46976 13469 46977
rect 0 46936 1612 46976
rect 1652 46936 1661 46976
rect 2851 46936 2860 46976
rect 2900 46936 13420 46976
rect 13460 46936 13469 46976
rect 0 46916 80 46936
rect 13411 46935 13469 46936
rect 18124 46936 19852 46976
rect 19892 46936 19901 46976
rect 18124 46893 18164 46936
rect 6595 46892 6653 46893
rect 18115 46892 18173 46893
rect 3679 46852 3688 46892
rect 3728 46852 3770 46892
rect 3810 46852 3852 46892
rect 3892 46852 3934 46892
rect 3974 46852 4016 46892
rect 4056 46852 4065 46892
rect 6307 46852 6316 46892
rect 6356 46852 6604 46892
rect 6644 46852 6653 46892
rect 8803 46852 8812 46892
rect 8852 46852 9292 46892
rect 9332 46852 10252 46892
rect 10292 46852 10301 46892
rect 10819 46852 10828 46892
rect 10868 46852 12556 46892
rect 12596 46852 12605 46892
rect 14083 46852 14092 46892
rect 14132 46852 16204 46892
rect 16244 46852 18124 46892
rect 18164 46852 18173 46892
rect 18799 46852 18808 46892
rect 18848 46852 18890 46892
rect 18930 46852 18972 46892
rect 19012 46852 19054 46892
rect 19094 46852 19136 46892
rect 19176 46852 19185 46892
rect 6595 46851 6653 46852
rect 18115 46851 18173 46852
rect 9571 46808 9629 46809
rect 21424 46808 21504 46828
rect 1411 46768 1420 46808
rect 1460 46768 1900 46808
rect 1940 46768 2540 46808
rect 2500 46724 2540 46768
rect 6604 46768 9580 46808
rect 9620 46768 9629 46808
rect 14371 46768 14380 46808
rect 14420 46768 21504 46808
rect 6604 46724 6644 46768
rect 9571 46767 9629 46768
rect 21424 46748 21504 46768
rect 18019 46724 18077 46725
rect 2500 46684 6644 46724
rect 6691 46684 6700 46724
rect 6740 46684 7564 46724
rect 7604 46684 7613 46724
rect 8611 46684 8620 46724
rect 8660 46684 14764 46724
rect 14804 46684 14813 46724
rect 18019 46684 18028 46724
rect 18068 46684 19796 46724
rect 18019 46683 18077 46684
rect 7075 46640 7133 46641
rect 8131 46640 8189 46641
rect 9187 46640 9245 46641
rect 19756 46640 19796 46684
rect 163 46600 172 46640
rect 212 46600 1324 46640
rect 1364 46600 1373 46640
rect 1699 46600 1708 46640
rect 1748 46600 2188 46640
rect 2228 46600 2237 46640
rect 5443 46600 5452 46640
rect 5492 46600 5501 46640
rect 6990 46600 7084 46640
rect 7124 46600 7133 46640
rect 8046 46600 8140 46640
rect 8180 46600 8189 46640
rect 9102 46600 9196 46640
rect 9236 46600 9245 46640
rect 11971 46600 11980 46640
rect 12020 46600 12029 46640
rect 19756 46600 20276 46640
rect 20899 46600 20908 46640
rect 20948 46600 20957 46640
rect 5452 46556 5492 46600
rect 7075 46599 7133 46600
rect 8131 46599 8189 46600
rect 9187 46599 9245 46600
rect 5827 46556 5885 46557
rect 11980 46556 12020 46600
rect 20236 46556 20276 46600
rect 20908 46556 20948 46600
rect 2500 46516 2860 46556
rect 2900 46516 2909 46556
rect 5452 46516 5836 46556
rect 5876 46516 5885 46556
rect 6211 46516 6220 46556
rect 6260 46516 6604 46556
rect 6644 46516 6653 46556
rect 7267 46516 7276 46556
rect 7316 46516 8236 46556
rect 8276 46516 8285 46556
rect 11587 46516 11596 46556
rect 11636 46516 12020 46556
rect 15139 46516 15148 46556
rect 15188 46516 20180 46556
rect 20236 46516 20948 46556
rect 0 46304 80 46324
rect 2500 46304 2540 46516
rect 5827 46515 5885 46516
rect 4675 46472 4733 46473
rect 18691 46472 18749 46473
rect 4675 46432 4684 46472
rect 4724 46432 4972 46472
rect 5012 46432 5021 46472
rect 6403 46432 6412 46472
rect 6452 46432 7180 46472
rect 7220 46432 7229 46472
rect 7843 46432 7852 46472
rect 7892 46432 11212 46472
rect 11252 46432 12076 46472
rect 12116 46432 12125 46472
rect 15331 46432 15340 46472
rect 15380 46432 16780 46472
rect 16820 46432 16829 46472
rect 17059 46432 17068 46472
rect 17108 46432 17452 46472
rect 17492 46432 17501 46472
rect 18595 46432 18604 46472
rect 18644 46432 18700 46472
rect 18740 46432 18749 46472
rect 4675 46431 4733 46432
rect 18691 46431 18749 46432
rect 19939 46472 19997 46473
rect 20140 46472 20180 46516
rect 21424 46472 21504 46492
rect 19939 46432 19948 46472
rect 19988 46432 20044 46472
rect 20084 46432 20093 46472
rect 20140 46432 21504 46472
rect 19939 46431 19997 46432
rect 21424 46412 21504 46432
rect 4579 46388 4637 46389
rect 20707 46388 20765 46389
rect 4579 46348 4588 46388
rect 4628 46348 5068 46388
rect 5108 46348 5117 46388
rect 6595 46348 6604 46388
rect 6644 46348 7756 46388
rect 7796 46348 7805 46388
rect 10243 46348 10252 46388
rect 10292 46348 10924 46388
rect 10964 46348 10973 46388
rect 12643 46348 12652 46388
rect 12692 46348 12940 46388
rect 12980 46348 13420 46388
rect 13460 46348 13469 46388
rect 14563 46348 14572 46388
rect 14612 46348 15052 46388
rect 15092 46348 15101 46388
rect 15235 46348 15244 46388
rect 15284 46348 15916 46388
rect 15956 46348 16588 46388
rect 16628 46348 17740 46388
rect 17780 46348 17789 46388
rect 20227 46348 20236 46388
rect 20276 46348 20716 46388
rect 20756 46348 20765 46388
rect 4579 46347 4637 46348
rect 4483 46304 4541 46305
rect 0 46264 2540 46304
rect 3523 46264 3532 46304
rect 3572 46264 4012 46304
rect 4052 46264 4061 46304
rect 4483 46264 4492 46304
rect 4532 46264 4684 46304
rect 4724 46264 4733 46304
rect 5836 46264 6796 46304
rect 6836 46264 6845 46304
rect 0 46244 80 46264
rect 4483 46263 4541 46264
rect 5836 46220 5876 46264
rect 6604 46220 6644 46264
rect 5827 46180 5836 46220
rect 5876 46180 5885 46220
rect 6595 46180 6604 46220
rect 6644 46180 6653 46220
rect 6988 46136 7028 46348
rect 20707 46347 20765 46348
rect 18115 46304 18173 46305
rect 21379 46304 21437 46305
rect 8419 46264 8428 46304
rect 8468 46264 15340 46304
rect 15380 46264 15389 46304
rect 16771 46264 16780 46304
rect 16820 46264 17068 46304
rect 17108 46264 17117 46304
rect 17251 46264 17260 46304
rect 17300 46264 17932 46304
rect 17972 46264 17981 46304
rect 18115 46264 18124 46304
rect 18164 46264 18604 46304
rect 18644 46264 18653 46304
rect 20140 46264 21388 46304
rect 21428 46264 21437 46304
rect 18115 46263 18173 46264
rect 20140 46220 20180 46264
rect 21379 46263 21437 46264
rect 9475 46180 9484 46220
rect 9524 46180 10060 46220
rect 10100 46180 10109 46220
rect 11320 46180 20180 46220
rect 11320 46136 11360 46180
rect 21424 46136 21504 46156
rect 4919 46096 4928 46136
rect 4968 46096 5010 46136
rect 5050 46096 5092 46136
rect 5132 46096 5174 46136
rect 5214 46096 5256 46136
rect 5296 46096 5305 46136
rect 6979 46096 6988 46136
rect 7028 46096 7037 46136
rect 7852 46096 11360 46136
rect 13219 46096 13228 46136
rect 13268 46096 17740 46136
rect 17780 46096 17789 46136
rect 18115 46096 18124 46136
rect 18164 46096 18412 46136
rect 18452 46096 18461 46136
rect 20039 46096 20048 46136
rect 20088 46096 20130 46136
rect 20170 46096 20212 46136
rect 20252 46096 20294 46136
rect 20334 46096 20376 46136
rect 20416 46096 20425 46136
rect 21292 46096 21504 46136
rect 7852 46052 7892 46096
rect 2659 46012 2668 46052
rect 2708 46012 3340 46052
rect 3380 46012 5204 46052
rect 5347 46012 5356 46052
rect 5396 46012 6316 46052
rect 6356 46012 7892 46052
rect 9571 46012 9580 46052
rect 9620 46012 9868 46052
rect 9908 46012 9917 46052
rect 12835 46012 12844 46052
rect 12884 46012 12893 46052
rect 13315 46012 13324 46052
rect 13364 46012 14764 46052
rect 14804 46012 16588 46052
rect 16628 46012 16637 46052
rect 4579 45968 4637 45969
rect 5164 45968 5204 46012
rect 12844 45968 12884 46012
rect 21292 45968 21332 46096
rect 21424 46076 21504 46096
rect 2851 45928 2860 45968
rect 2900 45928 4588 45968
rect 4628 45928 5068 45968
rect 5108 45928 5117 45968
rect 5164 45928 11360 45968
rect 12643 45928 12652 45968
rect 12692 45928 12884 45968
rect 13891 45928 13900 45968
rect 13940 45928 16108 45968
rect 16148 45928 16157 45968
rect 20140 45928 21332 45968
rect 4579 45927 4637 45928
rect 5827 45884 5885 45885
rect 6595 45884 6653 45885
rect 3331 45844 3340 45884
rect 3380 45844 4684 45884
rect 4724 45844 4733 45884
rect 5827 45844 5836 45884
rect 5876 45844 6220 45884
rect 6260 45844 6269 45884
rect 6403 45844 6412 45884
rect 6452 45844 6604 45884
rect 6644 45844 6653 45884
rect 5827 45843 5885 45844
rect 6595 45843 6653 45844
rect 7843 45884 7901 45885
rect 11320 45884 11360 45928
rect 20140 45884 20180 45928
rect 7843 45844 7852 45884
rect 7892 45844 7988 45884
rect 9667 45844 9676 45884
rect 9716 45844 9725 45884
rect 11320 45844 15244 45884
rect 15284 45844 15293 45884
rect 15436 45844 20180 45884
rect 7843 45843 7901 45844
rect 7948 45800 7988 45844
rect 9571 45800 9629 45801
rect 2092 45760 6932 45800
rect 7555 45760 7564 45800
rect 7604 45760 7756 45800
rect 7796 45760 7805 45800
rect 7939 45760 7948 45800
rect 7988 45760 8524 45800
rect 8564 45760 8573 45800
rect 9486 45760 9580 45800
rect 9620 45760 9629 45800
rect 9676 45800 9716 45844
rect 9676 45760 10828 45800
rect 10868 45760 12460 45800
rect 12500 45760 14092 45800
rect 14132 45760 14141 45800
rect 0 45632 80 45652
rect 2092 45632 2132 45760
rect 4579 45716 4637 45717
rect 4494 45676 4588 45716
rect 4628 45676 4637 45716
rect 4579 45675 4637 45676
rect 5923 45716 5981 45717
rect 6892 45716 6932 45760
rect 9571 45759 9629 45760
rect 5923 45676 5932 45716
rect 5972 45676 6028 45716
rect 6068 45676 6077 45716
rect 6892 45676 11596 45716
rect 11636 45676 11645 45716
rect 5923 45675 5981 45676
rect 0 45592 1228 45632
rect 1268 45592 2132 45632
rect 3043 45592 3052 45632
rect 3092 45592 4972 45632
rect 5012 45592 5021 45632
rect 5827 45592 5836 45632
rect 5876 45592 6316 45632
rect 6356 45592 6365 45632
rect 6691 45592 6700 45632
rect 6740 45592 8236 45632
rect 8276 45592 8285 45632
rect 11011 45592 11020 45632
rect 11060 45592 11692 45632
rect 11732 45592 11741 45632
rect 0 45572 80 45592
rect 4483 45508 4492 45548
rect 4532 45508 6412 45548
rect 6452 45508 6461 45548
rect 6979 45508 6988 45548
rect 7028 45508 7180 45548
rect 7220 45508 7372 45548
rect 7412 45508 7421 45548
rect 8707 45508 8716 45548
rect 8756 45508 9388 45548
rect 9428 45508 9437 45548
rect 7075 45464 7133 45465
rect 2947 45424 2956 45464
rect 2996 45424 4204 45464
rect 4244 45424 4253 45464
rect 6883 45424 6892 45464
rect 6932 45424 7084 45464
rect 7124 45424 7133 45464
rect 7075 45423 7133 45424
rect 8800 45424 10924 45464
rect 10964 45424 10973 45464
rect 13411 45424 13420 45464
rect 13460 45424 15244 45464
rect 15284 45424 15293 45464
rect 8800 45380 8840 45424
rect 15436 45380 15476 45844
rect 16099 45800 16157 45801
rect 21424 45800 21504 45820
rect 15619 45760 15628 45800
rect 15668 45760 15820 45800
rect 15860 45760 15869 45800
rect 16003 45760 16012 45800
rect 16052 45760 16108 45800
rect 16148 45760 16157 45800
rect 17059 45760 17068 45800
rect 17108 45760 18220 45800
rect 18260 45760 18269 45800
rect 20140 45760 21504 45800
rect 16099 45759 16157 45760
rect 17443 45716 17501 45717
rect 20140 45716 20180 45760
rect 21424 45740 21504 45760
rect 17443 45676 17452 45716
rect 17492 45676 20180 45716
rect 17443 45675 17501 45676
rect 16771 45592 16780 45632
rect 16820 45592 17932 45632
rect 17972 45592 17981 45632
rect 15523 45508 15532 45548
rect 15572 45508 16108 45548
rect 16148 45508 17452 45548
rect 17492 45508 17501 45548
rect 17731 45508 17740 45548
rect 17780 45508 18028 45548
rect 18068 45508 18077 45548
rect 18700 45508 19660 45548
rect 19700 45508 19709 45548
rect 15811 45424 15820 45464
rect 15860 45424 18412 45464
rect 18452 45424 18461 45464
rect 3679 45340 3688 45380
rect 3728 45340 3770 45380
rect 3810 45340 3852 45380
rect 3892 45340 3934 45380
rect 3974 45340 4016 45380
rect 4056 45340 4065 45380
rect 4963 45340 4972 45380
rect 5012 45340 5932 45380
rect 5972 45340 8840 45380
rect 9859 45340 9868 45380
rect 9908 45340 15476 45380
rect 13699 45296 13757 45297
rect 15043 45296 15101 45297
rect 15820 45296 15860 45424
rect 18700 45380 18740 45508
rect 19843 45464 19901 45465
rect 21424 45464 21504 45484
rect 19843 45424 19852 45464
rect 19892 45424 21504 45464
rect 19843 45423 19901 45424
rect 21424 45404 21504 45424
rect 17923 45340 17932 45380
rect 17972 45340 18740 45380
rect 18799 45340 18808 45380
rect 18848 45340 18890 45380
rect 18930 45340 18972 45380
rect 19012 45340 19054 45380
rect 19094 45340 19136 45380
rect 19176 45340 19185 45380
rect 4387 45256 4396 45296
rect 4436 45256 4445 45296
rect 4492 45256 11212 45296
rect 11252 45256 11261 45296
rect 11308 45256 13708 45296
rect 13748 45256 13757 45296
rect 14958 45256 15052 45296
rect 15092 45256 15101 45296
rect 15235 45256 15244 45296
rect 15284 45256 15860 45296
rect 4396 45212 4436 45256
rect 3907 45172 3916 45212
rect 3956 45172 4436 45212
rect 2755 45128 2813 45129
rect 4492 45128 4532 45256
rect 7651 45212 7709 45213
rect 11308 45212 11348 45256
rect 13699 45255 13757 45256
rect 15043 45255 15101 45256
rect 7267 45172 7276 45212
rect 7316 45172 7660 45212
rect 7700 45172 7709 45212
rect 9955 45172 9964 45212
rect 10004 45172 11348 45212
rect 11395 45212 11453 45213
rect 19843 45212 19901 45213
rect 11395 45172 11404 45212
rect 11444 45172 11538 45212
rect 12940 45172 16300 45212
rect 16340 45172 16349 45212
rect 18979 45172 18988 45212
rect 19028 45172 19852 45212
rect 19892 45172 19901 45212
rect 7651 45171 7709 45172
rect 11395 45171 11453 45172
rect 2500 45088 2764 45128
rect 2804 45088 4532 45128
rect 4675 45128 4733 45129
rect 12940 45128 12980 45172
rect 19843 45171 19901 45172
rect 21424 45128 21504 45148
rect 4675 45088 4684 45128
rect 4724 45088 4972 45128
rect 5012 45088 5021 45128
rect 7459 45088 7468 45128
rect 7508 45088 8140 45128
rect 8180 45088 8189 45128
rect 8323 45088 8332 45128
rect 8372 45088 8620 45128
rect 8660 45088 8669 45128
rect 9187 45088 9196 45128
rect 9236 45088 9868 45128
rect 9908 45088 12980 45128
rect 13036 45088 21504 45128
rect 0 44960 80 44980
rect 2500 44960 2540 45088
rect 2755 45087 2813 45088
rect 4675 45087 4733 45088
rect 4771 45044 4829 45045
rect 13036 45044 13076 45088
rect 21424 45068 21504 45088
rect 4771 45004 4780 45044
rect 4820 45004 9772 45044
rect 9812 45004 9821 45044
rect 10723 45004 10732 45044
rect 10772 45004 13076 45044
rect 13795 45004 13804 45044
rect 13844 45004 16972 45044
rect 17012 45004 17021 45044
rect 18883 45004 18892 45044
rect 18932 45004 19756 45044
rect 19796 45004 19805 45044
rect 4771 45003 4829 45004
rect 7267 44960 7325 44961
rect 0 44920 2540 44960
rect 4003 44920 4012 44960
rect 4052 44920 4780 44960
rect 4820 44920 4829 44960
rect 6499 44920 6508 44960
rect 6548 44920 6796 44960
rect 6836 44920 7276 44960
rect 7316 44920 7325 44960
rect 7747 44920 7756 44960
rect 7796 44920 8236 44960
rect 8276 44920 8285 44960
rect 9283 44920 9292 44960
rect 9332 44920 9676 44960
rect 9716 44920 9725 44960
rect 14956 44920 15572 44960
rect 0 44900 80 44920
rect 7267 44919 7325 44920
rect 4483 44876 4541 44877
rect 8899 44876 8957 44877
rect 4291 44836 4300 44876
rect 4340 44836 4492 44876
rect 4532 44836 4541 44876
rect 8611 44836 8620 44876
rect 8660 44836 8908 44876
rect 8948 44836 8957 44876
rect 4483 44835 4541 44836
rect 8899 44835 8957 44836
rect 9004 44836 13708 44876
rect 13748 44836 13757 44876
rect 7843 44792 7901 44793
rect 8131 44792 8189 44793
rect 2179 44752 2188 44792
rect 2228 44752 4204 44792
rect 4244 44752 4253 44792
rect 7758 44752 7852 44792
rect 7892 44752 7901 44792
rect 8035 44752 8044 44792
rect 8084 44752 8140 44792
rect 8180 44752 8189 44792
rect 7843 44751 7901 44752
rect 8131 44751 8189 44752
rect 9004 44708 9044 44836
rect 14956 44792 14996 44920
rect 10243 44752 10252 44792
rect 10292 44752 14996 44792
rect 15532 44792 15572 44920
rect 21424 44792 21504 44812
rect 15532 44752 21504 44792
rect 21424 44732 21504 44752
rect 19267 44708 19325 44709
rect 7459 44668 7468 44708
rect 7508 44668 9044 44708
rect 13891 44668 13900 44708
rect 13940 44668 19276 44708
rect 19316 44668 19468 44708
rect 19508 44668 19517 44708
rect 19267 44667 19325 44668
rect 9475 44624 9533 44625
rect 3235 44584 3244 44624
rect 3284 44584 4396 44624
rect 4436 44584 4445 44624
rect 4919 44584 4928 44624
rect 4968 44584 5010 44624
rect 5050 44584 5092 44624
rect 5132 44584 5174 44624
rect 5214 44584 5256 44624
rect 5296 44584 5305 44624
rect 7756 44584 9484 44624
rect 9524 44584 12940 44624
rect 12980 44584 12989 44624
rect 13315 44584 13324 44624
rect 13364 44584 13373 44624
rect 13795 44584 13804 44624
rect 13844 44584 13996 44624
rect 14036 44584 14668 44624
rect 14708 44584 14860 44624
rect 14900 44584 14909 44624
rect 20039 44584 20048 44624
rect 20088 44584 20130 44624
rect 20170 44584 20212 44624
rect 20252 44584 20294 44624
rect 20334 44584 20376 44624
rect 20416 44584 20425 44624
rect 7756 44540 7796 44584
rect 9475 44583 9533 44584
rect 13324 44540 13364 44584
rect 4300 44500 7796 44540
rect 8323 44500 8332 44540
rect 8372 44500 10348 44540
rect 10388 44500 10397 44540
rect 13324 44500 13708 44540
rect 13748 44500 14092 44540
rect 14132 44500 14141 44540
rect 355 44416 364 44456
rect 404 44416 3340 44456
rect 3380 44416 3389 44456
rect 4300 44372 4340 44500
rect 4579 44456 4637 44457
rect 18691 44456 18749 44457
rect 21424 44456 21504 44476
rect 4494 44416 4588 44456
rect 4628 44416 4637 44456
rect 4579 44415 4637 44416
rect 8140 44416 9100 44456
rect 9140 44416 9149 44456
rect 14275 44416 14284 44456
rect 14324 44416 15244 44456
rect 15284 44416 15293 44456
rect 16195 44416 16204 44456
rect 16244 44416 17164 44456
rect 17204 44416 17213 44456
rect 18606 44416 18700 44456
rect 18740 44416 21504 44456
rect 2500 44332 4340 44372
rect 4387 44372 4445 44373
rect 4387 44332 4396 44372
rect 4436 44332 6892 44372
rect 6932 44332 6941 44372
rect 0 44288 80 44308
rect 2500 44288 2540 44332
rect 4387 44331 4445 44332
rect 5347 44288 5405 44289
rect 8140 44288 8180 44416
rect 18691 44415 18749 44416
rect 21424 44396 21504 44416
rect 11320 44332 14668 44372
rect 14708 44332 17644 44372
rect 17684 44332 17693 44372
rect 0 44248 2540 44288
rect 4099 44248 4108 44288
rect 4148 44248 4876 44288
rect 4916 44248 5356 44288
rect 5396 44248 5405 44288
rect 6115 44248 6124 44288
rect 6164 44248 6508 44288
rect 6548 44248 6557 44288
rect 7075 44248 7084 44288
rect 7124 44248 8140 44288
rect 8180 44248 8189 44288
rect 9091 44248 9100 44288
rect 9140 44248 10252 44288
rect 10292 44248 10301 44288
rect 0 44228 80 44248
rect 5347 44247 5405 44248
rect 11320 44204 11360 44332
rect 11779 44248 11788 44288
rect 11828 44248 14380 44288
rect 14420 44248 14429 44288
rect 15139 44248 15148 44288
rect 15188 44248 15436 44288
rect 15476 44248 15485 44288
rect 16771 44248 16780 44288
rect 16820 44248 17260 44288
rect 17300 44248 17309 44288
rect 15043 44204 15101 44205
rect 6883 44164 6892 44204
rect 6932 44164 11360 44204
rect 13411 44164 13420 44204
rect 13460 44164 14284 44204
rect 14324 44164 14333 44204
rect 14958 44164 15052 44204
rect 15092 44164 15101 44204
rect 17635 44164 17644 44204
rect 17684 44164 19948 44204
rect 19988 44164 19997 44204
rect 15043 44163 15101 44164
rect 2275 44120 2333 44121
rect 8323 44120 8381 44121
rect 21424 44120 21504 44140
rect 2275 44080 2284 44120
rect 2324 44080 2572 44120
rect 2612 44080 2621 44120
rect 2755 44080 2764 44120
rect 2804 44080 3148 44120
rect 3188 44080 6796 44120
rect 6836 44080 7468 44120
rect 7508 44080 7517 44120
rect 8238 44080 8332 44120
rect 8372 44080 8381 44120
rect 17827 44080 17836 44120
rect 17876 44080 18316 44120
rect 18356 44080 21504 44120
rect 2275 44079 2333 44080
rect 8323 44079 8381 44080
rect 21424 44060 21504 44080
rect 1987 43996 1996 44036
rect 2036 43996 8236 44036
rect 8276 43996 8716 44036
rect 8756 43996 8765 44036
rect 12547 43996 12556 44036
rect 12596 43996 13228 44036
rect 13268 43996 13277 44036
rect 12835 43912 12844 43952
rect 12884 43912 13996 43952
rect 14036 43912 14045 43952
rect 14179 43912 14188 43952
rect 14228 43912 14956 43952
rect 14996 43912 15005 43952
rect 18307 43912 18316 43952
rect 18356 43912 18508 43952
rect 18548 43912 18557 43952
rect 3679 43828 3688 43868
rect 3728 43828 3770 43868
rect 3810 43828 3852 43868
rect 3892 43828 3934 43868
rect 3974 43828 4016 43868
rect 4056 43828 4065 43868
rect 8515 43828 8524 43868
rect 8564 43828 14668 43868
rect 14708 43828 17164 43868
rect 17204 43828 17213 43868
rect 18799 43828 18808 43868
rect 18848 43828 18890 43868
rect 18930 43828 18972 43868
rect 19012 43828 19054 43868
rect 19094 43828 19136 43868
rect 19176 43828 19185 43868
rect 21424 43784 21504 43804
rect 8803 43744 8812 43784
rect 8852 43744 9004 43784
rect 9044 43744 21504 43784
rect 21424 43724 21504 43744
rect 10915 43660 10924 43700
rect 10964 43660 20180 43700
rect 0 43616 80 43636
rect 4291 43616 4349 43617
rect 0 43576 4300 43616
rect 4340 43576 4349 43616
rect 13411 43576 13420 43616
rect 13460 43576 14092 43616
rect 14132 43576 14141 43616
rect 0 43556 80 43576
rect 4291 43575 4349 43576
rect 6499 43492 6508 43532
rect 6548 43492 8140 43532
rect 8180 43492 9964 43532
rect 10004 43492 11596 43532
rect 11636 43492 12556 43532
rect 12596 43492 17932 43532
rect 17972 43492 17981 43532
rect 20140 43448 20180 43660
rect 21424 43448 21504 43468
rect 3043 43408 3052 43448
rect 3092 43408 4876 43448
rect 4916 43408 4925 43448
rect 6211 43408 6220 43448
rect 6260 43408 11308 43448
rect 11348 43408 11357 43448
rect 13315 43408 13324 43448
rect 13364 43408 14476 43448
rect 14516 43408 14525 43448
rect 15331 43408 15340 43448
rect 15380 43408 16588 43448
rect 16628 43408 16637 43448
rect 20140 43408 21504 43448
rect 4876 43364 4916 43408
rect 21424 43388 21504 43408
rect 4876 43324 8044 43364
rect 8084 43324 8093 43364
rect 12835 43324 12844 43364
rect 12884 43324 13228 43364
rect 13268 43324 13277 43364
rect 12739 43240 12748 43280
rect 12788 43240 13612 43280
rect 13652 43240 13661 43280
rect 14371 43240 14380 43280
rect 14420 43240 16876 43280
rect 16916 43240 16925 43280
rect 11683 43156 11692 43196
rect 11732 43156 16780 43196
rect 16820 43156 16829 43196
rect 18307 43156 18316 43196
rect 18356 43156 20852 43196
rect 20812 43112 20852 43156
rect 21424 43112 21504 43132
rect 4919 43072 4928 43112
rect 4968 43072 5010 43112
rect 5050 43072 5092 43112
rect 5132 43072 5174 43112
rect 5214 43072 5256 43112
rect 5296 43072 5305 43112
rect 20039 43072 20048 43112
rect 20088 43072 20130 43112
rect 20170 43072 20212 43112
rect 20252 43072 20294 43112
rect 20334 43072 20376 43112
rect 20416 43072 20425 43112
rect 20812 43072 21504 43112
rect 21424 43052 21504 43072
rect 739 43028 797 43029
rect 739 42988 748 43028
rect 788 42988 7372 43028
rect 7412 42988 7421 43028
rect 739 42987 797 42988
rect 0 42944 80 42964
rect 0 42904 2092 42944
rect 2132 42904 2141 42944
rect 2668 42904 3052 42944
rect 3092 42904 3101 42944
rect 5347 42904 5356 42944
rect 5396 42904 5405 42944
rect 0 42884 80 42904
rect 2668 42776 2708 42904
rect 5356 42860 5396 42904
rect 10339 42860 10397 42861
rect 4195 42820 4204 42860
rect 4244 42820 5260 42860
rect 5300 42820 5309 42860
rect 5356 42820 5740 42860
rect 5780 42820 5789 42860
rect 9571 42820 9580 42860
rect 9620 42820 9772 42860
rect 9812 42820 10348 42860
rect 10388 42820 10397 42860
rect 5356 42776 5396 42820
rect 10339 42819 10397 42820
rect 15715 42860 15773 42861
rect 15715 42820 15724 42860
rect 15764 42820 16684 42860
rect 16724 42820 16733 42860
rect 15715 42819 15773 42820
rect 6595 42776 6653 42777
rect 10723 42776 10781 42777
rect 2659 42736 2668 42776
rect 2708 42736 2717 42776
rect 3235 42736 3244 42776
rect 3284 42736 4300 42776
rect 4340 42736 4349 42776
rect 4483 42736 4492 42776
rect 4532 42736 4541 42776
rect 5059 42736 5068 42776
rect 5108 42736 5396 42776
rect 5827 42736 5836 42776
rect 5876 42736 6604 42776
rect 6644 42736 6653 42776
rect 10638 42736 10732 42776
rect 10772 42736 10781 42776
rect 4492 42692 4532 42736
rect 6595 42735 6653 42736
rect 10723 42735 10781 42736
rect 12643 42776 12701 42777
rect 21424 42776 21504 42796
rect 12643 42736 12652 42776
rect 12692 42736 12748 42776
rect 12788 42736 12797 42776
rect 13219 42736 13228 42776
rect 13268 42736 13996 42776
rect 14036 42736 15916 42776
rect 15956 42736 16300 42776
rect 16340 42736 17548 42776
rect 17588 42736 17597 42776
rect 20227 42736 20236 42776
rect 20276 42736 21504 42776
rect 12643 42735 12701 42736
rect 13228 42692 13268 42736
rect 21424 42716 21504 42736
rect 3715 42652 3724 42692
rect 3764 42652 4396 42692
rect 4436 42652 4445 42692
rect 4492 42652 5356 42692
rect 5396 42652 5405 42692
rect 9091 42652 9100 42692
rect 9140 42652 10060 42692
rect 10100 42652 10109 42692
rect 11971 42652 11980 42692
rect 12020 42652 13268 42692
rect 11971 42608 12029 42609
rect 3619 42568 3628 42608
rect 3668 42568 4492 42608
rect 4532 42568 4541 42608
rect 11971 42568 11980 42608
rect 12020 42568 19756 42608
rect 19796 42568 20044 42608
rect 20084 42568 20093 42608
rect 11971 42567 12029 42568
rect 5155 42484 5164 42524
rect 5204 42484 5740 42524
rect 5780 42484 5789 42524
rect 6595 42484 6604 42524
rect 6644 42484 19564 42524
rect 19604 42484 19613 42524
rect 21424 42440 21504 42460
rect 2467 42400 2476 42440
rect 2516 42400 4340 42440
rect 5347 42400 5356 42440
rect 5396 42400 11980 42440
rect 12020 42400 12029 42440
rect 18115 42400 18124 42440
rect 18164 42400 21504 42440
rect 4300 42356 4340 42400
rect 21424 42380 21504 42400
rect 3679 42316 3688 42356
rect 3728 42316 3770 42356
rect 3810 42316 3852 42356
rect 3892 42316 3934 42356
rect 3974 42316 4016 42356
rect 4056 42316 4065 42356
rect 4300 42316 6700 42356
rect 6740 42316 6749 42356
rect 18799 42316 18808 42356
rect 18848 42316 18890 42356
rect 18930 42316 18972 42356
rect 19012 42316 19054 42356
rect 19094 42316 19136 42356
rect 19176 42316 19185 42356
rect 0 42272 80 42292
rect 11587 42272 11645 42273
rect 0 42232 5548 42272
rect 5588 42232 5597 42272
rect 10243 42232 10252 42272
rect 10292 42232 11596 42272
rect 11636 42232 20524 42272
rect 20564 42232 20573 42272
rect 0 42212 80 42232
rect 11587 42231 11645 42232
rect 3907 42148 3916 42188
rect 3956 42148 4684 42188
rect 4724 42148 4733 42188
rect 10723 42104 10781 42105
rect 21424 42104 21504 42124
rect 3043 42064 3052 42104
rect 3092 42064 3724 42104
rect 3764 42064 5356 42104
rect 5396 42064 5405 42104
rect 10723 42064 10732 42104
rect 10772 42064 14668 42104
rect 14708 42064 17932 42104
rect 17972 42064 17981 42104
rect 19843 42064 19852 42104
rect 19892 42064 21504 42104
rect 10723 42063 10781 42064
rect 21424 42044 21504 42064
rect 4387 41980 4396 42020
rect 4436 41980 4780 42020
rect 4820 41980 4829 42020
rect 12835 41980 12844 42020
rect 12884 41980 13036 42020
rect 13076 41980 14956 42020
rect 14996 41980 15724 42020
rect 15764 41980 15773 42020
rect 18115 41980 18124 42020
rect 18164 41980 19660 42020
rect 19700 41980 19709 42020
rect 10147 41936 10205 41937
rect 11011 41936 11069 41937
rect 1795 41896 1804 41936
rect 1844 41896 2476 41936
rect 2516 41896 2525 41936
rect 3235 41896 3244 41936
rect 3284 41896 4204 41936
rect 4244 41896 4253 41936
rect 9763 41896 9772 41936
rect 9812 41896 9964 41936
rect 10004 41896 10013 41936
rect 10062 41896 10156 41936
rect 10196 41896 10205 41936
rect 10723 41896 10732 41936
rect 10772 41896 11020 41936
rect 11060 41896 11069 41936
rect 12739 41896 12748 41936
rect 12788 41896 14860 41936
rect 14900 41896 14909 41936
rect 16291 41896 16300 41936
rect 16340 41896 16492 41936
rect 16532 41896 16541 41936
rect 17251 41896 17260 41936
rect 17300 41896 17740 41936
rect 17780 41896 18700 41936
rect 18740 41896 18988 41936
rect 19028 41896 19037 41936
rect 10147 41895 10205 41896
rect 11011 41895 11069 41896
rect 2500 41812 8140 41852
rect 8180 41812 8189 41852
rect 8803 41812 8812 41852
rect 8852 41812 9676 41852
rect 9716 41812 9725 41852
rect 10051 41812 10060 41852
rect 10100 41812 16396 41852
rect 16436 41812 16445 41852
rect 2500 41768 2540 41812
rect 21424 41768 21504 41788
rect 739 41728 748 41768
rect 788 41728 2540 41768
rect 4492 41728 5068 41768
rect 5108 41728 5117 41768
rect 5251 41728 5260 41768
rect 5300 41728 5309 41768
rect 12355 41728 12364 41768
rect 12404 41728 14476 41768
rect 14516 41728 14525 41768
rect 15619 41728 15628 41768
rect 15668 41728 16108 41768
rect 16148 41728 16157 41768
rect 19459 41728 19468 41768
rect 19508 41728 21504 41768
rect 4492 41684 4532 41728
rect 5260 41684 5300 41728
rect 21424 41708 21504 41728
rect 460 41644 4532 41684
rect 4780 41644 11500 41684
rect 11540 41644 11549 41684
rect 13219 41644 13228 41684
rect 13268 41644 13900 41684
rect 13940 41644 13949 41684
rect 0 41600 80 41620
rect 460 41600 500 41644
rect 3523 41600 3581 41601
rect 4780 41600 4820 41644
rect 6892 41600 6932 41644
rect 11971 41600 12029 41601
rect 0 41560 500 41600
rect 2668 41560 3532 41600
rect 3572 41560 3581 41600
rect 3811 41560 3820 41600
rect 3860 41560 4108 41600
rect 4148 41560 4300 41600
rect 4340 41560 4349 41600
rect 4771 41560 4780 41600
rect 4820 41560 4829 41600
rect 4919 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 5305 41600
rect 5635 41560 5644 41600
rect 5684 41560 5932 41600
rect 5972 41560 5981 41600
rect 6307 41560 6316 41600
rect 6356 41560 6700 41600
rect 6740 41560 6749 41600
rect 6883 41560 6892 41600
rect 6932 41560 6972 41600
rect 8035 41560 8044 41600
rect 8084 41560 8620 41600
rect 8660 41560 8669 41600
rect 11779 41560 11788 41600
rect 11828 41560 11980 41600
rect 12020 41560 12029 41600
rect 20039 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20425 41600
rect 0 41540 80 41560
rect 2179 41516 2237 41517
rect 1315 41476 1324 41516
rect 1364 41476 2188 41516
rect 2228 41476 2572 41516
rect 2612 41476 2621 41516
rect 2179 41475 2237 41476
rect 2668 41432 2708 41560
rect 3523 41559 3581 41560
rect 11971 41559 12029 41560
rect 13987 41516 14045 41517
rect 14851 41516 14909 41517
rect 6787 41476 6796 41516
rect 6836 41476 7660 41516
rect 7700 41476 7709 41516
rect 13315 41476 13324 41516
rect 13364 41476 13516 41516
rect 13556 41476 13996 41516
rect 14036 41476 14860 41516
rect 14900 41476 15436 41516
rect 15476 41476 15485 41516
rect 13987 41475 14045 41476
rect 14851 41475 14909 41476
rect 21424 41432 21504 41452
rect 931 41392 940 41432
rect 980 41392 2708 41432
rect 2755 41392 2764 41432
rect 2804 41392 3148 41432
rect 3188 41392 3197 41432
rect 5731 41392 5740 41432
rect 5780 41392 6220 41432
rect 6260 41392 6269 41432
rect 13411 41392 13420 41432
rect 13460 41392 13804 41432
rect 13844 41392 13853 41432
rect 19843 41392 19852 41432
rect 19892 41392 21504 41432
rect 21424 41372 21504 41392
rect 8227 41308 8236 41348
rect 8276 41308 10060 41348
rect 10100 41308 10109 41348
rect 11587 41308 11596 41348
rect 11636 41308 12076 41348
rect 12116 41308 12125 41348
rect 1795 41264 1853 41265
rect 9859 41264 9917 41265
rect 1710 41224 1804 41264
rect 1844 41224 1853 41264
rect 2851 41224 2860 41264
rect 2900 41224 3724 41264
rect 3764 41224 3773 41264
rect 8611 41224 8620 41264
rect 8660 41224 9868 41264
rect 9908 41224 9917 41264
rect 1795 41223 1853 41224
rect 9859 41223 9917 41224
rect 14083 41264 14141 41265
rect 14083 41224 14092 41264
rect 14132 41224 14476 41264
rect 14516 41224 14525 41264
rect 14083 41223 14141 41224
rect 1804 41180 1844 41223
rect 1804 41140 19276 41180
rect 19316 41140 19325 41180
rect 21424 41096 21504 41116
rect 2500 41056 4148 41096
rect 4195 41056 4204 41096
rect 4244 41056 4492 41096
rect 4532 41056 4541 41096
rect 19459 41056 19468 41096
rect 19508 41056 21504 41096
rect 355 41012 413 41013
rect 2500 41012 2540 41056
rect 4108 41012 4148 41056
rect 21424 41036 21504 41056
rect 355 40972 364 41012
rect 404 40972 2540 41012
rect 4003 40972 4012 41012
rect 4052 40972 4061 41012
rect 4108 40972 5164 41012
rect 5204 40972 5213 41012
rect 7555 40972 7564 41012
rect 7604 40972 11116 41012
rect 11156 40972 11165 41012
rect 355 40971 413 40972
rect 0 40928 80 40948
rect 4012 40928 4052 40972
rect 0 40888 4052 40928
rect 6403 40888 6412 40928
rect 6452 40888 8044 40928
rect 8084 40888 8093 40928
rect 0 40868 80 40888
rect 3679 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 4065 40844
rect 18799 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 19185 40844
rect 14467 40760 14525 40761
rect 14755 40760 14813 40761
rect 21424 40760 21504 40780
rect 4771 40720 4780 40760
rect 4820 40720 7564 40760
rect 7604 40720 7613 40760
rect 8140 40720 8812 40760
rect 8852 40720 8861 40760
rect 14467 40720 14476 40760
rect 14516 40720 14764 40760
rect 14804 40720 19372 40760
rect 19412 40720 19421 40760
rect 19555 40720 19564 40760
rect 19604 40720 21504 40760
rect 547 40676 605 40677
rect 8140 40676 8180 40720
rect 14467 40719 14525 40720
rect 14755 40719 14813 40720
rect 21424 40700 21504 40720
rect 13795 40676 13853 40677
rect 547 40636 556 40676
rect 596 40636 6796 40676
rect 6836 40636 8180 40676
rect 8227 40636 8236 40676
rect 8276 40636 11212 40676
rect 11252 40636 11261 40676
rect 13795 40636 13804 40676
rect 13844 40636 17836 40676
rect 17876 40636 17885 40676
rect 547 40635 605 40636
rect 13795 40635 13853 40636
rect 5539 40592 5597 40593
rect 3331 40552 3340 40592
rect 3380 40552 5356 40592
rect 5396 40552 5405 40592
rect 5539 40552 5548 40592
rect 5588 40552 7276 40592
rect 7316 40552 11360 40592
rect 5539 40551 5597 40552
rect 2563 40468 2572 40508
rect 2612 40468 3532 40508
rect 3572 40468 7660 40508
rect 7700 40468 7709 40508
rect 9091 40468 9100 40508
rect 9140 40468 9149 40508
rect 8899 40424 8957 40425
rect 9100 40424 9140 40468
rect 11320 40424 11360 40552
rect 12652 40552 15820 40592
rect 15860 40552 15869 40592
rect 12652 40424 12692 40552
rect 14947 40468 14956 40508
rect 14996 40468 16012 40508
rect 16052 40468 16061 40508
rect 14851 40424 14909 40425
rect 21424 40424 21504 40444
rect 835 40384 844 40424
rect 884 40384 1900 40424
rect 1940 40384 1949 40424
rect 5155 40384 5164 40424
rect 5204 40384 5644 40424
rect 5684 40384 5693 40424
rect 6019 40384 6028 40424
rect 6068 40384 6700 40424
rect 6740 40384 6749 40424
rect 8035 40384 8044 40424
rect 8084 40384 8620 40424
rect 8660 40384 8669 40424
rect 8899 40384 8908 40424
rect 8948 40384 9004 40424
rect 9044 40384 9053 40424
rect 9100 40384 10484 40424
rect 11320 40384 12652 40424
rect 12692 40384 12701 40424
rect 14766 40384 14860 40424
rect 14900 40384 14909 40424
rect 15907 40384 15916 40424
rect 15956 40384 17164 40424
rect 17204 40384 17213 40424
rect 18019 40384 18028 40424
rect 18068 40384 21504 40424
rect 8899 40383 8957 40384
rect 1795 40340 1853 40341
rect 1987 40340 2045 40341
rect 10444 40340 10484 40384
rect 14851 40383 14909 40384
rect 21424 40364 21504 40384
rect 10915 40340 10973 40341
rect 13795 40340 13853 40341
rect 1795 40300 1804 40340
rect 1844 40300 1996 40340
rect 2036 40300 2045 40340
rect 2467 40300 2476 40340
rect 2516 40300 3148 40340
rect 3188 40300 3197 40340
rect 4963 40300 4972 40340
rect 5012 40300 6316 40340
rect 6356 40300 6365 40340
rect 6595 40300 6604 40340
rect 6644 40300 9388 40340
rect 9428 40300 9437 40340
rect 10444 40300 10924 40340
rect 10964 40300 11884 40340
rect 11924 40300 11933 40340
rect 12652 40300 13804 40340
rect 13844 40300 13853 40340
rect 13987 40300 13996 40340
rect 14036 40300 15148 40340
rect 15188 40300 15197 40340
rect 1795 40299 1853 40300
rect 1987 40299 2045 40300
rect 10915 40299 10973 40300
rect 0 40256 80 40276
rect 4675 40256 4733 40257
rect 0 40216 4684 40256
rect 4724 40216 4733 40256
rect 0 40196 80 40216
rect 4675 40215 4733 40216
rect 8323 40256 8381 40257
rect 8323 40216 8332 40256
rect 8372 40216 8428 40256
rect 8468 40216 8477 40256
rect 8323 40215 8381 40216
rect 12652 40172 12692 40300
rect 13795 40299 13853 40300
rect 12931 40216 12940 40256
rect 12980 40216 14476 40256
rect 14516 40216 15052 40256
rect 15092 40216 15101 40256
rect 2500 40132 6124 40172
rect 6164 40132 6173 40172
rect 12643 40132 12652 40172
rect 12692 40132 12701 40172
rect 14659 40132 14668 40172
rect 14708 40132 14717 40172
rect 14947 40132 14956 40172
rect 14996 40132 15244 40172
rect 15284 40132 15293 40172
rect 2500 40004 2540 40132
rect 14668 40088 14708 40132
rect 21424 40088 21504 40108
rect 2659 40048 2668 40088
rect 2708 40048 3148 40088
rect 3188 40048 3197 40088
rect 4919 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 5305 40088
rect 14668 40048 15052 40088
rect 15092 40048 15101 40088
rect 20039 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20425 40088
rect 20812 40048 21504 40088
rect 20812 40004 20852 40048
rect 21424 40028 21504 40048
rect 20 39964 2540 40004
rect 5164 39964 12844 40004
rect 12884 39964 12893 40004
rect 14371 39964 14380 40004
rect 14420 39964 14668 40004
rect 14708 39964 14717 40004
rect 19171 39964 19180 40004
rect 19220 39964 20852 40004
rect 20 39752 60 39964
rect 5164 39920 5204 39964
rect 835 39880 844 39920
rect 884 39880 5204 39920
rect 11395 39880 11404 39920
rect 11444 39880 15532 39920
rect 15572 39880 15581 39920
rect 16099 39880 16108 39920
rect 16148 39880 20044 39920
rect 20084 39880 20093 39920
rect 1795 39836 1853 39837
rect 1795 39796 1804 39836
rect 1844 39796 6988 39836
rect 7028 39796 7037 39836
rect 8131 39796 8140 39836
rect 8180 39796 19564 39836
rect 19604 39796 19613 39836
rect 1795 39795 1853 39796
rect 10531 39752 10589 39753
rect 21424 39752 21504 39772
rect 20 39712 212 39752
rect 2659 39712 2668 39752
rect 2708 39712 3820 39752
rect 3860 39712 3869 39752
rect 5155 39712 5164 39752
rect 5204 39712 5740 39752
rect 5780 39712 5789 39752
rect 9955 39712 9964 39752
rect 10004 39712 10156 39752
rect 10196 39712 10540 39752
rect 10580 39712 10589 39752
rect 12163 39712 12172 39752
rect 12212 39712 12460 39752
rect 12500 39712 12509 39752
rect 14851 39712 14860 39752
rect 14900 39712 16684 39752
rect 16724 39712 17452 39752
rect 17492 39712 17501 39752
rect 19843 39712 19852 39752
rect 19892 39712 21504 39752
rect 0 39584 80 39604
rect 172 39584 212 39712
rect 10531 39711 10589 39712
rect 21424 39692 21504 39712
rect 8995 39668 9053 39669
rect 12931 39668 12989 39669
rect 16483 39668 16541 39669
rect 2275 39628 2284 39668
rect 2324 39628 4300 39668
rect 4340 39628 6508 39668
rect 6548 39628 6557 39668
rect 8995 39628 9004 39668
rect 9044 39628 9868 39668
rect 9908 39628 9917 39668
rect 12846 39628 12940 39668
rect 12980 39628 12989 39668
rect 15811 39628 15820 39668
rect 15860 39628 16108 39668
rect 16148 39628 16492 39668
rect 16532 39628 19660 39668
rect 19700 39628 19709 39668
rect 8995 39627 9053 39628
rect 12931 39627 12989 39628
rect 16483 39627 16541 39628
rect 14083 39584 14141 39585
rect 0 39544 212 39584
rect 8803 39544 8812 39584
rect 8852 39544 9100 39584
rect 9140 39544 9149 39584
rect 12547 39544 12556 39584
rect 12596 39544 14092 39584
rect 14132 39544 14141 39584
rect 0 39524 80 39544
rect 14083 39543 14141 39544
rect 6115 39460 6124 39500
rect 6164 39460 7372 39500
rect 7412 39460 7421 39500
rect 19459 39460 19468 39500
rect 19508 39460 20180 39500
rect 20140 39416 20180 39460
rect 21424 39416 21504 39436
rect 20140 39376 21504 39416
rect 21424 39356 21504 39376
rect 3679 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 4065 39332
rect 18799 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 19185 39332
rect 5923 39248 5981 39249
rect 4195 39208 4204 39248
rect 4244 39208 5932 39248
rect 5972 39208 7468 39248
rect 7508 39208 7517 39248
rect 5923 39207 5981 39208
rect 835 39164 893 39165
rect 6019 39164 6077 39165
rect 835 39124 844 39164
rect 884 39124 6028 39164
rect 6068 39124 6077 39164
rect 6883 39124 6892 39164
rect 6932 39124 7564 39164
rect 7604 39124 7613 39164
rect 14179 39124 14188 39164
rect 14228 39124 14237 39164
rect 835 39123 893 39124
rect 6019 39123 6077 39124
rect 4771 39080 4829 39081
rect 14188 39080 14228 39124
rect 21424 39080 21504 39100
rect 4099 39040 4108 39080
rect 4148 39040 4780 39080
rect 4820 39040 4829 39080
rect 5731 39040 5740 39080
rect 5780 39040 6028 39080
rect 6068 39040 6316 39080
rect 6356 39040 6365 39080
rect 6979 39040 6988 39080
rect 7028 39040 7037 39080
rect 7171 39040 7180 39080
rect 7220 39040 7948 39080
rect 7988 39040 7997 39080
rect 8803 39040 8812 39080
rect 8852 39040 10156 39080
rect 10196 39040 10205 39080
rect 12451 39040 12460 39080
rect 12500 39040 13996 39080
rect 14036 39040 14045 39080
rect 14188 39040 14668 39080
rect 14708 39040 14717 39080
rect 19843 39040 19852 39080
rect 19892 39040 21504 39080
rect 4771 39039 4829 39040
rect 6988 38996 7028 39040
rect 21424 39020 21504 39040
rect 2500 38956 4628 38996
rect 4675 38956 4684 38996
rect 4724 38956 7468 38996
rect 7508 38956 7517 38996
rect 8611 38956 8620 38996
rect 8660 38956 10252 38996
rect 10292 38956 10301 38996
rect 11320 38956 19660 38996
rect 19700 38956 19709 38996
rect 0 38912 80 38932
rect 2500 38912 2540 38956
rect 4588 38912 4628 38956
rect 11320 38912 11360 38956
rect 0 38872 2540 38912
rect 2947 38872 2956 38912
rect 2996 38872 3340 38912
rect 3380 38872 3389 38912
rect 4588 38872 5164 38912
rect 5204 38872 5213 38912
rect 5347 38872 5356 38912
rect 5396 38872 5644 38912
rect 5684 38872 11360 38912
rect 14947 38912 15005 38913
rect 16387 38912 16445 38913
rect 14947 38872 14956 38912
rect 14996 38872 16396 38912
rect 16436 38872 16445 38912
rect 0 38852 80 38872
rect 14947 38871 15005 38872
rect 16387 38871 16445 38872
rect 7372 38788 19276 38828
rect 19316 38788 19325 38828
rect 7372 38744 7412 38788
rect 21424 38744 21504 38764
rect 3043 38704 3052 38744
rect 3092 38704 3532 38744
rect 3572 38704 3581 38744
rect 6019 38704 6028 38744
rect 6068 38704 7412 38744
rect 10435 38704 10444 38744
rect 10484 38704 11692 38744
rect 11732 38704 11741 38744
rect 13411 38704 13420 38744
rect 13460 38704 14956 38744
rect 14996 38704 15724 38744
rect 15764 38704 15773 38744
rect 16291 38704 16300 38744
rect 16340 38704 16492 38744
rect 16532 38704 17260 38744
rect 17300 38704 18700 38744
rect 18740 38704 18988 38744
rect 19028 38704 19037 38744
rect 19459 38704 19468 38744
rect 19508 38704 21504 38744
rect 21424 38684 21504 38704
rect 13027 38620 13036 38660
rect 13076 38620 13900 38660
rect 13940 38620 13949 38660
rect 2563 38536 2572 38576
rect 2612 38536 3052 38576
rect 3092 38536 3101 38576
rect 4919 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 5305 38576
rect 6691 38536 6700 38576
rect 6740 38536 9676 38576
rect 9716 38536 9725 38576
rect 10243 38536 10252 38576
rect 10292 38536 11360 38576
rect 13987 38536 13996 38576
rect 14036 38536 15916 38576
rect 15956 38536 15965 38576
rect 16099 38536 16108 38576
rect 16148 38536 16300 38576
rect 16340 38536 16349 38576
rect 20039 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20425 38576
rect 163 38452 172 38492
rect 212 38452 2540 38492
rect 2500 38324 2540 38452
rect 7276 38452 10828 38492
rect 10868 38452 10877 38492
rect 7276 38408 7316 38452
rect 10723 38408 10781 38409
rect 5443 38368 5452 38408
rect 5492 38368 6604 38408
rect 6644 38368 7276 38408
rect 7316 38368 7325 38408
rect 10638 38368 10732 38408
rect 10772 38368 10781 38408
rect 11320 38408 11360 38536
rect 11971 38492 12029 38493
rect 11971 38452 11980 38492
rect 12020 38452 17644 38492
rect 17684 38452 17693 38492
rect 11971 38451 12029 38452
rect 21424 38408 21504 38428
rect 11320 38368 12076 38408
rect 12116 38368 12125 38408
rect 14659 38368 14668 38408
rect 14708 38368 16436 38408
rect 19459 38368 19468 38408
rect 19508 38368 21504 38408
rect 10723 38367 10781 38368
rect 12739 38324 12797 38325
rect 2500 38284 12748 38324
rect 12788 38284 12797 38324
rect 12739 38283 12797 38284
rect 0 38240 80 38260
rect 3139 38240 3197 38241
rect 10243 38240 10301 38241
rect 0 38200 3148 38240
rect 3188 38200 3197 38240
rect 3331 38200 3340 38240
rect 3380 38200 6316 38240
rect 6356 38200 6365 38240
rect 7555 38200 7564 38240
rect 7604 38200 8140 38240
rect 8180 38200 8189 38240
rect 8899 38200 8908 38240
rect 8948 38200 9676 38240
rect 9716 38200 9725 38240
rect 10158 38200 10252 38240
rect 10292 38200 10301 38240
rect 0 38180 80 38200
rect 3139 38199 3197 38200
rect 10243 38199 10301 38200
rect 11107 38240 11165 38241
rect 13315 38240 13373 38241
rect 14755 38240 14813 38241
rect 16396 38240 16436 38368
rect 21424 38348 21504 38368
rect 11107 38200 11116 38240
rect 11156 38200 11212 38240
rect 11252 38200 11261 38240
rect 13230 38200 13324 38240
rect 13364 38200 13373 38240
rect 13987 38200 13996 38240
rect 14036 38200 14612 38240
rect 14659 38200 14668 38240
rect 14708 38200 14764 38240
rect 14804 38200 14813 38240
rect 16387 38200 16396 38240
rect 16436 38200 16445 38240
rect 11107 38199 11165 38200
rect 13315 38199 13373 38200
rect 10627 38156 10685 38157
rect 14083 38156 14141 38157
rect 14572 38156 14612 38200
rect 14755 38199 14813 38200
rect 18307 38156 18365 38157
rect 19843 38156 19901 38157
rect 3619 38116 3628 38156
rect 3668 38116 4052 38156
rect 5443 38116 5452 38156
rect 5492 38116 5836 38156
rect 5876 38116 5885 38156
rect 10542 38116 10636 38156
rect 10676 38116 10685 38156
rect 12835 38116 12844 38156
rect 12884 38116 13420 38156
rect 13460 38116 13469 38156
rect 14083 38116 14092 38156
rect 14132 38116 14476 38156
rect 14516 38116 14525 38156
rect 14572 38116 15340 38156
rect 15380 38116 16492 38156
rect 16532 38116 16541 38156
rect 18307 38116 18316 38156
rect 18356 38116 18604 38156
rect 18644 38116 18653 38156
rect 19267 38116 19276 38156
rect 19316 38116 19325 38156
rect 19843 38116 19852 38156
rect 19892 38116 20044 38156
rect 20084 38116 20093 38156
rect 4012 38072 4052 38116
rect 10627 38115 10685 38116
rect 14083 38115 14141 38116
rect 18307 38115 18365 38116
rect 4291 38072 4349 38073
rect 4003 38032 4012 38072
rect 4052 38032 4300 38072
rect 4340 38032 6700 38072
rect 6740 38032 6749 38072
rect 11875 38032 11884 38072
rect 11924 38032 18220 38072
rect 18260 38032 18269 38072
rect 4291 38031 4349 38032
rect 11971 37988 12029 37989
rect 19276 37988 19316 38116
rect 19843 38115 19901 38116
rect 21424 38072 21504 38092
rect 20227 38032 20236 38072
rect 20276 38032 21504 38072
rect 21424 38012 21504 38032
rect 4099 37948 4108 37988
rect 4148 37948 4492 37988
rect 4532 37948 4541 37988
rect 7267 37948 7276 37988
rect 7316 37948 8140 37988
rect 8180 37948 8189 37988
rect 10723 37948 10732 37988
rect 10772 37948 11980 37988
rect 12020 37948 12029 37988
rect 11971 37947 12029 37948
rect 12076 37948 19316 37988
rect 19555 37988 19613 37989
rect 19555 37948 19564 37988
rect 19604 37948 19852 37988
rect 19892 37948 19901 37988
rect 1219 37864 1228 37904
rect 1268 37864 6508 37904
rect 6548 37864 6557 37904
rect 3679 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 4065 37820
rect 12076 37736 12116 37948
rect 19555 37947 19613 37948
rect 15811 37904 15869 37905
rect 13315 37864 13324 37904
rect 13364 37864 13940 37904
rect 12739 37820 12797 37821
rect 12654 37780 12748 37820
rect 12788 37780 12797 37820
rect 12739 37779 12797 37780
rect 2083 37696 2092 37736
rect 2132 37696 5932 37736
rect 5972 37696 5981 37736
rect 7651 37696 7660 37736
rect 7700 37696 12116 37736
rect 13900 37736 13940 37864
rect 14188 37864 14572 37904
rect 14612 37864 14621 37904
rect 15726 37864 15820 37904
rect 15860 37864 15869 37904
rect 18211 37864 18220 37904
rect 18260 37864 18604 37904
rect 18644 37864 18653 37904
rect 14188 37820 14228 37864
rect 15811 37863 15869 37864
rect 15139 37820 15197 37821
rect 14179 37780 14188 37820
rect 14228 37780 14237 37820
rect 15054 37780 15148 37820
rect 15188 37780 15197 37820
rect 18799 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 19185 37820
rect 15139 37779 15197 37780
rect 21424 37736 21504 37756
rect 13900 37696 14284 37736
rect 14324 37696 15436 37736
rect 15476 37696 15820 37736
rect 15860 37696 16300 37736
rect 16340 37696 16349 37736
rect 18691 37696 18700 37736
rect 18740 37696 21504 37736
rect 21424 37676 21504 37696
rect 12739 37652 12797 37653
rect 15139 37652 15197 37653
rect 5539 37612 5548 37652
rect 5588 37612 6220 37652
rect 6260 37612 6269 37652
rect 7171 37612 7180 37652
rect 7220 37612 7756 37652
rect 7796 37612 7805 37652
rect 8803 37612 8812 37652
rect 8852 37612 10924 37652
rect 10964 37612 10973 37652
rect 12739 37612 12748 37652
rect 12788 37612 14860 37652
rect 14900 37612 14909 37652
rect 15139 37612 15148 37652
rect 15188 37612 15916 37652
rect 15956 37612 15965 37652
rect 12739 37611 12797 37612
rect 0 37568 80 37588
rect 14860 37568 14900 37612
rect 15139 37611 15197 37612
rect 0 37528 1708 37568
rect 1748 37528 1757 37568
rect 14860 37528 15436 37568
rect 15476 37528 15485 37568
rect 0 37508 80 37528
rect 7939 37444 7948 37484
rect 7988 37444 19276 37484
rect 19316 37444 19325 37484
rect 20035 37444 20044 37484
rect 20084 37444 20093 37484
rect 7267 37400 7325 37401
rect 20044 37400 20084 37444
rect 21424 37400 21504 37420
rect 2371 37360 2380 37400
rect 2420 37360 3724 37400
rect 3764 37360 4588 37400
rect 4628 37360 4637 37400
rect 5347 37360 5356 37400
rect 5396 37360 6988 37400
rect 7028 37360 7276 37400
rect 7316 37360 7325 37400
rect 9187 37360 9196 37400
rect 9236 37360 9388 37400
rect 9428 37360 9437 37400
rect 11875 37360 11884 37400
rect 11924 37360 13516 37400
rect 13556 37360 13565 37400
rect 14179 37360 14188 37400
rect 14228 37360 20084 37400
rect 20227 37360 20236 37400
rect 20276 37360 21504 37400
rect 7267 37359 7325 37360
rect 12259 37316 12317 37317
rect 14188 37316 14228 37360
rect 21424 37340 21504 37360
rect 643 37276 652 37316
rect 692 37276 11360 37316
rect 11779 37276 11788 37316
rect 11828 37276 12172 37316
rect 12212 37276 12268 37316
rect 12308 37276 12317 37316
rect 12835 37276 12844 37316
rect 12884 37276 14228 37316
rect 17059 37276 17068 37316
rect 17108 37276 19660 37316
rect 19700 37276 19709 37316
rect 1891 37232 1949 37233
rect 4099 37232 4157 37233
rect 11320 37232 11360 37276
rect 12259 37275 12317 37276
rect 1315 37192 1324 37232
rect 1364 37192 1900 37232
rect 1940 37192 2540 37232
rect 4014 37192 4108 37232
rect 4148 37192 5260 37232
rect 5300 37192 5309 37232
rect 11320 37192 16588 37232
rect 16628 37192 16637 37232
rect 1891 37191 1949 37192
rect 2500 37148 2540 37192
rect 4099 37191 4157 37192
rect 2500 37108 5740 37148
rect 5780 37108 7372 37148
rect 7412 37108 11212 37148
rect 11252 37108 19372 37148
rect 19412 37108 19421 37148
rect 21424 37064 21504 37084
rect 3427 37024 3436 37064
rect 3476 37024 3628 37064
rect 3668 37024 3677 37064
rect 4919 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 5305 37064
rect 20039 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20425 37064
rect 20524 37024 21504 37064
rect 1507 36980 1565 36981
rect 5635 36980 5693 36981
rect 6595 36980 6653 36981
rect 20524 36980 20564 37024
rect 21424 37004 21504 37024
rect 1507 36940 1516 36980
rect 1556 36940 2476 36980
rect 2516 36940 5548 36980
rect 5588 36940 5644 36980
rect 5684 36940 5712 36980
rect 6499 36940 6508 36980
rect 6548 36940 6604 36980
rect 6644 36940 6653 36980
rect 13411 36940 13420 36980
rect 13460 36940 13804 36980
rect 13844 36940 13853 36980
rect 16963 36940 16972 36980
rect 17012 36940 17548 36980
rect 17588 36940 17597 36980
rect 19747 36940 19756 36980
rect 19796 36940 20564 36980
rect 1507 36939 1565 36940
rect 5635 36939 5693 36940
rect 6595 36939 6653 36940
rect 0 36896 80 36916
rect 7075 36896 7133 36897
rect 0 36856 1996 36896
rect 2036 36856 2045 36896
rect 2659 36856 2668 36896
rect 2708 36856 3532 36896
rect 3572 36856 3581 36896
rect 6787 36856 6796 36896
rect 6836 36856 7084 36896
rect 7124 36856 7133 36896
rect 10723 36856 10732 36896
rect 10772 36856 11020 36896
rect 11060 36856 11069 36896
rect 11320 36856 18124 36896
rect 18164 36856 18173 36896
rect 0 36836 80 36856
rect 7075 36855 7133 36856
rect 5635 36812 5693 36813
rect 11320 36812 11360 36856
rect 5635 36772 5644 36812
rect 5684 36772 11360 36812
rect 11491 36772 11500 36812
rect 11540 36772 16588 36812
rect 16628 36772 16637 36812
rect 16963 36772 16972 36812
rect 17012 36772 18220 36812
rect 18260 36772 18269 36812
rect 5635 36771 5693 36772
rect 1123 36728 1181 36729
rect 9763 36728 9821 36729
rect 21424 36728 21504 36748
rect 1104 36688 1132 36728
rect 1172 36688 1228 36728
rect 1268 36688 1516 36728
rect 1556 36688 1565 36728
rect 6787 36688 6796 36728
rect 6836 36688 7084 36728
rect 7124 36688 7133 36728
rect 9678 36688 9772 36728
rect 9812 36688 9821 36728
rect 10339 36688 10348 36728
rect 10388 36688 11020 36728
rect 11060 36688 11069 36728
rect 12739 36688 12748 36728
rect 12788 36688 14092 36728
rect 14132 36688 14141 36728
rect 15427 36688 15436 36728
rect 15476 36688 15724 36728
rect 15764 36688 15773 36728
rect 20131 36688 20140 36728
rect 20180 36688 21504 36728
rect 1123 36687 1181 36688
rect 9763 36687 9821 36688
rect 21424 36668 21504 36688
rect 12739 36644 12797 36645
rect 67 36604 76 36644
rect 116 36604 3340 36644
rect 3380 36604 3389 36644
rect 6115 36604 6124 36644
rect 6164 36604 11500 36644
rect 11540 36604 11549 36644
rect 12739 36604 12748 36644
rect 12788 36604 13708 36644
rect 13748 36604 13757 36644
rect 15907 36604 15916 36644
rect 15956 36604 17068 36644
rect 17108 36604 17117 36644
rect 12739 36603 12797 36604
rect 10051 36560 10109 36561
rect 4867 36520 4876 36560
rect 4916 36520 6988 36560
rect 7028 36520 8332 36560
rect 8372 36520 8381 36560
rect 8803 36520 8812 36560
rect 8852 36520 9388 36560
rect 9428 36520 9868 36560
rect 9908 36520 9917 36560
rect 9966 36520 10060 36560
rect 10100 36520 10109 36560
rect 10051 36519 10109 36520
rect 10723 36560 10781 36561
rect 13219 36560 13277 36561
rect 10723 36520 10732 36560
rect 10772 36520 10924 36560
rect 10964 36520 10973 36560
rect 12355 36520 12364 36560
rect 12404 36520 13228 36560
rect 13268 36520 13324 36560
rect 13364 36520 14380 36560
rect 14420 36520 15340 36560
rect 15380 36520 15389 36560
rect 16387 36520 16396 36560
rect 16436 36520 16972 36560
rect 17012 36520 17021 36560
rect 10723 36519 10781 36520
rect 13219 36519 13277 36520
rect 931 36476 989 36477
rect 6211 36476 6269 36477
rect 13027 36476 13085 36477
rect 15811 36476 15869 36477
rect 931 36436 940 36476
rect 980 36436 6220 36476
rect 6260 36436 6269 36476
rect 11299 36436 11308 36476
rect 11348 36436 11500 36476
rect 11540 36436 11549 36476
rect 13027 36436 13036 36476
rect 13076 36436 13228 36476
rect 13268 36436 13277 36476
rect 15715 36436 15724 36476
rect 15764 36436 15820 36476
rect 15860 36436 15869 36476
rect 931 36435 989 36436
rect 6211 36435 6269 36436
rect 13027 36435 13085 36436
rect 15811 36435 15869 36436
rect 10819 36392 10877 36393
rect 3331 36352 3340 36392
rect 3380 36352 10828 36392
rect 10868 36352 10877 36392
rect 0 36224 80 36244
rect 0 36184 3148 36224
rect 3188 36184 3197 36224
rect 0 36164 80 36184
rect 3532 36140 3572 36352
rect 10819 36351 10877 36352
rect 19651 36392 19709 36393
rect 21424 36392 21504 36412
rect 19651 36352 19660 36392
rect 19700 36352 21504 36392
rect 19651 36351 19709 36352
rect 21424 36332 21504 36352
rect 11779 36308 11837 36309
rect 19459 36308 19517 36309
rect 3679 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 4065 36308
rect 11683 36268 11692 36308
rect 11732 36268 11788 36308
rect 11828 36268 11837 36308
rect 18799 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 19185 36308
rect 19374 36268 19468 36308
rect 19508 36268 19517 36308
rect 11779 36267 11837 36268
rect 19459 36267 19517 36268
rect 6595 36224 6653 36225
rect 6595 36184 6604 36224
rect 6644 36184 7372 36224
rect 7412 36184 7421 36224
rect 11299 36184 11308 36224
rect 11348 36184 11980 36224
rect 12020 36184 12029 36224
rect 14188 36184 19948 36224
rect 19988 36184 19997 36224
rect 6595 36183 6653 36184
rect 4291 36140 4349 36141
rect 7171 36140 7229 36141
rect 3532 36100 3724 36140
rect 3764 36100 3773 36140
rect 4003 36100 4012 36140
rect 4052 36100 4300 36140
rect 4340 36100 4349 36140
rect 7086 36100 7180 36140
rect 7220 36100 7229 36140
rect 4291 36099 4349 36100
rect 7171 36099 7229 36100
rect 9667 36140 9725 36141
rect 14188 36140 14228 36184
rect 19843 36140 19901 36141
rect 9667 36100 9676 36140
rect 9716 36100 14228 36140
rect 14275 36100 14284 36140
rect 14324 36100 15244 36140
rect 15284 36100 15293 36140
rect 18979 36100 18988 36140
rect 19028 36100 19852 36140
rect 19892 36100 19901 36140
rect 9667 36099 9725 36100
rect 19843 36099 19901 36100
rect 12643 36056 12701 36057
rect 17347 36056 17405 36057
rect 21424 36056 21504 36076
rect 1987 36016 1996 36056
rect 2036 36016 7372 36056
rect 7412 36016 7421 36056
rect 8803 36016 8812 36056
rect 8852 36016 9196 36056
rect 9236 36016 12172 36056
rect 12212 36016 12221 36056
rect 12643 36016 12652 36056
rect 12692 36016 17356 36056
rect 17396 36016 19604 36056
rect 20035 36016 20044 36056
rect 20084 36016 21504 36056
rect 12643 36015 12701 36016
rect 17347 36015 17405 36016
rect 19564 35972 19604 36016
rect 21424 35996 21504 36016
rect 2467 35932 2476 35972
rect 2516 35932 3340 35972
rect 3380 35932 8620 35972
rect 8660 35932 8669 35972
rect 10531 35932 10540 35972
rect 10580 35932 11404 35972
rect 11444 35932 11692 35972
rect 11732 35932 11741 35972
rect 14947 35932 14956 35972
rect 14996 35932 15820 35972
rect 15860 35932 18124 35972
rect 18164 35932 18173 35972
rect 19555 35932 19564 35972
rect 19604 35932 19613 35972
rect 9091 35888 9149 35889
rect 2500 35848 9100 35888
rect 9140 35848 9676 35888
rect 9716 35848 9725 35888
rect 10051 35848 10060 35888
rect 10100 35848 11980 35888
rect 12020 35848 12029 35888
rect 17347 35848 17356 35888
rect 17396 35848 17740 35888
rect 17780 35848 17789 35888
rect 739 35804 797 35805
rect 2500 35804 2540 35848
rect 9091 35847 9149 35848
rect 739 35764 748 35804
rect 788 35764 2540 35804
rect 9475 35804 9533 35805
rect 10819 35804 10877 35805
rect 9475 35764 9484 35804
rect 9524 35764 9772 35804
rect 9812 35764 9821 35804
rect 10819 35764 10828 35804
rect 10868 35764 19852 35804
rect 19892 35764 19901 35804
rect 739 35763 797 35764
rect 9475 35763 9533 35764
rect 10819 35763 10877 35764
rect 18307 35720 18365 35721
rect 21424 35720 21504 35740
rect 10339 35680 10348 35720
rect 10388 35680 12652 35720
rect 12692 35680 12701 35720
rect 16579 35680 16588 35720
rect 16628 35680 18316 35720
rect 18356 35680 18365 35720
rect 19747 35680 19756 35720
rect 19796 35680 21504 35720
rect 18307 35679 18365 35680
rect 21424 35660 21504 35680
rect 7363 35596 7372 35636
rect 7412 35596 19852 35636
rect 19892 35596 19901 35636
rect 0 35552 80 35572
rect 0 35512 76 35552
rect 116 35512 125 35552
rect 4919 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 5305 35552
rect 6124 35512 10156 35552
rect 10196 35512 10205 35552
rect 11491 35512 11500 35552
rect 11540 35512 12460 35552
rect 12500 35512 12509 35552
rect 20039 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20425 35552
rect 0 35492 80 35512
rect 6124 35468 6164 35512
rect 1219 35428 1228 35468
rect 1268 35428 6164 35468
rect 6211 35468 6269 35469
rect 6211 35428 6220 35468
rect 6260 35428 10732 35468
rect 10772 35428 10781 35468
rect 11779 35428 11788 35468
rect 11828 35428 12652 35468
rect 12692 35428 12701 35468
rect 6211 35427 6269 35428
rect 7267 35384 7325 35385
rect 20707 35384 20765 35385
rect 21424 35384 21504 35404
rect 5827 35344 5836 35384
rect 5876 35344 5885 35384
rect 6979 35344 6988 35384
rect 7028 35344 7276 35384
rect 7316 35344 7325 35384
rect 15235 35344 15244 35384
rect 15284 35344 16684 35384
rect 16724 35344 17740 35384
rect 17780 35344 17789 35384
rect 19171 35344 19180 35384
rect 19220 35344 20524 35384
rect 20564 35344 20573 35384
rect 20707 35344 20716 35384
rect 20756 35344 21504 35384
rect 5836 35301 5876 35344
rect 7267 35343 7325 35344
rect 20707 35343 20765 35344
rect 21424 35324 21504 35344
rect 5827 35300 5885 35301
rect 7075 35300 7133 35301
rect 16099 35300 16157 35301
rect 16675 35300 16733 35301
rect 18307 35300 18365 35301
rect 3043 35260 3052 35300
rect 3092 35260 3101 35300
rect 5796 35260 5836 35300
rect 5876 35260 5885 35300
rect 6211 35260 6220 35300
rect 6260 35260 6269 35300
rect 7075 35260 7084 35300
rect 7124 35260 8236 35300
rect 8276 35260 8620 35300
rect 8660 35260 9772 35300
rect 9812 35260 9821 35300
rect 15427 35260 15436 35300
rect 15476 35260 15628 35300
rect 15668 35260 15677 35300
rect 16099 35260 16108 35300
rect 16148 35260 16684 35300
rect 16724 35260 16733 35300
rect 18222 35260 18316 35300
rect 18356 35260 18365 35300
rect 2947 35216 3005 35217
rect 3052 35216 3092 35260
rect 5827 35259 5885 35260
rect 6220 35216 6260 35260
rect 7075 35259 7133 35260
rect 16099 35259 16157 35260
rect 16675 35259 16733 35260
rect 18307 35259 18365 35260
rect 2659 35176 2668 35216
rect 2708 35176 2956 35216
rect 2996 35176 3092 35216
rect 3619 35176 3628 35216
rect 3668 35176 4012 35216
rect 4052 35176 4061 35216
rect 5836 35176 6260 35216
rect 6691 35176 6700 35216
rect 6740 35176 7372 35216
rect 7412 35176 7852 35216
rect 7892 35176 7901 35216
rect 9091 35176 9100 35216
rect 9140 35176 9868 35216
rect 9908 35176 9917 35216
rect 10243 35176 10252 35216
rect 10292 35176 12172 35216
rect 12212 35176 12221 35216
rect 14083 35176 14092 35216
rect 14132 35176 14380 35216
rect 14420 35176 16204 35216
rect 16244 35176 16253 35216
rect 2947 35175 3005 35176
rect 3139 35132 3197 35133
rect 3043 35092 3052 35132
rect 3092 35092 3148 35132
rect 3188 35092 3436 35132
rect 3476 35092 3485 35132
rect 3139 35091 3197 35092
rect 5836 35049 5876 35176
rect 18019 35132 18077 35133
rect 9187 35092 9196 35132
rect 9236 35092 12076 35132
rect 12116 35092 12125 35132
rect 13123 35092 13132 35132
rect 13172 35092 18028 35132
rect 18068 35092 18988 35132
rect 19028 35092 19037 35132
rect 2755 35048 2813 35049
rect 4483 35048 4541 35049
rect 2755 35008 2764 35048
rect 2804 35008 3148 35048
rect 3188 35008 3532 35048
rect 3572 35008 3581 35048
rect 4398 35008 4492 35048
rect 4532 35008 4541 35048
rect 2755 35007 2813 35008
rect 4483 35007 4541 35008
rect 5827 35048 5885 35049
rect 8227 35048 8285 35049
rect 13132 35048 13172 35092
rect 18019 35091 18077 35092
rect 15043 35048 15101 35049
rect 19651 35048 19709 35049
rect 5827 35008 5836 35048
rect 5876 35008 5885 35048
rect 8142 35008 8236 35048
rect 8276 35008 9676 35048
rect 9716 35008 9725 35048
rect 9859 35008 9868 35048
rect 9908 35008 13172 35048
rect 13603 35008 13612 35048
rect 13652 35008 14956 35048
rect 14996 35008 15052 35048
rect 15092 35008 15101 35048
rect 15619 35008 15628 35048
rect 15668 35008 17260 35048
rect 17300 35008 17309 35048
rect 19566 35008 19660 35048
rect 19700 35008 19709 35048
rect 5827 35007 5885 35008
rect 8227 35007 8285 35008
rect 3523 34964 3581 34965
rect 5539 34964 5597 34965
rect 9676 34964 9716 35008
rect 15043 35007 15101 35008
rect 19651 35007 19709 35008
rect 19939 35048 19997 35049
rect 21424 35048 21504 35068
rect 19939 35008 19948 35048
rect 19988 35008 21504 35048
rect 19939 35007 19997 35008
rect 21424 34988 21504 35008
rect 11395 34964 11453 34965
rect 1891 34924 1900 34964
rect 1940 34924 1949 34964
rect 3523 34924 3532 34964
rect 3572 34924 3724 34964
rect 3764 34924 3773 34964
rect 5059 34924 5068 34964
rect 5108 34924 5548 34964
rect 5588 34924 5597 34964
rect 7843 34924 7852 34964
rect 7892 34924 8524 34964
rect 8564 34924 8573 34964
rect 9676 34924 10444 34964
rect 10484 34924 10493 34964
rect 11395 34924 11404 34964
rect 11444 34924 11692 34964
rect 11732 34924 11741 34964
rect 11971 34924 11980 34964
rect 12020 34924 12364 34964
rect 12404 34924 12413 34964
rect 12835 34924 12844 34964
rect 12884 34924 13228 34964
rect 13268 34924 13277 34964
rect 0 34880 80 34900
rect 1900 34880 1940 34924
rect 3523 34923 3581 34924
rect 5539 34923 5597 34924
rect 11395 34923 11453 34924
rect 15331 34880 15389 34881
rect 0 34840 1940 34880
rect 5443 34840 5452 34880
rect 5492 34840 5932 34880
rect 5972 34840 10348 34880
rect 10388 34840 10397 34880
rect 10723 34840 10732 34880
rect 10772 34840 15340 34880
rect 15380 34840 16684 34880
rect 16724 34840 16733 34880
rect 0 34820 80 34840
rect 15331 34839 15389 34840
rect 1699 34796 1757 34797
rect 5347 34796 5405 34797
rect 10339 34796 10397 34797
rect 1699 34756 1708 34796
rect 1748 34756 2540 34796
rect 3679 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 4065 34796
rect 5347 34756 5356 34796
rect 5396 34756 6892 34796
rect 6932 34756 6941 34796
rect 9667 34756 9676 34796
rect 9716 34756 9964 34796
rect 10004 34756 10013 34796
rect 10339 34756 10348 34796
rect 10388 34756 11212 34796
rect 11252 34756 11261 34796
rect 11320 34756 15476 34796
rect 18799 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 19185 34796
rect 1699 34755 1757 34756
rect 2500 34712 2540 34756
rect 5347 34755 5405 34756
rect 10339 34755 10397 34756
rect 5539 34712 5597 34713
rect 6595 34712 6653 34713
rect 11320 34712 11360 34756
rect 15436 34712 15476 34756
rect 21424 34712 21504 34732
rect 2500 34672 5260 34712
rect 5300 34672 5309 34712
rect 5539 34672 5548 34712
rect 5588 34672 6548 34712
rect 5539 34671 5597 34672
rect 2371 34628 2429 34629
rect 6508 34628 6548 34672
rect 6595 34672 6604 34712
rect 6644 34672 11360 34712
rect 11971 34672 11980 34712
rect 12020 34672 12268 34712
rect 12308 34672 12317 34712
rect 15436 34672 19468 34712
rect 19508 34672 19517 34712
rect 20140 34672 21504 34712
rect 6595 34671 6653 34672
rect 11779 34628 11837 34629
rect 13123 34628 13181 34629
rect 20140 34628 20180 34672
rect 21424 34652 21504 34672
rect 2371 34588 2380 34628
rect 2420 34588 6124 34628
rect 6164 34588 6173 34628
rect 6508 34588 6796 34628
rect 6836 34588 6845 34628
rect 8515 34588 8524 34628
rect 8564 34588 11788 34628
rect 11828 34588 13132 34628
rect 13172 34588 13181 34628
rect 16867 34588 16876 34628
rect 16916 34588 20180 34628
rect 2371 34587 2429 34588
rect 11779 34587 11837 34588
rect 13123 34587 13181 34588
rect 5539 34544 5597 34545
rect 6019 34544 6077 34545
rect 17443 34544 17501 34545
rect 5539 34504 5548 34544
rect 5588 34504 5740 34544
rect 5780 34504 5789 34544
rect 5934 34504 6028 34544
rect 6068 34504 6077 34544
rect 6403 34504 6412 34544
rect 6452 34504 6700 34544
rect 6740 34504 6749 34544
rect 7363 34504 7372 34544
rect 7412 34504 9772 34544
rect 9812 34504 11404 34544
rect 11444 34504 11692 34544
rect 11732 34504 11741 34544
rect 15052 34504 15436 34544
rect 15476 34504 15485 34544
rect 17443 34504 17452 34544
rect 17492 34504 17548 34544
rect 17588 34504 17597 34544
rect 19363 34504 19372 34544
rect 19412 34504 19421 34544
rect 5539 34503 5597 34504
rect 6019 34503 6077 34504
rect 6211 34460 6269 34461
rect 11107 34460 11165 34461
rect 15052 34460 15092 34504
rect 17443 34503 17501 34504
rect 1411 34420 1420 34460
rect 1460 34420 4300 34460
rect 4340 34420 4349 34460
rect 5251 34420 5260 34460
rect 5300 34420 6124 34460
rect 6164 34420 6220 34460
rect 6260 34420 6288 34460
rect 9379 34420 9388 34460
rect 9428 34420 9964 34460
rect 10004 34420 10252 34460
rect 10292 34420 10636 34460
rect 10676 34420 10685 34460
rect 11107 34420 11116 34460
rect 11156 34420 12940 34460
rect 12980 34420 12989 34460
rect 13699 34420 13708 34460
rect 13748 34420 15052 34460
rect 15092 34420 15101 34460
rect 16675 34420 16684 34460
rect 16724 34420 17164 34460
rect 17204 34420 17213 34460
rect 6211 34419 6269 34420
rect 11107 34419 11165 34420
rect 1315 34376 1373 34377
rect 10723 34376 10781 34377
rect 12835 34376 12893 34377
rect 1219 34336 1228 34376
rect 1268 34336 1324 34376
rect 1364 34336 1373 34376
rect 3043 34336 3052 34376
rect 3092 34336 4588 34376
rect 4628 34336 5740 34376
rect 5780 34336 6604 34376
rect 6644 34336 6653 34376
rect 7747 34336 7756 34376
rect 7796 34336 9580 34376
rect 9620 34336 9629 34376
rect 10638 34336 10732 34376
rect 10772 34336 10781 34376
rect 12739 34336 12748 34376
rect 12788 34336 12844 34376
rect 12884 34336 12893 34376
rect 14947 34336 14956 34376
rect 14996 34336 15916 34376
rect 15956 34336 15965 34376
rect 16963 34336 16972 34376
rect 17012 34336 18124 34376
rect 18164 34336 18173 34376
rect 1315 34335 1373 34336
rect 10723 34335 10781 34336
rect 12835 34335 12893 34336
rect 7651 34292 7709 34293
rect 19372 34292 19412 34504
rect 21424 34376 21504 34396
rect 20140 34336 21504 34376
rect 20140 34292 20180 34336
rect 21424 34316 21504 34336
rect 4483 34252 4492 34292
rect 4532 34252 6700 34292
rect 6740 34252 6749 34292
rect 7566 34252 7660 34292
rect 7700 34252 7709 34292
rect 9379 34252 9388 34292
rect 9428 34252 19412 34292
rect 19651 34252 19660 34292
rect 19700 34252 20180 34292
rect 7651 34251 7709 34252
rect 0 34208 80 34228
rect 12355 34208 12413 34209
rect 19843 34208 19901 34209
rect 0 34168 2764 34208
rect 2804 34168 2813 34208
rect 5539 34168 5548 34208
rect 5588 34168 6412 34208
rect 6452 34168 6461 34208
rect 6883 34168 6892 34208
rect 6932 34168 10636 34208
rect 10676 34168 11212 34208
rect 11252 34168 11261 34208
rect 11320 34168 11924 34208
rect 12270 34168 12364 34208
rect 12404 34168 12413 34208
rect 13987 34168 13996 34208
rect 14036 34168 14572 34208
rect 14612 34168 17644 34208
rect 17684 34168 17693 34208
rect 19843 34168 19852 34208
rect 19892 34168 20044 34208
rect 20084 34168 20093 34208
rect 0 34148 80 34168
rect 2851 34124 2909 34125
rect 11320 34124 11360 34168
rect 2851 34084 2860 34124
rect 2900 34084 3244 34124
rect 3284 34084 3293 34124
rect 4291 34084 4300 34124
rect 4340 34084 7756 34124
rect 7796 34084 7805 34124
rect 8035 34084 8044 34124
rect 8084 34084 9196 34124
rect 9236 34084 9484 34124
rect 9524 34084 9533 34124
rect 10147 34084 10156 34124
rect 10196 34084 11360 34124
rect 11884 34124 11924 34168
rect 12355 34167 12413 34168
rect 19843 34167 19901 34168
rect 11884 34084 12460 34124
rect 12500 34084 12509 34124
rect 14083 34084 14092 34124
rect 14132 34084 14141 34124
rect 17539 34084 17548 34124
rect 17588 34084 18028 34124
rect 18068 34084 18077 34124
rect 19843 34084 19852 34124
rect 19892 34084 20564 34124
rect 2851 34083 2909 34084
rect 1315 34040 1373 34041
rect 2083 34040 2141 34041
rect 14092 34040 14132 34084
rect 20524 34040 20564 34084
rect 21424 34040 21504 34060
rect 1315 34000 1324 34040
rect 1364 34000 2092 34040
rect 2132 34000 4492 34040
rect 4532 34000 4541 34040
rect 4919 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 5305 34040
rect 5635 34000 5644 34040
rect 5684 34000 9772 34040
rect 9812 34000 9821 34040
rect 10051 34000 10060 34040
rect 10100 34000 12212 34040
rect 12259 34000 12268 34040
rect 12308 34000 12748 34040
rect 12788 34000 12797 34040
rect 13996 34000 14132 34040
rect 20039 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20425 34040
rect 20524 34000 21504 34040
rect 1315 33999 1373 34000
rect 2083 33999 2141 34000
rect 10339 33956 10397 33957
rect 3043 33916 3052 33956
rect 3092 33916 4204 33956
rect 4244 33916 4253 33956
rect 5443 33916 5452 33956
rect 5492 33916 5932 33956
rect 5972 33916 5981 33956
rect 10254 33916 10348 33956
rect 10388 33916 10397 33956
rect 12172 33956 12212 34000
rect 12172 33916 12556 33956
rect 12596 33916 12605 33956
rect 10339 33915 10397 33916
rect 3235 33872 3293 33873
rect 13996 33872 14036 34000
rect 21424 33980 21504 34000
rect 20707 33956 20765 33957
rect 14083 33916 14092 33956
rect 14132 33916 15244 33956
rect 15284 33916 15293 33956
rect 19267 33916 19276 33956
rect 19316 33916 19325 33956
rect 19555 33916 19564 33956
rect 19604 33916 20716 33956
rect 20756 33916 20765 33956
rect 2947 33832 2956 33872
rect 2996 33832 3005 33872
rect 3150 33832 3244 33872
rect 3284 33832 3293 33872
rect 4387 33832 4396 33872
rect 4436 33832 7660 33872
rect 7700 33832 7709 33872
rect 11395 33832 11404 33872
rect 11444 33832 15724 33872
rect 15764 33832 15773 33872
rect 17731 33832 17740 33872
rect 17780 33832 18604 33872
rect 18644 33832 18653 33872
rect 2956 33788 2996 33832
rect 3235 33831 3293 33832
rect 8131 33788 8189 33789
rect 18115 33788 18173 33789
rect 19276 33788 19316 33916
rect 20707 33915 20765 33916
rect 19939 33872 19997 33873
rect 19854 33832 19948 33872
rect 19988 33832 19997 33872
rect 19939 33831 19997 33832
rect 739 33748 748 33788
rect 788 33748 1036 33788
rect 1076 33748 1085 33788
rect 2956 33748 3436 33788
rect 3476 33748 3485 33788
rect 5155 33748 5164 33788
rect 5204 33748 6124 33788
rect 6164 33748 6173 33788
rect 7555 33748 7564 33788
rect 7604 33748 8140 33788
rect 8180 33748 8189 33788
rect 11779 33748 11788 33788
rect 11828 33748 12364 33788
rect 12404 33748 12413 33788
rect 12931 33748 12940 33788
rect 12980 33748 12989 33788
rect 18115 33748 18124 33788
rect 18164 33748 18220 33788
rect 18260 33748 18269 33788
rect 19276 33748 20044 33788
rect 20084 33748 20093 33788
rect 8131 33747 8189 33748
rect 3427 33704 3485 33705
rect 10819 33704 10877 33705
rect 2947 33664 2956 33704
rect 2996 33664 3436 33704
rect 3476 33664 3485 33704
rect 3907 33664 3916 33704
rect 3956 33664 4204 33704
rect 4244 33664 6892 33704
rect 6932 33664 6941 33704
rect 8803 33664 8812 33704
rect 8852 33664 9004 33704
rect 9044 33664 9053 33704
rect 10734 33664 10828 33704
rect 10868 33664 10877 33704
rect 3427 33663 3485 33664
rect 10819 33663 10877 33664
rect 4291 33620 4349 33621
rect 12940 33620 12980 33748
rect 18115 33747 18173 33748
rect 21424 33705 21504 33724
rect 18691 33704 18749 33705
rect 15715 33664 15724 33704
rect 15764 33664 18412 33704
rect 18452 33664 18700 33704
rect 18740 33664 18749 33704
rect 18691 33663 18749 33664
rect 21379 33704 21504 33705
rect 21379 33664 21388 33704
rect 21428 33664 21504 33704
rect 21379 33663 21504 33664
rect 21424 33644 21504 33663
rect 16579 33620 16637 33621
rect 4272 33580 4300 33620
rect 4340 33580 4396 33620
rect 4436 33580 10732 33620
rect 10772 33580 10781 33620
rect 12835 33580 12844 33620
rect 12884 33580 12980 33620
rect 14467 33580 14476 33620
rect 14516 33580 14525 33620
rect 16579 33580 16588 33620
rect 16628 33580 19468 33620
rect 19508 33580 19517 33620
rect 4291 33579 4349 33580
rect 0 33536 80 33556
rect 1219 33536 1277 33537
rect 6211 33536 6269 33537
rect 14476 33536 14516 33580
rect 16579 33579 16637 33580
rect 17251 33536 17309 33537
rect 0 33496 1228 33536
rect 1268 33496 1277 33536
rect 4867 33496 4876 33536
rect 4916 33496 5932 33536
rect 5972 33496 5981 33536
rect 6211 33496 6220 33536
rect 6260 33496 6412 33536
rect 6452 33496 6461 33536
rect 10531 33496 10540 33536
rect 10580 33496 17260 33536
rect 17300 33496 17309 33536
rect 0 33476 80 33496
rect 1219 33495 1277 33496
rect 6211 33495 6269 33496
rect 17251 33495 17309 33496
rect 5827 33452 5885 33453
rect 6220 33452 6260 33495
rect 2659 33412 2668 33452
rect 2708 33412 4108 33452
rect 4148 33412 4157 33452
rect 4483 33412 4492 33452
rect 4532 33412 5452 33452
rect 5492 33412 5836 33452
rect 5876 33412 6260 33452
rect 14275 33412 14284 33452
rect 14324 33412 18220 33452
rect 18260 33412 18269 33452
rect 5827 33411 5885 33412
rect 13315 33368 13373 33369
rect 21424 33368 21504 33388
rect 5347 33328 5356 33368
rect 5396 33328 7180 33368
rect 7220 33328 7229 33368
rect 13315 33328 13324 33368
rect 13364 33328 13804 33368
rect 13844 33328 13853 33368
rect 18691 33328 18700 33368
rect 18740 33328 21504 33368
rect 13315 33327 13373 33328
rect 21424 33308 21504 33328
rect 16867 33284 16925 33285
rect 3679 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 4065 33284
rect 4387 33244 4396 33284
rect 4436 33244 4972 33284
rect 5012 33244 5021 33284
rect 12163 33244 12172 33284
rect 12212 33244 13420 33284
rect 13460 33244 14092 33284
rect 14132 33244 14572 33284
rect 14612 33244 14621 33284
rect 14947 33244 14956 33284
rect 14996 33244 16876 33284
rect 16916 33244 17260 33284
rect 17300 33244 17309 33284
rect 18799 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 19185 33284
rect 16867 33243 16925 33244
rect 21379 33200 21437 33201
rect 12643 33160 12652 33200
rect 12692 33160 21388 33200
rect 21428 33160 21437 33200
rect 21379 33159 21437 33160
rect 4675 33116 4733 33117
rect 4675 33076 4684 33116
rect 4724 33076 4876 33116
rect 4916 33076 4925 33116
rect 11971 33076 11980 33116
rect 12020 33076 13228 33116
rect 13268 33076 17972 33116
rect 19171 33076 19180 33116
rect 19220 33076 19852 33116
rect 19892 33076 19901 33116
rect 4675 33075 4733 33076
rect 17932 33033 17972 33076
rect 3235 33032 3293 33033
rect 15043 33032 15101 33033
rect 16579 33032 16637 33033
rect 17443 33032 17501 33033
rect 3235 32992 3244 33032
rect 3284 32992 3340 33032
rect 3380 32992 3389 33032
rect 7939 32992 7948 33032
rect 7988 32992 8332 33032
rect 8372 32992 8381 33032
rect 8428 32992 10924 33032
rect 10964 32992 10973 33032
rect 13228 32992 13420 33032
rect 13460 32992 13469 33032
rect 13603 32992 13612 33032
rect 13652 32992 15052 33032
rect 15092 32992 16588 33032
rect 16628 32992 16637 33032
rect 17347 32992 17356 33032
rect 17396 32992 17452 33032
rect 17492 32992 17501 33032
rect 3235 32991 3293 32992
rect 1603 32948 1661 32949
rect 1603 32908 1612 32948
rect 1652 32908 4148 32948
rect 4675 32908 4684 32948
rect 4724 32908 6796 32948
rect 6836 32908 8044 32948
rect 8084 32908 8093 32948
rect 1603 32907 1661 32908
rect 0 32864 80 32884
rect 2563 32864 2621 32865
rect 4108 32864 4148 32908
rect 8428 32864 8468 32992
rect 13228 32948 13268 32992
rect 15043 32991 15101 32992
rect 16579 32991 16637 32992
rect 17443 32991 17501 32992
rect 17923 33032 17981 33033
rect 21424 33032 21504 33052
rect 17923 32992 17932 33032
rect 17972 32992 19756 33032
rect 19796 32992 19805 33032
rect 19939 32992 19948 33032
rect 19988 32992 21504 33032
rect 17923 32991 17981 32992
rect 21424 32972 21504 32992
rect 10627 32908 10636 32948
rect 10676 32908 11212 32948
rect 11252 32908 11261 32948
rect 13219 32908 13228 32948
rect 13268 32908 13277 32948
rect 13507 32908 13516 32948
rect 13556 32908 18604 32948
rect 18644 32908 18653 32948
rect 14083 32864 14141 32865
rect 0 32824 2572 32864
rect 2612 32824 2621 32864
rect 2851 32824 2860 32864
rect 2900 32824 3820 32864
rect 3860 32824 3869 32864
rect 4099 32824 4108 32864
rect 4148 32824 8468 32864
rect 10147 32824 10156 32864
rect 10196 32824 10732 32864
rect 10772 32824 10781 32864
rect 10915 32824 10924 32864
rect 10964 32824 14092 32864
rect 14132 32824 18028 32864
rect 18068 32824 18796 32864
rect 18836 32824 19372 32864
rect 19412 32824 19421 32864
rect 0 32804 80 32824
rect 2563 32823 2621 32824
rect 14083 32823 14141 32824
rect 1123 32780 1181 32781
rect 17443 32780 17501 32781
rect 1123 32740 1132 32780
rect 1172 32740 1228 32780
rect 1268 32740 2092 32780
rect 2132 32740 2141 32780
rect 7171 32740 7180 32780
rect 7220 32740 7468 32780
rect 7508 32740 7517 32780
rect 7651 32740 7660 32780
rect 7700 32740 7948 32780
rect 7988 32740 7997 32780
rect 8515 32740 8524 32780
rect 8564 32740 11020 32780
rect 11060 32740 11308 32780
rect 11348 32740 11357 32780
rect 11779 32740 11788 32780
rect 11828 32740 17452 32780
rect 17492 32740 17501 32780
rect 18403 32740 18412 32780
rect 18452 32740 19852 32780
rect 19892 32740 19901 32780
rect 1123 32739 1181 32740
rect 17443 32739 17501 32740
rect 3235 32696 3293 32697
rect 13411 32696 13469 32697
rect 17635 32696 17693 32697
rect 3139 32656 3148 32696
rect 3188 32656 3244 32696
rect 3284 32656 3293 32696
rect 13326 32656 13420 32696
rect 13460 32656 13469 32696
rect 16771 32656 16780 32696
rect 16820 32656 17548 32696
rect 17588 32656 17644 32696
rect 17684 32656 17693 32696
rect 3235 32655 3293 32656
rect 13411 32655 13469 32656
rect 17635 32655 17693 32656
rect 18211 32696 18269 32697
rect 21424 32696 21504 32716
rect 18211 32656 18220 32696
rect 18260 32656 18316 32696
rect 18356 32656 18365 32696
rect 20419 32656 20428 32696
rect 20468 32656 21004 32696
rect 21044 32656 21053 32696
rect 18211 32655 18269 32656
rect 21388 32636 21504 32696
rect 2851 32612 2909 32613
rect 21388 32612 21428 32636
rect 2851 32572 2860 32612
rect 2900 32572 5644 32612
rect 5684 32572 6028 32612
rect 6068 32572 8840 32612
rect 19651 32572 19660 32612
rect 19700 32572 21428 32612
rect 2851 32571 2909 32572
rect 8800 32528 8840 32572
rect 3523 32488 3532 32528
rect 3572 32488 4780 32528
rect 4820 32488 4829 32528
rect 4919 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 5305 32528
rect 8800 32488 12940 32528
rect 12980 32488 13516 32528
rect 13556 32488 13565 32528
rect 13612 32488 18988 32528
rect 19028 32488 19037 32528
rect 20039 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20425 32528
rect 13612 32444 13652 32488
rect 1507 32404 1516 32444
rect 1556 32404 8428 32444
rect 8468 32404 12652 32444
rect 12692 32404 13652 32444
rect 13699 32404 13708 32444
rect 13748 32404 16780 32444
rect 16820 32404 16829 32444
rect 4099 32360 4157 32361
rect 13411 32360 13469 32361
rect 20707 32360 20765 32361
rect 21424 32360 21504 32380
rect 1315 32320 1324 32360
rect 1364 32320 4108 32360
rect 4148 32320 4157 32360
rect 7075 32320 7084 32360
rect 7124 32320 8044 32360
rect 8084 32320 8093 32360
rect 9859 32320 9868 32360
rect 9908 32320 10060 32360
rect 10100 32320 10109 32360
rect 13219 32320 13228 32360
rect 13268 32320 13420 32360
rect 13460 32320 13469 32360
rect 15715 32320 15724 32360
rect 15764 32320 16108 32360
rect 16148 32320 16157 32360
rect 20707 32320 20716 32360
rect 20756 32320 21504 32360
rect 4099 32319 4157 32320
rect 13411 32319 13469 32320
rect 20707 32319 20765 32320
rect 21424 32300 21504 32320
rect 16963 32276 17021 32277
rect 1123 32236 1132 32276
rect 1172 32236 16972 32276
rect 17012 32236 17021 32276
rect 16963 32235 17021 32236
rect 18691 32276 18749 32277
rect 18691 32236 18700 32276
rect 18740 32236 20044 32276
rect 20084 32236 20093 32276
rect 18691 32235 18749 32236
rect 0 32192 80 32212
rect 2851 32192 2909 32193
rect 18211 32192 18269 32193
rect 0 32152 2188 32192
rect 2228 32152 2237 32192
rect 2766 32152 2860 32192
rect 2900 32152 2909 32192
rect 3523 32152 3532 32192
rect 3572 32152 4492 32192
rect 4532 32152 4541 32192
rect 6115 32152 6124 32192
rect 6164 32152 7756 32192
rect 7796 32152 7805 32192
rect 10060 32152 11404 32192
rect 11444 32152 11453 32192
rect 13315 32152 13324 32192
rect 13364 32152 13996 32192
rect 14036 32152 14045 32192
rect 14275 32152 14284 32192
rect 14324 32152 15148 32192
rect 15188 32152 16300 32192
rect 16340 32152 16349 32192
rect 16483 32152 16492 32192
rect 16532 32152 17356 32192
rect 17396 32152 17405 32192
rect 18211 32152 18220 32192
rect 18260 32152 18604 32192
rect 18644 32152 18653 32192
rect 0 32132 80 32152
rect 2851 32151 2909 32152
rect 2947 32108 3005 32109
rect 10060 32108 10100 32152
rect 1891 32068 1900 32108
rect 1940 32068 2476 32108
rect 2516 32068 2525 32108
rect 2755 32068 2764 32108
rect 2804 32068 2956 32108
rect 2996 32068 3005 32108
rect 3235 32068 3244 32108
rect 3284 32068 4588 32108
rect 4628 32068 4637 32108
rect 6979 32068 6988 32108
rect 7028 32068 8812 32108
rect 8852 32068 9676 32108
rect 9716 32068 10100 32108
rect 13996 32108 14036 32152
rect 18211 32151 18269 32152
rect 13996 32068 14380 32108
rect 14420 32068 14429 32108
rect 2947 32067 3005 32068
rect 19843 32024 19901 32025
rect 21424 32024 21504 32044
rect 19843 31984 19852 32024
rect 19892 31984 21504 32024
rect 19843 31983 19901 31984
rect 21424 31964 21504 31984
rect 4771 31940 4829 31941
rect 2467 31900 2476 31940
rect 2516 31900 4780 31940
rect 4820 31900 4829 31940
rect 4771 31899 4829 31900
rect 3679 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 4065 31772
rect 18799 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 19185 31772
rect 4675 31688 4733 31689
rect 21424 31688 21504 31708
rect 4590 31648 4684 31688
rect 4724 31648 4733 31688
rect 17347 31648 17356 31688
rect 17396 31648 17405 31688
rect 20515 31648 20524 31688
rect 20564 31648 21504 31688
rect 4675 31647 4733 31648
rect 17356 31604 17396 31648
rect 21424 31628 21504 31648
rect 4579 31564 4588 31604
rect 4628 31564 6988 31604
rect 7028 31564 7037 31604
rect 12643 31564 12652 31604
rect 12692 31564 13420 31604
rect 13460 31564 13469 31604
rect 17356 31564 19084 31604
rect 19124 31564 19133 31604
rect 0 31520 80 31540
rect 13123 31520 13181 31521
rect 0 31480 652 31520
rect 692 31480 701 31520
rect 5443 31480 5452 31520
rect 5492 31480 5932 31520
rect 5972 31480 5981 31520
rect 6691 31480 6700 31520
rect 6740 31480 7276 31520
rect 7316 31480 7325 31520
rect 8803 31480 8812 31520
rect 8852 31480 11116 31520
rect 11156 31480 11165 31520
rect 13038 31480 13132 31520
rect 13172 31480 13324 31520
rect 13364 31480 13373 31520
rect 14755 31480 14764 31520
rect 14804 31480 15244 31520
rect 15284 31480 15293 31520
rect 16195 31480 16204 31520
rect 16244 31480 19372 31520
rect 19412 31480 19421 31520
rect 0 31460 80 31480
rect 13123 31479 13181 31480
rect 18115 31436 18173 31437
rect 2500 31396 9004 31436
rect 9044 31396 9053 31436
rect 9187 31396 9196 31436
rect 9236 31396 17164 31436
rect 17204 31396 17213 31436
rect 17731 31396 17740 31436
rect 17780 31396 18124 31436
rect 18164 31396 18173 31436
rect 2083 31312 2092 31352
rect 2132 31312 2380 31352
rect 2420 31312 2429 31352
rect 0 30848 80 30868
rect 0 30808 1132 30848
rect 1172 30808 1181 30848
rect 0 30788 80 30808
rect 2500 30764 2540 31396
rect 18115 31395 18173 31396
rect 5347 31352 5405 31353
rect 13987 31352 14045 31353
rect 14755 31352 14813 31353
rect 21424 31352 21504 31372
rect 5059 31312 5068 31352
rect 5108 31312 5356 31352
rect 5396 31312 5405 31352
rect 6883 31312 6892 31352
rect 6932 31312 8044 31352
rect 8084 31312 8524 31352
rect 8564 31312 10156 31352
rect 10196 31312 10205 31352
rect 13987 31312 13996 31352
rect 14036 31312 14764 31352
rect 14804 31312 15532 31352
rect 15572 31312 15581 31352
rect 17443 31312 17452 31352
rect 17492 31312 21504 31352
rect 5347 31311 5405 31312
rect 10156 31268 10196 31312
rect 13987 31311 14045 31312
rect 14755 31311 14813 31312
rect 21424 31292 21504 31312
rect 5155 31228 5164 31268
rect 5204 31228 8140 31268
rect 8180 31228 8189 31268
rect 10156 31228 14572 31268
rect 14612 31228 14621 31268
rect 15331 31228 15340 31268
rect 15380 31228 17836 31268
rect 17876 31228 18124 31268
rect 18164 31228 18173 31268
rect 5635 31184 5693 31185
rect 5550 31144 5644 31184
rect 5684 31144 5693 31184
rect 7075 31144 7084 31184
rect 7124 31144 7660 31184
rect 7700 31144 7709 31184
rect 8707 31144 8716 31184
rect 8756 31144 9196 31184
rect 9236 31144 9245 31184
rect 12355 31144 12364 31184
rect 12404 31144 16780 31184
rect 16820 31144 16829 31184
rect 19555 31144 19564 31184
rect 19604 31144 21332 31184
rect 5635 31143 5693 31144
rect 2851 31100 2909 31101
rect 2766 31060 2860 31100
rect 2900 31060 16340 31100
rect 16387 31060 16396 31100
rect 16436 31060 16684 31100
rect 16724 31060 16733 31100
rect 2851 31059 2909 31060
rect 5539 31016 5597 31017
rect 16300 31016 16340 31060
rect 17059 31016 17117 31017
rect 21292 31016 21332 31144
rect 21424 31016 21504 31036
rect 4919 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 5305 31016
rect 5443 30976 5452 31016
rect 5492 30976 5548 31016
rect 5588 30976 5597 31016
rect 8131 30976 8140 31016
rect 8180 30976 8620 31016
rect 8660 30976 11212 31016
rect 11252 30976 11261 31016
rect 16300 30976 17068 31016
rect 17108 30976 17356 31016
rect 17396 30976 17405 31016
rect 20039 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20425 31016
rect 21292 30976 21504 31016
rect 5539 30975 5597 30976
rect 17059 30975 17117 30976
rect 21424 30956 21504 30976
rect 13795 30932 13853 30933
rect 4483 30892 4492 30932
rect 4532 30892 13804 30932
rect 13844 30892 13853 30932
rect 13795 30891 13853 30892
rect 14476 30892 19756 30932
rect 19796 30892 19805 30932
rect 12259 30848 12317 30849
rect 14476 30848 14516 30892
rect 7843 30808 7852 30848
rect 7892 30808 12268 30848
rect 12308 30808 14516 30848
rect 14755 30808 14764 30848
rect 14804 30808 17260 30848
rect 17300 30808 17309 30848
rect 12259 30807 12317 30808
rect 1795 30724 1804 30764
rect 1844 30724 2540 30764
rect 3427 30724 3436 30764
rect 3476 30724 7892 30764
rect 2467 30680 2525 30681
rect 3523 30680 3581 30681
rect 5827 30680 5885 30681
rect 7852 30680 7892 30724
rect 18019 30680 18077 30681
rect 21424 30680 21504 30700
rect 2382 30640 2476 30680
rect 2516 30640 2525 30680
rect 3331 30640 3340 30680
rect 3380 30640 3532 30680
rect 3572 30640 3581 30680
rect 4387 30640 4396 30680
rect 4436 30640 4780 30680
rect 4820 30640 5068 30680
rect 5108 30640 5117 30680
rect 5827 30640 5836 30680
rect 5876 30640 7276 30680
rect 7316 30640 7325 30680
rect 7843 30640 7852 30680
rect 7892 30640 10828 30680
rect 10868 30640 11116 30680
rect 11156 30640 11165 30680
rect 14563 30640 14572 30680
rect 14612 30640 16204 30680
rect 16244 30640 16876 30680
rect 16916 30640 16925 30680
rect 17827 30640 17836 30680
rect 17876 30640 18028 30680
rect 18068 30640 18077 30680
rect 20611 30640 20620 30680
rect 20660 30640 21504 30680
rect 2467 30639 2525 30640
rect 3523 30639 3581 30640
rect 5827 30639 5885 30640
rect 18019 30639 18077 30640
rect 21424 30620 21504 30640
rect 5539 30596 5597 30597
rect 9667 30596 9725 30597
rect 5454 30556 5548 30596
rect 5588 30556 5597 30596
rect 7363 30556 7372 30596
rect 7412 30556 9676 30596
rect 9716 30556 9725 30596
rect 5539 30555 5597 30556
rect 9667 30555 9725 30556
rect 12835 30596 12893 30597
rect 12835 30556 12844 30596
rect 12884 30556 15532 30596
rect 15572 30556 19372 30596
rect 19412 30556 19421 30596
rect 12835 30555 12893 30556
rect 7267 30512 7325 30513
rect 5347 30472 5356 30512
rect 5396 30472 5644 30512
rect 5684 30472 7276 30512
rect 7316 30472 7325 30512
rect 8323 30472 8332 30512
rect 8372 30472 11692 30512
rect 11732 30472 11741 30512
rect 16195 30472 16204 30512
rect 16244 30472 17932 30512
rect 17972 30472 17981 30512
rect 7267 30471 7325 30472
rect 5155 30388 5164 30428
rect 5204 30388 5740 30428
rect 5780 30388 6412 30428
rect 6452 30388 6461 30428
rect 17827 30388 17836 30428
rect 17876 30388 18124 30428
rect 18164 30388 18173 30428
rect 18979 30388 18988 30428
rect 19028 30388 19468 30428
rect 19508 30388 19517 30428
rect 20611 30344 20669 30345
rect 21424 30344 21504 30364
rect 6691 30304 6700 30344
rect 6740 30304 8084 30344
rect 15427 30304 15436 30344
rect 15476 30304 18740 30344
rect 8044 30260 8084 30304
rect 11011 30260 11069 30261
rect 18700 30260 18740 30304
rect 20611 30304 20620 30344
rect 20660 30304 21504 30344
rect 20611 30303 20669 30304
rect 21424 30284 21504 30304
rect 3679 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 4065 30260
rect 4771 30220 4780 30260
rect 4820 30220 6028 30260
rect 6068 30220 6988 30260
rect 7028 30220 7037 30260
rect 8035 30220 8044 30260
rect 8084 30220 8564 30260
rect 8899 30220 8908 30260
rect 8948 30220 9484 30260
rect 9524 30220 11020 30260
rect 11060 30220 11069 30260
rect 15043 30220 15052 30260
rect 15092 30220 16492 30260
rect 16532 30220 16541 30260
rect 17059 30220 17068 30260
rect 17108 30220 17740 30260
rect 17780 30220 17789 30260
rect 18691 30220 18700 30260
rect 18740 30220 18749 30260
rect 18799 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 19185 30260
rect 0 30176 80 30196
rect 5443 30176 5501 30177
rect 8524 30176 8564 30220
rect 11011 30219 11069 30220
rect 0 30136 5452 30176
rect 5492 30136 5501 30176
rect 6211 30136 6220 30176
rect 6260 30136 7180 30176
rect 7220 30136 7229 30176
rect 8515 30136 8524 30176
rect 8564 30136 8573 30176
rect 14851 30136 14860 30176
rect 14900 30136 19756 30176
rect 19796 30136 19805 30176
rect 0 30116 80 30136
rect 5443 30135 5501 30136
rect 7651 30092 7709 30093
rect 20707 30092 20765 30093
rect 1987 30052 1996 30092
rect 2036 30052 2668 30092
rect 2708 30052 2717 30092
rect 6403 30052 6412 30092
rect 6452 30052 7084 30092
rect 7124 30052 7133 30092
rect 7651 30052 7660 30092
rect 7700 30052 8620 30092
rect 8660 30052 8669 30092
rect 11971 30052 11980 30092
rect 12020 30052 17164 30092
rect 17204 30052 17213 30092
rect 17539 30052 17548 30092
rect 17588 30052 18316 30092
rect 18356 30052 18365 30092
rect 19843 30052 19852 30092
rect 19892 30052 20716 30092
rect 20756 30052 20765 30092
rect 7651 30051 7709 30052
rect 20707 30051 20765 30052
rect 21424 30008 21504 30028
rect 3139 29968 3148 30008
rect 3188 29968 4108 30008
rect 4148 29968 8908 30008
rect 8948 29968 8957 30008
rect 15811 29968 15820 30008
rect 15860 29968 16300 30008
rect 16340 29968 16349 30008
rect 20707 29968 20716 30008
rect 20756 29968 21504 30008
rect 21424 29948 21504 29968
rect 5635 29924 5693 29925
rect 17443 29924 17501 29925
rect 1987 29884 1996 29924
rect 2036 29884 5452 29924
rect 5492 29884 5501 29924
rect 5635 29884 5644 29924
rect 5684 29884 10540 29924
rect 10580 29884 11020 29924
rect 11060 29884 11069 29924
rect 14851 29884 14860 29924
rect 14900 29884 16588 29924
rect 16628 29884 16820 29924
rect 5635 29883 5693 29884
rect 9667 29840 9725 29841
rect 2179 29800 2188 29840
rect 2228 29800 3148 29840
rect 3188 29800 3197 29840
rect 3811 29800 3820 29840
rect 3860 29800 3869 29840
rect 4579 29800 4588 29840
rect 4628 29800 5356 29840
rect 5396 29800 5405 29840
rect 5539 29800 5548 29840
rect 5588 29800 5836 29840
rect 5876 29800 6604 29840
rect 6644 29800 6653 29840
rect 7843 29800 7852 29840
rect 7892 29800 8716 29840
rect 8756 29800 8765 29840
rect 9091 29800 9100 29840
rect 9140 29800 9676 29840
rect 9716 29800 9725 29840
rect 10339 29800 10348 29840
rect 10388 29800 11596 29840
rect 11636 29800 11645 29840
rect 12163 29800 12172 29840
rect 12212 29800 13708 29840
rect 13748 29800 13757 29840
rect 13987 29800 13996 29840
rect 14036 29800 15916 29840
rect 15956 29800 15965 29840
rect 3820 29756 3860 29800
rect 9667 29799 9725 29800
rect 13603 29756 13661 29757
rect 16780 29756 16820 29884
rect 17443 29884 17452 29924
rect 17492 29884 20044 29924
rect 20084 29884 20093 29924
rect 17443 29883 17501 29884
rect 17059 29840 17117 29841
rect 17059 29800 17068 29840
rect 17108 29800 17740 29840
rect 17780 29800 17789 29840
rect 19363 29800 19372 29840
rect 19412 29800 19852 29840
rect 19892 29800 19901 29840
rect 17059 29799 17117 29800
rect 3820 29716 8236 29756
rect 8276 29716 8285 29756
rect 13603 29716 13612 29756
rect 13652 29716 13900 29756
rect 13940 29716 13949 29756
rect 14755 29716 14764 29756
rect 14804 29716 16148 29756
rect 16771 29716 16780 29756
rect 16820 29716 16829 29756
rect 13603 29715 13661 29716
rect 6019 29672 6077 29673
rect 14371 29672 14429 29673
rect 1411 29632 1420 29672
rect 1460 29632 3628 29672
rect 3668 29632 3677 29672
rect 4099 29632 4108 29672
rect 4148 29632 4684 29672
rect 4724 29632 4733 29672
rect 6019 29632 6028 29672
rect 6068 29632 6220 29672
rect 6260 29632 6269 29672
rect 11320 29632 14380 29672
rect 14420 29632 14429 29672
rect 15331 29632 15340 29672
rect 15380 29632 15724 29672
rect 15764 29632 15773 29672
rect 6019 29631 6077 29632
rect 4003 29548 4012 29588
rect 4052 29548 4396 29588
rect 4436 29548 4445 29588
rect 0 29504 80 29524
rect 2275 29504 2333 29505
rect 6211 29504 6269 29505
rect 0 29464 2284 29504
rect 2324 29464 2333 29504
rect 3811 29464 3820 29504
rect 3860 29464 4588 29504
rect 4628 29464 4637 29504
rect 4919 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 5305 29504
rect 5347 29464 5356 29504
rect 5396 29464 6220 29504
rect 6260 29464 10924 29504
rect 10964 29464 10973 29504
rect 0 29444 80 29464
rect 2275 29463 2333 29464
rect 6211 29463 6269 29464
rect 2659 29380 2668 29420
rect 2708 29380 5204 29420
rect 5923 29380 5932 29420
rect 5972 29380 7276 29420
rect 7316 29380 7325 29420
rect 2275 29336 2333 29337
rect 5164 29336 5204 29380
rect 10819 29336 10877 29337
rect 2190 29296 2284 29336
rect 2324 29296 2333 29336
rect 3715 29296 3724 29336
rect 3764 29296 4972 29336
rect 5012 29296 5021 29336
rect 5155 29296 5164 29336
rect 5204 29296 5213 29336
rect 8227 29296 8236 29336
rect 8276 29296 10828 29336
rect 10868 29296 10877 29336
rect 2275 29295 2333 29296
rect 10819 29295 10877 29296
rect 11320 29252 11360 29632
rect 14371 29631 14429 29632
rect 16108 29588 16148 29716
rect 16963 29672 17021 29673
rect 17068 29672 17108 29799
rect 17251 29756 17309 29757
rect 17251 29716 17260 29756
rect 17300 29716 19660 29756
rect 19700 29716 19709 29756
rect 17251 29715 17309 29716
rect 19363 29672 19421 29673
rect 21424 29672 21504 29692
rect 16579 29632 16588 29672
rect 16628 29632 16972 29672
rect 17012 29632 17108 29672
rect 17347 29632 17356 29672
rect 17396 29632 19372 29672
rect 19412 29632 19421 29672
rect 19939 29632 19948 29672
rect 19988 29632 21504 29672
rect 16963 29631 17021 29632
rect 19363 29631 19421 29632
rect 21424 29612 21504 29632
rect 17635 29588 17693 29589
rect 18307 29588 18365 29589
rect 12355 29548 12364 29588
rect 12404 29548 15244 29588
rect 15284 29548 15293 29588
rect 16108 29548 17644 29588
rect 17684 29548 18316 29588
rect 18356 29548 18365 29588
rect 17635 29547 17693 29548
rect 18307 29547 18365 29548
rect 15427 29464 15436 29504
rect 15476 29464 15820 29504
rect 15860 29464 15869 29504
rect 18115 29464 18124 29504
rect 18164 29464 18508 29504
rect 18548 29464 18557 29504
rect 20039 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20425 29504
rect 15043 29380 15052 29420
rect 15092 29380 17548 29420
rect 17588 29380 17597 29420
rect 17932 29380 18220 29420
rect 18260 29380 18269 29420
rect 14851 29336 14909 29337
rect 17932 29336 17972 29380
rect 21424 29336 21504 29356
rect 14083 29296 14092 29336
rect 14132 29296 14476 29336
rect 14516 29296 14525 29336
rect 14851 29296 14860 29336
rect 14900 29296 14956 29336
rect 14996 29296 15005 29336
rect 16291 29296 16300 29336
rect 16340 29296 17972 29336
rect 18019 29296 18028 29336
rect 18068 29296 18412 29336
rect 18452 29296 18461 29336
rect 19267 29296 19276 29336
rect 19316 29296 19852 29336
rect 19892 29296 19901 29336
rect 21379 29296 21388 29336
rect 21428 29296 21504 29336
rect 14851 29295 14909 29296
rect 21424 29276 21504 29296
rect 19267 29252 19325 29253
rect 259 29212 268 29252
rect 308 29212 11360 29252
rect 11587 29212 11596 29252
rect 11636 29212 12268 29252
rect 12308 29212 13996 29252
rect 14036 29212 15148 29252
rect 15188 29212 15197 29252
rect 17059 29212 17068 29252
rect 17108 29212 19276 29252
rect 19316 29212 19325 29252
rect 19267 29211 19325 29212
rect 19459 29252 19517 29253
rect 19459 29212 19468 29252
rect 19508 29212 20180 29252
rect 19459 29211 19517 29212
rect 8227 29168 8285 29169
rect 2179 29128 2188 29168
rect 2228 29128 3380 29168
rect 3907 29128 3916 29168
rect 3956 29128 5164 29168
rect 5204 29128 5213 29168
rect 6307 29128 6316 29168
rect 6356 29128 6700 29168
rect 6740 29128 6749 29168
rect 6979 29128 6988 29168
rect 7028 29128 7180 29168
rect 7220 29128 7229 29168
rect 7459 29128 7468 29168
rect 7508 29128 7660 29168
rect 7700 29128 7709 29168
rect 8142 29128 8236 29168
rect 8276 29128 8285 29168
rect 15907 29128 15916 29168
rect 15956 29128 16492 29168
rect 16532 29128 16541 29168
rect 17923 29128 17932 29168
rect 17972 29128 18508 29168
rect 18548 29128 19700 29168
rect 19747 29128 19756 29168
rect 19796 29128 20044 29168
rect 20084 29128 20093 29168
rect 3340 29084 3380 29128
rect 2275 29044 2284 29084
rect 2324 29044 3052 29084
rect 3092 29044 3101 29084
rect 3331 29044 3340 29084
rect 3380 29044 4485 29084
rect 4525 29044 4534 29084
rect 4588 29000 4628 29128
rect 8227 29127 8285 29128
rect 19660 29084 19700 29128
rect 5059 29044 5068 29084
rect 5108 29044 5644 29084
rect 5684 29044 5693 29084
rect 13795 29044 13804 29084
rect 13844 29044 15092 29084
rect 15331 29044 15340 29084
rect 15380 29044 16972 29084
rect 17012 29044 17021 29084
rect 17068 29044 17836 29084
rect 17876 29044 17885 29084
rect 19651 29044 19660 29084
rect 19700 29044 19709 29084
rect 15052 29000 15092 29044
rect 4579 28960 4588 29000
rect 4628 28960 4637 29000
rect 15012 28960 15052 29000
rect 15092 28960 15101 29000
rect 10819 28916 10877 28917
rect 17068 28916 17108 29044
rect 20140 29000 20180 29212
rect 21424 29000 21504 29020
rect 19555 28960 19564 29000
rect 19604 28960 19613 29000
rect 20140 28960 21504 29000
rect 19564 28916 19604 28960
rect 21424 28940 21504 28960
rect 2947 28876 2956 28916
rect 2996 28876 3724 28916
rect 3764 28876 3773 28916
rect 10723 28876 10732 28916
rect 10772 28876 10828 28916
rect 10868 28876 10877 28916
rect 17059 28876 17068 28916
rect 17108 28876 17117 28916
rect 17923 28876 17932 28916
rect 17972 28876 18316 28916
rect 18356 28876 18365 28916
rect 19564 28876 19660 28916
rect 19700 28876 19709 28916
rect 10819 28875 10877 28876
rect 0 28832 80 28852
rect 547 28832 605 28833
rect 2467 28832 2525 28833
rect 0 28792 556 28832
rect 596 28792 605 28832
rect 2371 28792 2380 28832
rect 2420 28792 2476 28832
rect 2516 28792 2525 28832
rect 9379 28792 9388 28832
rect 9428 28792 19564 28832
rect 19604 28792 19613 28832
rect 0 28772 80 28792
rect 547 28791 605 28792
rect 2467 28791 2525 28792
rect 3679 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 4065 28748
rect 11491 28708 11500 28748
rect 11540 28708 11980 28748
rect 12020 28708 12029 28748
rect 18799 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 19185 28748
rect 19555 28664 19613 28665
rect 21424 28664 21504 28684
rect 4291 28624 4300 28664
rect 4340 28624 4492 28664
rect 4532 28624 4541 28664
rect 11875 28624 11884 28664
rect 11924 28624 12556 28664
rect 12596 28624 12605 28664
rect 13027 28624 13036 28664
rect 13076 28624 13228 28664
rect 13268 28624 15628 28664
rect 15668 28624 17356 28664
rect 17396 28624 17405 28664
rect 18307 28624 18316 28664
rect 18356 28624 18700 28664
rect 18740 28624 18749 28664
rect 19555 28624 19564 28664
rect 19604 28624 21504 28664
rect 19555 28623 19613 28624
rect 21424 28604 21504 28624
rect 20611 28580 20669 28581
rect 8899 28540 8908 28580
rect 8948 28540 11360 28580
rect 12643 28540 12652 28580
rect 12692 28540 13420 28580
rect 13460 28540 13469 28580
rect 18595 28540 18604 28580
rect 18644 28540 18988 28580
rect 19028 28540 19037 28580
rect 19747 28540 19756 28580
rect 19796 28540 20620 28580
rect 20660 28540 20669 28580
rect 11320 28496 11360 28540
rect 20611 28539 20669 28540
rect 3139 28456 3148 28496
rect 3188 28456 4108 28496
rect 4148 28456 4300 28496
rect 4340 28456 4349 28496
rect 6883 28456 6892 28496
rect 6932 28456 7564 28496
rect 7604 28456 7613 28496
rect 9859 28456 9868 28496
rect 9908 28456 10252 28496
rect 10292 28456 10301 28496
rect 11320 28456 19852 28496
rect 19892 28456 19901 28496
rect 10723 28412 10781 28413
rect 3523 28372 3532 28412
rect 3572 28372 10732 28412
rect 10772 28372 10781 28412
rect 11280 28372 11308 28412
rect 11348 28372 11444 28412
rect 17251 28372 17260 28412
rect 17300 28372 19948 28412
rect 19988 28372 19997 28412
rect 10723 28371 10781 28372
rect 3235 28328 3293 28329
rect 4483 28328 4541 28329
rect 11404 28328 11444 28372
rect 13987 28328 14045 28329
rect 16291 28328 16349 28329
rect 3235 28288 3244 28328
rect 3284 28288 3628 28328
rect 3668 28288 3677 28328
rect 4099 28288 4108 28328
rect 4148 28288 4492 28328
rect 4532 28288 4541 28328
rect 6979 28288 6988 28328
rect 7028 28288 7276 28328
rect 7316 28288 7325 28328
rect 10243 28288 10252 28328
rect 10292 28288 10444 28328
rect 10484 28288 10493 28328
rect 11395 28288 11404 28328
rect 11444 28288 11453 28328
rect 12163 28288 12172 28328
rect 12212 28288 12221 28328
rect 12931 28288 12940 28328
rect 12980 28288 13804 28328
rect 13844 28288 13853 28328
rect 13987 28288 13996 28328
rect 14036 28288 14130 28328
rect 15235 28288 15244 28328
rect 15284 28288 16108 28328
rect 16148 28288 16300 28328
rect 16340 28288 16349 28328
rect 3235 28287 3293 28288
rect 4483 28287 4541 28288
rect 12172 28244 12212 28288
rect 13987 28287 14045 28288
rect 16291 28287 16349 28288
rect 17251 28328 17309 28329
rect 21424 28328 21504 28348
rect 17251 28288 17260 28328
rect 17300 28288 17548 28328
rect 17588 28288 17597 28328
rect 19651 28288 19660 28328
rect 19700 28288 21504 28328
rect 17251 28287 17309 28288
rect 21424 28268 21504 28288
rect 19747 28244 19805 28245
rect 20707 28244 20765 28245
rect 5731 28204 5740 28244
rect 5780 28204 7180 28244
rect 7220 28204 7229 28244
rect 12172 28204 16588 28244
rect 16628 28204 16637 28244
rect 19747 28204 19756 28244
rect 19796 28204 20716 28244
rect 20756 28204 20765 28244
rect 19747 28203 19805 28204
rect 20707 28203 20765 28204
rect 0 28160 80 28180
rect 0 28120 1228 28160
rect 1268 28120 1277 28160
rect 11875 28120 11884 28160
rect 11924 28120 12364 28160
rect 12404 28120 16108 28160
rect 16148 28120 16157 28160
rect 16867 28120 16876 28160
rect 16916 28120 17356 28160
rect 17396 28120 17405 28160
rect 0 28100 80 28120
rect 14371 28036 14380 28076
rect 14420 28036 19084 28076
rect 19124 28036 19133 28076
rect 21424 27992 21504 28012
rect 2851 27952 2860 27992
rect 2900 27952 3244 27992
rect 3284 27952 3293 27992
rect 4919 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 5305 27992
rect 16675 27952 16684 27992
rect 16724 27952 17396 27992
rect 20039 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20425 27992
rect 20524 27952 21504 27992
rect 1507 27868 1516 27908
rect 1556 27868 1996 27908
rect 2036 27868 2045 27908
rect 14467 27868 14476 27908
rect 14516 27868 15436 27908
rect 15476 27868 16724 27908
rect 6019 27824 6077 27825
rect 3139 27784 3148 27824
rect 3188 27784 4588 27824
rect 4628 27784 4637 27824
rect 5731 27784 5740 27824
rect 5780 27784 6028 27824
rect 6068 27784 6077 27824
rect 6019 27783 6077 27784
rect 15331 27824 15389 27825
rect 16684 27824 16724 27868
rect 15331 27784 15340 27824
rect 15380 27784 15820 27824
rect 15860 27784 15869 27824
rect 16675 27784 16684 27824
rect 16724 27784 16733 27824
rect 15331 27783 15389 27784
rect 3523 27740 3581 27741
rect 6979 27740 7037 27741
rect 3523 27700 3532 27740
rect 3572 27700 3628 27740
rect 3668 27700 3677 27740
rect 6499 27700 6508 27740
rect 6548 27700 6988 27740
rect 7028 27700 7037 27740
rect 17356 27740 17396 27952
rect 20524 27908 20564 27952
rect 21424 27932 21504 27952
rect 19651 27868 19660 27908
rect 19700 27868 20564 27908
rect 20035 27784 20044 27824
rect 20084 27784 20180 27824
rect 20140 27740 20180 27784
rect 17356 27700 18836 27740
rect 20140 27700 20716 27740
rect 20756 27700 20765 27740
rect 3523 27699 3581 27700
rect 6979 27699 7037 27700
rect 1315 27656 1373 27657
rect 6595 27656 6653 27657
rect 7075 27656 7133 27657
rect 12259 27656 12317 27657
rect 18307 27656 18365 27657
rect 18796 27656 18836 27700
rect 21424 27656 21504 27676
rect 1219 27616 1228 27656
rect 1268 27616 1324 27656
rect 1364 27616 1373 27656
rect 2947 27616 2956 27656
rect 2996 27616 3188 27656
rect 3523 27616 3532 27656
rect 3572 27616 4108 27656
rect 4148 27616 4157 27656
rect 6595 27616 6604 27656
rect 6644 27616 6796 27656
rect 6836 27616 7084 27656
rect 7124 27616 7133 27656
rect 7267 27616 7276 27656
rect 7316 27616 8044 27656
rect 8084 27616 8093 27656
rect 12067 27616 12076 27656
rect 12116 27616 12268 27656
rect 12308 27616 12317 27656
rect 13987 27616 13996 27656
rect 14036 27616 15532 27656
rect 15572 27616 15581 27656
rect 18307 27616 18316 27656
rect 18356 27616 18700 27656
rect 18740 27616 18749 27656
rect 18796 27616 21504 27656
rect 1315 27615 1373 27616
rect 3148 27572 3188 27616
rect 6595 27615 6653 27616
rect 7075 27615 7133 27616
rect 12259 27615 12317 27616
rect 18307 27615 18365 27616
rect 4099 27572 4157 27573
rect 3139 27532 3148 27572
rect 3188 27532 3197 27572
rect 4099 27532 4108 27572
rect 4148 27532 8468 27572
rect 12163 27532 12172 27572
rect 12212 27532 12556 27572
rect 12596 27532 13324 27572
rect 13364 27532 15244 27572
rect 15284 27532 15293 27572
rect 17059 27532 17068 27572
rect 17108 27532 18220 27572
rect 18260 27532 18269 27572
rect 4099 27531 4157 27532
rect 0 27488 80 27508
rect 8428 27488 8468 27532
rect 18700 27488 18740 27616
rect 21424 27596 21504 27616
rect 19459 27572 19517 27573
rect 19075 27532 19084 27572
rect 19124 27532 19468 27572
rect 19508 27532 19517 27572
rect 19459 27531 19517 27532
rect 20995 27488 21053 27489
rect 0 27448 2956 27488
rect 2996 27448 3005 27488
rect 3331 27448 3340 27488
rect 3380 27448 5164 27488
rect 5204 27448 5356 27488
rect 5396 27448 5405 27488
rect 8419 27448 8428 27488
rect 8468 27448 10348 27488
rect 10388 27448 10397 27488
rect 10723 27448 10732 27488
rect 10772 27448 11212 27488
rect 11252 27448 11261 27488
rect 14563 27448 14572 27488
rect 14612 27448 15916 27488
rect 15956 27448 15965 27488
rect 18700 27448 21004 27488
rect 21044 27448 21053 27488
rect 0 27428 80 27448
rect 20995 27447 21053 27448
rect 11395 27404 11453 27405
rect 3523 27364 3532 27404
rect 3572 27364 6604 27404
rect 6644 27364 6653 27404
rect 8707 27364 8716 27404
rect 8756 27364 10060 27404
rect 10100 27364 10109 27404
rect 11395 27364 11404 27404
rect 11444 27364 12556 27404
rect 12596 27364 12605 27404
rect 16195 27364 16204 27404
rect 16244 27364 19756 27404
rect 19796 27364 19805 27404
rect 11395 27363 11453 27364
rect 1987 27320 2045 27321
rect 2467 27320 2525 27321
rect 11107 27320 11165 27321
rect 21424 27320 21504 27340
rect 1987 27280 1996 27320
rect 2036 27280 2476 27320
rect 2516 27280 5932 27320
rect 5972 27280 5981 27320
rect 6499 27280 6508 27320
rect 6548 27280 11116 27320
rect 11156 27280 11165 27320
rect 1987 27279 2045 27280
rect 2467 27279 2525 27280
rect 11107 27279 11165 27280
rect 15436 27280 21504 27320
rect 15436 27236 15476 27280
rect 21424 27260 21504 27280
rect 16867 27236 16925 27237
rect 3679 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 4065 27236
rect 5731 27196 5740 27236
rect 5780 27196 6604 27236
rect 6644 27196 7756 27236
rect 7796 27196 8236 27236
rect 8276 27196 8285 27236
rect 10051 27196 10060 27236
rect 10100 27196 12364 27236
rect 12404 27196 12652 27236
rect 12692 27196 12701 27236
rect 14755 27196 14764 27236
rect 14804 27196 15188 27236
rect 15427 27196 15436 27236
rect 15476 27196 15485 27236
rect 16579 27196 16588 27236
rect 16628 27196 16876 27236
rect 16916 27196 18412 27236
rect 18452 27196 18461 27236
rect 18799 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 19185 27236
rect 8227 27152 8285 27153
rect 15043 27152 15101 27153
rect 7939 27112 7948 27152
rect 7988 27112 8236 27152
rect 8276 27112 8285 27152
rect 14947 27112 14956 27152
rect 14996 27112 15052 27152
rect 15092 27112 15101 27152
rect 15148 27152 15188 27196
rect 16588 27152 16628 27196
rect 16867 27195 16925 27196
rect 15148 27112 16628 27152
rect 17251 27112 17260 27152
rect 17300 27112 17452 27152
rect 17492 27112 17501 27152
rect 8227 27111 8285 27112
rect 15043 27111 15101 27112
rect 14851 27068 14909 27069
rect 17443 27068 17501 27069
rect 2500 27028 4396 27068
rect 4436 27028 4445 27068
rect 5635 27028 5644 27068
rect 5684 27028 6316 27068
rect 6356 27028 6365 27068
rect 11320 27028 14860 27068
rect 14900 27028 17452 27068
rect 17492 27028 17501 27068
rect 2500 26984 2540 27028
rect 11320 26984 11360 27028
rect 14851 27027 14909 27028
rect 17443 27027 17501 27028
rect 21424 26984 21504 27004
rect 1315 26944 1324 26984
rect 1364 26944 2540 26984
rect 3619 26944 3628 26984
rect 3668 26944 11360 26984
rect 12451 26944 12460 26984
rect 12500 26944 19412 26984
rect 20515 26944 20524 26984
rect 20564 26944 21504 26984
rect 16963 26900 17021 26901
rect 19372 26900 19412 26944
rect 21424 26924 21504 26944
rect 7276 26860 7468 26900
rect 7508 26860 7517 26900
rect 8515 26860 8524 26900
rect 8564 26860 15244 26900
rect 15284 26860 15293 26900
rect 16963 26860 16972 26900
rect 17012 26860 17356 26900
rect 17396 26860 17405 26900
rect 19363 26860 19372 26900
rect 19412 26860 19421 26900
rect 0 26816 80 26836
rect 2467 26816 2525 26817
rect 5635 26816 5693 26817
rect 0 26776 1228 26816
rect 1268 26776 1277 26816
rect 1987 26776 1996 26816
rect 2036 26776 2476 26816
rect 2516 26776 2525 26816
rect 4579 26776 4588 26816
rect 4628 26776 4876 26816
rect 4916 26776 4925 26816
rect 5635 26776 5644 26816
rect 5684 26776 6028 26816
rect 6068 26776 6077 26816
rect 0 26756 80 26776
rect 2467 26775 2525 26776
rect 5635 26775 5693 26776
rect 2563 26692 2572 26732
rect 2612 26692 2860 26732
rect 2900 26692 3244 26732
rect 3284 26692 3293 26732
rect 7276 26648 7316 26860
rect 16963 26859 17021 26860
rect 7363 26776 7372 26816
rect 7412 26776 8332 26816
rect 8372 26776 8381 26816
rect 14851 26776 14860 26816
rect 14900 26776 15148 26816
rect 15188 26776 15197 26816
rect 16675 26776 16684 26816
rect 16724 26776 16876 26816
rect 16916 26776 16925 26816
rect 11320 26692 12748 26732
rect 12788 26692 12797 26732
rect 14755 26692 14764 26732
rect 14804 26692 14813 26732
rect 19459 26692 19468 26732
rect 19508 26692 20948 26732
rect 3043 26608 3052 26648
rect 3092 26608 3628 26648
rect 3668 26608 3677 26648
rect 5827 26608 5836 26648
rect 5876 26608 7276 26648
rect 7316 26608 7325 26648
rect 2275 26480 2333 26481
rect 2190 26440 2284 26480
rect 2324 26440 2333 26480
rect 4919 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 5305 26480
rect 6883 26440 6892 26480
rect 6932 26440 7852 26480
rect 7892 26440 7901 26480
rect 9091 26440 9100 26480
rect 9140 26440 10636 26480
rect 10676 26440 10685 26480
rect 2275 26439 2333 26440
rect 9187 26396 9245 26397
rect 11320 26396 11360 26692
rect 14764 26648 14804 26692
rect 20908 26648 20948 26692
rect 21424 26648 21504 26668
rect 12835 26608 12844 26648
rect 12884 26608 13516 26648
rect 13556 26608 13900 26648
rect 13940 26608 14804 26648
rect 16387 26608 16396 26648
rect 16436 26608 16724 26648
rect 16867 26608 16876 26648
rect 16916 26608 18124 26648
rect 18164 26608 18173 26648
rect 19555 26608 19564 26648
rect 19604 26608 19613 26648
rect 19939 26608 19948 26648
rect 19988 26608 20812 26648
rect 20852 26608 20861 26648
rect 20908 26608 21504 26648
rect 16684 26564 16724 26608
rect 19564 26564 19604 26608
rect 21424 26588 21504 26608
rect 12355 26524 12364 26564
rect 12404 26524 13804 26564
rect 13844 26524 13853 26564
rect 14083 26524 14092 26564
rect 14132 26524 16492 26564
rect 16532 26524 16541 26564
rect 16675 26524 16684 26564
rect 16724 26524 17740 26564
rect 17780 26524 17789 26564
rect 19564 26524 20524 26564
rect 20564 26524 20573 26564
rect 13411 26480 13469 26481
rect 13699 26480 13757 26481
rect 13326 26440 13420 26480
rect 13460 26440 13469 26480
rect 13614 26440 13708 26480
rect 13748 26440 13757 26480
rect 14563 26440 14572 26480
rect 14612 26440 14956 26480
rect 14996 26440 15005 26480
rect 16963 26440 16972 26480
rect 17012 26440 18988 26480
rect 19028 26440 19037 26480
rect 20039 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20425 26480
rect 13411 26439 13469 26440
rect 13699 26439 13757 26440
rect 1987 26356 1996 26396
rect 2036 26356 2540 26396
rect 3139 26356 3148 26396
rect 3188 26356 3820 26396
rect 3860 26356 3869 26396
rect 5068 26356 9196 26396
rect 9236 26356 11360 26396
rect 12643 26356 12652 26396
rect 12692 26356 13324 26396
rect 13364 26356 13373 26396
rect 18403 26356 18412 26396
rect 18452 26356 19276 26396
rect 19316 26356 19325 26396
rect 1411 26312 1469 26313
rect 1326 26272 1420 26312
rect 1460 26272 1469 26312
rect 1411 26271 1469 26272
rect 2500 26228 2540 26356
rect 5068 26312 5108 26356
rect 9187 26355 9245 26356
rect 21424 26312 21504 26332
rect 3427 26272 3436 26312
rect 3476 26272 4204 26312
rect 4244 26272 4253 26312
rect 5059 26272 5068 26312
rect 5108 26272 5117 26312
rect 8515 26272 8524 26312
rect 8564 26272 9292 26312
rect 9332 26272 9341 26312
rect 17059 26272 17068 26312
rect 17108 26272 17260 26312
rect 17300 26272 17309 26312
rect 18691 26272 18700 26312
rect 18740 26272 18892 26312
rect 18932 26272 18941 26312
rect 20140 26272 21504 26312
rect 7075 26228 7133 26229
rect 20140 26228 20180 26272
rect 21424 26252 21504 26272
rect 1219 26188 1228 26228
rect 1268 26188 1900 26228
rect 1940 26188 1949 26228
rect 2500 26188 7084 26228
rect 7124 26188 7133 26228
rect 15715 26188 15724 26228
rect 15764 26188 20180 26228
rect 7075 26187 7133 26188
rect 0 26144 80 26164
rect 259 26144 317 26145
rect 19747 26144 19805 26145
rect 0 26104 268 26144
rect 308 26104 317 26144
rect 1315 26104 1324 26144
rect 1364 26104 3148 26144
rect 3188 26104 3197 26144
rect 8323 26104 8332 26144
rect 8372 26104 9964 26144
rect 10004 26104 11308 26144
rect 11348 26104 11357 26144
rect 11779 26104 11788 26144
rect 11828 26104 12844 26144
rect 12884 26104 12893 26144
rect 13603 26104 13612 26144
rect 13652 26104 13996 26144
rect 14036 26104 17068 26144
rect 17108 26104 17117 26144
rect 18115 26104 18124 26144
rect 18164 26104 18892 26144
rect 18932 26104 18941 26144
rect 19662 26104 19756 26144
rect 19796 26104 19805 26144
rect 0 26084 80 26104
rect 259 26103 317 26104
rect 19747 26103 19805 26104
rect 3523 26060 3581 26061
rect 16291 26060 16349 26061
rect 2851 26020 2860 26060
rect 2900 26020 3244 26060
rect 3284 26020 3293 26060
rect 3523 26020 3532 26060
rect 3572 26020 15668 26060
rect 3244 25976 3284 26020
rect 3523 26019 3581 26020
rect 4579 25976 4637 25977
rect 8035 25976 8093 25977
rect 15628 25976 15668 26020
rect 16291 26020 16300 26060
rect 16340 26020 16876 26060
rect 16916 26020 16925 26060
rect 16291 26019 16349 26020
rect 16675 25976 16733 25977
rect 17059 25976 17117 25977
rect 20515 25976 20573 25977
rect 21424 25976 21504 25996
rect 3244 25936 3532 25976
rect 3572 25936 3581 25976
rect 4579 25936 4588 25976
rect 4628 25936 7084 25976
rect 7124 25936 8044 25976
rect 8084 25936 12076 25976
rect 12116 25936 12125 25976
rect 15628 25936 16684 25976
rect 16724 25936 17068 25976
rect 17108 25936 17260 25976
rect 17300 25936 17309 25976
rect 20515 25936 20524 25976
rect 20564 25936 21504 25976
rect 4579 25935 4637 25936
rect 8035 25935 8093 25936
rect 16675 25935 16733 25936
rect 17059 25935 17117 25936
rect 20515 25935 20573 25936
rect 21424 25916 21504 25936
rect 19555 25892 19613 25893
rect 1507 25852 1516 25892
rect 1556 25852 2540 25892
rect 3235 25852 3244 25892
rect 3284 25852 3820 25892
rect 3860 25852 3869 25892
rect 11587 25852 11596 25892
rect 11636 25852 13132 25892
rect 13172 25852 13181 25892
rect 15811 25852 15820 25892
rect 15860 25852 19180 25892
rect 19220 25852 19229 25892
rect 19470 25852 19564 25892
rect 19604 25852 19613 25892
rect 2500 25556 2540 25852
rect 19555 25851 19613 25852
rect 5923 25808 5981 25809
rect 7459 25808 7517 25809
rect 5923 25768 5932 25808
rect 5972 25768 7468 25808
rect 7508 25768 8332 25808
rect 8372 25768 8381 25808
rect 16387 25768 16396 25808
rect 16436 25768 17932 25808
rect 17972 25768 17981 25808
rect 5923 25767 5981 25768
rect 7459 25767 7517 25768
rect 18691 25724 18749 25725
rect 3679 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 4065 25724
rect 6019 25684 6028 25724
rect 6068 25684 6412 25724
rect 6452 25684 6461 25724
rect 12739 25684 12748 25724
rect 12788 25684 13324 25724
rect 13364 25684 13373 25724
rect 16867 25684 16876 25724
rect 16916 25684 18700 25724
rect 18740 25684 18749 25724
rect 18799 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 19185 25724
rect 18691 25683 18749 25684
rect 13027 25640 13085 25641
rect 6220 25600 7124 25640
rect 12931 25600 12940 25640
rect 12980 25600 13036 25640
rect 13076 25600 13085 25640
rect 2500 25516 4012 25556
rect 4052 25516 4780 25556
rect 4820 25516 4829 25556
rect 0 25472 80 25492
rect 6220 25472 6260 25600
rect 7084 25472 7124 25600
rect 13027 25599 13085 25600
rect 16867 25640 16925 25641
rect 17443 25640 17501 25641
rect 19267 25640 19325 25641
rect 21424 25640 21504 25660
rect 16867 25600 16876 25640
rect 16916 25600 17452 25640
rect 17492 25600 17740 25640
rect 17780 25600 17789 25640
rect 18019 25600 18028 25640
rect 18068 25600 19124 25640
rect 16867 25599 16925 25600
rect 17443 25599 17501 25600
rect 19084 25556 19124 25600
rect 19267 25600 19276 25640
rect 19316 25600 21504 25640
rect 19267 25599 19325 25600
rect 21424 25580 21504 25600
rect 10819 25516 10828 25556
rect 10868 25516 12556 25556
rect 12596 25516 15148 25556
rect 15188 25516 15197 25556
rect 17164 25516 18316 25556
rect 18356 25516 18365 25556
rect 19075 25516 19084 25556
rect 19124 25516 19133 25556
rect 14851 25472 14909 25473
rect 0 25432 6260 25472
rect 6316 25432 6988 25472
rect 7028 25432 7037 25472
rect 7084 25432 12460 25472
rect 12500 25432 12509 25472
rect 13036 25432 14860 25472
rect 14900 25432 14909 25472
rect 0 25412 80 25432
rect 2179 25348 2188 25388
rect 2228 25348 2860 25388
rect 2900 25348 2909 25388
rect 3139 25348 3148 25388
rect 3188 25348 5548 25388
rect 5588 25348 5836 25388
rect 5876 25348 5885 25388
rect 6316 25304 6356 25432
rect 13036 25388 13076 25432
rect 14851 25431 14909 25432
rect 8707 25348 8716 25388
rect 8756 25348 8765 25388
rect 13027 25348 13036 25388
rect 13076 25348 13085 25388
rect 13507 25348 13516 25388
rect 13556 25348 13565 25388
rect 13795 25348 13804 25388
rect 13844 25348 14092 25388
rect 14132 25348 14141 25388
rect 1603 25264 1612 25304
rect 1652 25264 2540 25304
rect 2659 25264 2668 25304
rect 2708 25264 3436 25304
rect 3476 25264 3485 25304
rect 3532 25264 4492 25304
rect 4532 25264 6356 25304
rect 7075 25264 7084 25304
rect 7124 25264 7756 25304
rect 7796 25264 7805 25304
rect 2500 25220 2540 25264
rect 3532 25220 3572 25264
rect 5443 25220 5501 25221
rect 2500 25180 2804 25220
rect 2851 25180 2860 25220
rect 2900 25180 3244 25220
rect 3284 25180 3293 25220
rect 3340 25180 3572 25220
rect 4387 25180 4396 25220
rect 4436 25180 5068 25220
rect 5108 25180 5117 25220
rect 5347 25180 5356 25220
rect 5396 25180 5452 25220
rect 5492 25180 5501 25220
rect 2764 25136 2804 25180
rect 3340 25136 3380 25180
rect 5443 25179 5501 25180
rect 5347 25136 5405 25137
rect 1315 25096 1324 25136
rect 1364 25096 1900 25136
rect 1940 25096 1949 25136
rect 2764 25096 3380 25136
rect 4963 25096 4972 25136
rect 5012 25096 5356 25136
rect 5396 25096 5405 25136
rect 5347 25095 5405 25096
rect 6316 25052 6356 25264
rect 7555 25180 7564 25220
rect 7604 25180 8428 25220
rect 8468 25180 8477 25220
rect 8716 25052 8756 25348
rect 13411 25304 13469 25305
rect 13326 25264 13420 25304
rect 13460 25264 13469 25304
rect 13411 25263 13469 25264
rect 13516 25220 13556 25348
rect 14083 25304 14141 25305
rect 13987 25264 13996 25304
rect 14036 25264 14092 25304
rect 14132 25264 14141 25304
rect 17164 25304 17204 25516
rect 17251 25432 17260 25472
rect 17300 25432 17309 25472
rect 17635 25432 17644 25472
rect 17684 25432 18028 25472
rect 18068 25432 18077 25472
rect 19171 25432 19180 25472
rect 19220 25432 19468 25472
rect 19508 25432 19517 25472
rect 19651 25432 19660 25472
rect 19700 25432 19852 25472
rect 19892 25432 19901 25472
rect 17260 25388 17300 25432
rect 17260 25348 17452 25388
rect 17492 25348 17501 25388
rect 17923 25348 17932 25388
rect 17972 25348 19756 25388
rect 19796 25348 19805 25388
rect 21424 25304 21504 25324
rect 17164 25264 17253 25304
rect 17293 25264 17302 25304
rect 17347 25264 17356 25304
rect 17396 25264 21504 25304
rect 14083 25263 14141 25264
rect 21424 25244 21504 25264
rect 18595 25220 18653 25221
rect 11491 25180 11500 25220
rect 11540 25180 14284 25220
rect 14324 25180 14333 25220
rect 15427 25180 15436 25220
rect 15476 25180 17548 25220
rect 17588 25180 18124 25220
rect 18164 25180 18173 25220
rect 18403 25180 18412 25220
rect 18452 25180 18604 25220
rect 18644 25180 18653 25220
rect 18595 25179 18653 25180
rect 18787 25220 18845 25221
rect 18787 25180 18796 25220
rect 18836 25180 18892 25220
rect 18932 25180 18941 25220
rect 18787 25179 18845 25180
rect 12643 25096 12652 25136
rect 12692 25096 13228 25136
rect 13268 25096 13277 25136
rect 14083 25096 14092 25136
rect 14132 25096 14476 25136
rect 14516 25096 14525 25136
rect 16003 25096 16012 25136
rect 16052 25096 16300 25136
rect 16340 25096 16349 25136
rect 19459 25096 19468 25136
rect 19508 25096 20044 25136
rect 20084 25096 20093 25136
rect 18115 25052 18173 25053
rect 20899 25052 20957 25053
rect 6307 25012 6316 25052
rect 6356 25012 6365 25052
rect 8716 25012 16780 25052
rect 16820 25012 16829 25052
rect 18115 25012 18124 25052
rect 18164 25012 20908 25052
rect 20948 25012 20957 25052
rect 18115 25011 18173 25012
rect 20899 25011 20957 25012
rect 6979 24968 7037 24969
rect 15331 24968 15389 24969
rect 21424 24968 21504 24988
rect 1411 24928 1420 24968
rect 1460 24928 4108 24968
rect 4148 24928 4157 24968
rect 4919 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 5305 24968
rect 5443 24928 5452 24968
rect 5492 24928 6988 24968
rect 7028 24928 7037 24968
rect 12931 24928 12940 24968
rect 12980 24928 15340 24968
rect 15380 24928 15389 24968
rect 20039 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20425 24968
rect 20515 24928 20524 24968
rect 20564 24928 21504 24968
rect 6979 24927 7037 24928
rect 15331 24927 15389 24928
rect 21424 24908 21504 24928
rect 13027 24884 13085 24885
rect 3523 24844 3532 24884
rect 3572 24844 5740 24884
rect 5780 24844 5789 24884
rect 13027 24844 13036 24884
rect 13076 24844 16108 24884
rect 16148 24844 18604 24884
rect 18644 24844 18653 24884
rect 19267 24844 19276 24884
rect 19316 24844 19852 24884
rect 19892 24844 19901 24884
rect 13027 24843 13085 24844
rect 0 24800 80 24820
rect 19555 24800 19613 24801
rect 19852 24800 19892 24844
rect 0 24760 3052 24800
rect 3092 24760 3101 24800
rect 7555 24760 7564 24800
rect 7604 24760 8524 24800
rect 8564 24760 8573 24800
rect 11971 24760 11980 24800
rect 12020 24760 13036 24800
rect 13076 24760 13228 24800
rect 13268 24760 13277 24800
rect 15427 24760 15436 24800
rect 15476 24760 15724 24800
rect 15764 24760 15773 24800
rect 15907 24760 15916 24800
rect 15956 24760 15965 24800
rect 18211 24760 18220 24800
rect 18260 24760 19372 24800
rect 19412 24760 19421 24800
rect 19555 24760 19564 24800
rect 19604 24760 19660 24800
rect 19700 24760 19709 24800
rect 19852 24760 20044 24800
rect 20084 24760 20093 24800
rect 0 24740 80 24760
rect 2467 24716 2525 24717
rect 6595 24716 6653 24717
rect 1123 24676 1132 24716
rect 1172 24676 2476 24716
rect 2516 24676 6124 24716
rect 6164 24676 6604 24716
rect 6644 24676 6653 24716
rect 12067 24676 12076 24716
rect 12116 24676 15244 24716
rect 15284 24676 15293 24716
rect 2467 24675 2525 24676
rect 6595 24675 6653 24676
rect 2947 24632 3005 24633
rect 5347 24632 5405 24633
rect 7363 24632 7421 24633
rect 8227 24632 8285 24633
rect 1219 24592 1228 24632
rect 1268 24592 2956 24632
rect 2996 24592 3916 24632
rect 3956 24592 3965 24632
rect 5262 24592 5356 24632
rect 5396 24592 5405 24632
rect 6691 24592 6700 24632
rect 6740 24592 7372 24632
rect 7412 24592 7421 24632
rect 7747 24592 7756 24632
rect 7796 24592 7948 24632
rect 7988 24592 8236 24632
rect 8276 24592 8285 24632
rect 2947 24591 3005 24592
rect 5347 24591 5405 24592
rect 7363 24591 7421 24592
rect 8227 24591 8285 24592
rect 9283 24632 9341 24633
rect 10147 24632 10205 24633
rect 15916 24632 15956 24760
rect 19555 24759 19613 24760
rect 19267 24632 19325 24633
rect 21424 24632 21504 24652
rect 9283 24592 9292 24632
rect 9332 24592 10156 24632
rect 10196 24592 10205 24632
rect 13507 24592 13516 24632
rect 13556 24592 14476 24632
rect 14516 24592 14525 24632
rect 15715 24592 15724 24632
rect 15764 24592 15956 24632
rect 16483 24592 16492 24632
rect 16532 24592 18988 24632
rect 19028 24592 19037 24632
rect 19267 24592 19276 24632
rect 19316 24592 21504 24632
rect 9283 24591 9341 24592
rect 10147 24591 10205 24592
rect 19267 24591 19325 24592
rect 21424 24572 21504 24592
rect 4771 24548 4829 24549
rect 13987 24548 14045 24549
rect 20899 24548 20957 24549
rect 4771 24508 4780 24548
rect 4820 24508 4876 24548
rect 4916 24508 4925 24548
rect 6892 24508 13996 24548
rect 14036 24508 14045 24548
rect 14755 24508 14764 24548
rect 14804 24508 17932 24548
rect 17972 24508 17981 24548
rect 19075 24508 19084 24548
rect 19124 24508 20908 24548
rect 20948 24508 20957 24548
rect 4771 24507 4829 24508
rect 6892 24464 6932 24508
rect 13987 24507 14045 24508
rect 20899 24507 20957 24508
rect 9955 24464 10013 24465
rect 1987 24424 1996 24464
rect 2036 24424 6932 24464
rect 9870 24424 9964 24464
rect 10004 24424 10013 24464
rect 11203 24424 11212 24464
rect 11252 24424 12844 24464
rect 12884 24424 12893 24464
rect 9955 24423 10013 24424
rect 6019 24380 6077 24381
rect 13996 24380 14036 24507
rect 14851 24424 14860 24464
rect 14900 24424 17356 24464
rect 17396 24424 17405 24464
rect 20035 24424 20044 24464
rect 20084 24424 20524 24464
rect 20564 24424 20573 24464
rect 21187 24380 21245 24381
rect 20 24340 4244 24380
rect 4387 24340 4396 24380
rect 4436 24340 5836 24380
rect 5876 24340 5885 24380
rect 6019 24340 6028 24380
rect 6068 24340 6124 24380
rect 6164 24340 6173 24380
rect 8611 24340 8620 24380
rect 8660 24340 11596 24380
rect 11636 24340 11645 24380
rect 13987 24340 13996 24380
rect 14036 24340 14045 24380
rect 16003 24340 16012 24380
rect 16052 24340 17932 24380
rect 17972 24340 17981 24380
rect 18979 24340 18988 24380
rect 19028 24340 21196 24380
rect 21236 24340 21245 24380
rect 20 24296 60 24340
rect 20 24256 116 24296
rect 76 24148 116 24256
rect 4204 24212 4244 24340
rect 6019 24339 6077 24340
rect 21187 24339 21245 24340
rect 21424 24296 21504 24316
rect 4963 24256 4972 24296
rect 5012 24256 14092 24296
rect 14132 24256 14141 24296
rect 16588 24256 19564 24296
rect 19604 24256 19613 24296
rect 20803 24256 20812 24296
rect 20852 24256 21504 24296
rect 5827 24212 5885 24213
rect 16588 24212 16628 24256
rect 21424 24236 21504 24256
rect 3679 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 4065 24212
rect 4204 24172 5836 24212
rect 5876 24172 5885 24212
rect 7939 24172 7948 24212
rect 7988 24172 8620 24212
rect 8660 24172 8669 24212
rect 13507 24172 13516 24212
rect 13556 24172 16588 24212
rect 16628 24172 16637 24212
rect 18799 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 19185 24212
rect 5827 24171 5885 24172
rect 0 24088 116 24148
rect 9763 24088 9772 24128
rect 9812 24088 11692 24128
rect 11732 24088 11741 24128
rect 0 24068 80 24088
rect 9859 24044 9917 24045
rect 10723 24044 10781 24045
rect 3043 24004 3052 24044
rect 3092 24004 3628 24044
rect 3668 24004 3677 24044
rect 9187 24004 9196 24044
rect 9236 24004 9868 24044
rect 9908 24004 9917 24044
rect 10339 24004 10348 24044
rect 10388 24004 10732 24044
rect 10772 24004 10781 24044
rect 15811 24004 15820 24044
rect 15860 24004 16108 24044
rect 16148 24004 16157 24044
rect 9859 24003 9917 24004
rect 10723 24003 10781 24004
rect 9091 23960 9149 23961
rect 14083 23960 14141 23961
rect 18691 23960 18749 23961
rect 21424 23960 21504 23980
rect 4579 23920 4588 23960
rect 4628 23920 5644 23960
rect 5684 23920 5693 23960
rect 6883 23920 6892 23960
rect 6932 23920 7276 23960
rect 7316 23920 7325 23960
rect 7459 23920 7468 23960
rect 7508 23920 7852 23960
rect 7892 23920 7901 23960
rect 9091 23920 9100 23960
rect 9140 23920 9292 23960
rect 9332 23920 9341 23960
rect 9571 23920 9580 23960
rect 9620 23920 9964 23960
rect 10004 23920 10013 23960
rect 10147 23920 10156 23960
rect 10196 23920 10636 23960
rect 10676 23920 10685 23960
rect 13219 23920 13228 23960
rect 13268 23920 14092 23960
rect 14132 23920 15148 23960
rect 15188 23920 15197 23960
rect 15331 23920 15340 23960
rect 15380 23920 15916 23960
rect 15956 23920 16588 23960
rect 16628 23920 16637 23960
rect 17347 23920 17356 23960
rect 17396 23920 17548 23960
rect 17588 23920 17597 23960
rect 18595 23920 18604 23960
rect 18644 23920 18700 23960
rect 18740 23920 18749 23960
rect 19651 23920 19660 23960
rect 19700 23920 20180 23960
rect 9091 23919 9149 23920
rect 7363 23876 7421 23877
rect 1795 23836 1804 23876
rect 1844 23836 1996 23876
rect 2036 23836 5972 23876
rect 2755 23752 2764 23792
rect 2804 23752 3148 23792
rect 3188 23752 3197 23792
rect 3523 23752 3532 23792
rect 3572 23752 4012 23792
rect 4052 23752 4061 23792
rect 1891 23668 1900 23708
rect 1940 23668 3916 23708
rect 3956 23668 3965 23708
rect 2083 23584 2092 23624
rect 2132 23584 4588 23624
rect 4628 23584 4637 23624
rect 5059 23584 5068 23624
rect 5108 23584 5117 23624
rect 4099 23540 4157 23541
rect 5068 23540 5108 23584
rect 1987 23500 1996 23540
rect 2036 23500 2380 23540
rect 2420 23500 2429 23540
rect 3331 23500 3340 23540
rect 3380 23500 4108 23540
rect 4148 23500 4492 23540
rect 4532 23500 4541 23540
rect 4588 23500 5108 23540
rect 5932 23540 5972 23836
rect 7363 23836 7372 23876
rect 7412 23836 9196 23876
rect 9236 23836 9676 23876
rect 9716 23836 9725 23876
rect 7363 23835 7421 23836
rect 10156 23792 10196 23920
rect 14083 23919 14141 23920
rect 18691 23919 18749 23920
rect 20140 23876 20180 23920
rect 21004 23920 21504 23960
rect 21004 23876 21044 23920
rect 21424 23900 21504 23920
rect 13603 23836 13612 23876
rect 13652 23836 13900 23876
rect 13940 23836 16396 23876
rect 16436 23836 16445 23876
rect 20140 23836 21044 23876
rect 11011 23792 11069 23793
rect 17059 23792 17117 23793
rect 6019 23752 6028 23792
rect 6068 23752 6220 23792
rect 6260 23752 10196 23792
rect 10926 23752 11020 23792
rect 11060 23752 11069 23792
rect 11011 23751 11069 23752
rect 11116 23752 11308 23792
rect 11348 23752 11357 23792
rect 12643 23752 12652 23792
rect 12692 23752 14476 23792
rect 14516 23752 14525 23792
rect 17059 23752 17068 23792
rect 17108 23752 19276 23792
rect 19316 23752 19564 23792
rect 19604 23752 19613 23792
rect 7363 23708 7421 23709
rect 11116 23708 11156 23752
rect 17059 23751 17117 23752
rect 12259 23708 12317 23709
rect 7267 23668 7276 23708
rect 7316 23668 7372 23708
rect 7412 23668 7421 23708
rect 9667 23668 9676 23708
rect 9716 23668 11156 23708
rect 11212 23668 12268 23708
rect 12308 23668 12317 23708
rect 7363 23667 7421 23668
rect 11212 23624 11252 23668
rect 12259 23667 12317 23668
rect 9475 23584 9484 23624
rect 9524 23584 11252 23624
rect 11299 23624 11357 23625
rect 19363 23624 19421 23625
rect 21424 23624 21504 23644
rect 11299 23584 11308 23624
rect 11348 23584 11596 23624
rect 11636 23584 11645 23624
rect 15235 23584 15244 23624
rect 15284 23584 17164 23624
rect 17204 23584 17213 23624
rect 19363 23584 19372 23624
rect 19412 23584 21504 23624
rect 11299 23583 11357 23584
rect 19363 23583 19421 23584
rect 21424 23564 21504 23584
rect 13123 23540 13181 23541
rect 5932 23500 12556 23540
rect 12596 23500 13132 23540
rect 13172 23500 13181 23540
rect 4099 23499 4157 23500
rect 0 23456 80 23476
rect 163 23456 221 23457
rect 4588 23456 4628 23500
rect 13123 23499 13181 23500
rect 0 23416 172 23456
rect 212 23416 221 23456
rect 4579 23416 4588 23456
rect 4628 23416 4637 23456
rect 4919 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 5305 23456
rect 9571 23416 9580 23456
rect 9620 23416 9629 23456
rect 11299 23416 11308 23456
rect 11348 23416 11500 23456
rect 11540 23416 11549 23456
rect 20039 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20425 23456
rect 0 23396 80 23416
rect 163 23415 221 23416
rect 7555 23372 7613 23373
rect 9580 23372 9620 23416
rect 11299 23372 11357 23373
rect 7555 23332 7564 23372
rect 7604 23332 7948 23372
rect 7988 23332 7997 23372
rect 9379 23332 9388 23372
rect 9428 23332 11020 23372
rect 11060 23332 11308 23372
rect 11348 23332 11357 23372
rect 7555 23331 7613 23332
rect 11299 23331 11357 23332
rect 19363 23288 19421 23289
rect 21424 23288 21504 23308
rect 3427 23248 3436 23288
rect 3476 23248 6604 23288
rect 6644 23248 6796 23288
rect 6836 23248 6845 23288
rect 9283 23248 9292 23288
rect 9332 23248 11212 23288
rect 11252 23248 11261 23288
rect 14179 23248 14188 23288
rect 14228 23248 14476 23288
rect 14516 23248 14525 23288
rect 16387 23248 16396 23288
rect 16436 23248 16876 23288
rect 16916 23248 19121 23288
rect 19161 23248 19372 23288
rect 19412 23248 19421 23288
rect 19843 23248 19852 23288
rect 19892 23248 20140 23288
rect 20180 23248 20189 23288
rect 20236 23248 21504 23288
rect 19363 23247 19421 23248
rect 4579 23204 4637 23205
rect 7363 23204 7421 23205
rect 16483 23204 16541 23205
rect 17347 23204 17405 23205
rect 20236 23204 20276 23248
rect 21424 23228 21504 23248
rect 1315 23164 1324 23204
rect 1364 23164 2540 23204
rect 3619 23164 3628 23204
rect 3668 23164 4204 23204
rect 4244 23164 4253 23204
rect 4483 23164 4492 23204
rect 4532 23164 4588 23204
rect 4628 23164 4637 23204
rect 5923 23164 5932 23204
rect 5972 23164 6508 23204
rect 6548 23164 7372 23204
rect 7412 23164 7421 23204
rect 7555 23164 7564 23204
rect 7604 23164 10348 23204
rect 10388 23164 10397 23204
rect 12835 23164 12844 23204
rect 12884 23164 13132 23204
rect 13172 23164 13181 23204
rect 16483 23164 16492 23204
rect 16532 23164 17356 23204
rect 17396 23164 17452 23204
rect 17492 23164 17501 23204
rect 20140 23164 20276 23204
rect 2500 23120 2540 23164
rect 4579 23163 4637 23164
rect 7363 23163 7421 23164
rect 16483 23163 16541 23164
rect 17347 23163 17405 23164
rect 11107 23120 11165 23121
rect 2500 23080 3148 23120
rect 3188 23080 3820 23120
rect 3860 23080 5548 23120
rect 5588 23080 5597 23120
rect 7075 23080 7084 23120
rect 7124 23080 7948 23120
rect 7988 23080 7997 23120
rect 8515 23080 8524 23120
rect 8564 23080 8716 23120
rect 8756 23080 8765 23120
rect 8995 23080 9004 23120
rect 9044 23080 9772 23120
rect 9812 23080 9821 23120
rect 11022 23080 11116 23120
rect 11156 23080 11165 23120
rect 13411 23080 13420 23120
rect 13460 23080 13612 23120
rect 13652 23080 13661 23120
rect 16195 23080 16204 23120
rect 16244 23080 17644 23120
rect 17684 23080 17693 23120
rect 18115 23080 18124 23120
rect 18164 23080 18508 23120
rect 18548 23080 19852 23120
rect 19892 23080 19901 23120
rect 11107 23079 11165 23080
rect 17443 23036 17501 23037
rect 20140 23036 20180 23164
rect 7171 22996 7180 23036
rect 7220 22996 7508 23036
rect 11683 22996 11692 23036
rect 11732 22996 15244 23036
rect 15284 22996 15293 23036
rect 16483 22996 16492 23036
rect 16532 22996 16876 23036
rect 16916 22996 16925 23036
rect 17443 22996 17452 23036
rect 17492 22996 20180 23036
rect 7468 22952 7508 22996
rect 17443 22995 17501 22996
rect 13027 22952 13085 22953
rect 21424 22952 21504 22972
rect 4099 22912 4108 22952
rect 4148 22912 6892 22952
rect 6932 22912 6941 22952
rect 7459 22912 7468 22952
rect 7508 22912 7517 22952
rect 8515 22912 8524 22952
rect 8564 22912 12652 22952
rect 12692 22912 12701 22952
rect 12942 22912 13036 22952
rect 13076 22912 13085 22952
rect 17251 22912 17260 22952
rect 17300 22912 18220 22952
rect 18260 22912 18269 22952
rect 21379 22912 21388 22952
rect 21428 22912 21504 22952
rect 13027 22911 13085 22912
rect 21424 22892 21504 22912
rect 19651 22868 19709 22869
rect 4771 22828 4780 22868
rect 4820 22828 6028 22868
rect 6068 22828 6077 22868
rect 9379 22828 9388 22868
rect 9428 22828 9868 22868
rect 9908 22828 9917 22868
rect 19566 22828 19660 22868
rect 19700 22828 19709 22868
rect 19651 22827 19709 22828
rect 0 22784 80 22804
rect 0 22744 11884 22784
rect 11924 22744 11933 22784
rect 13219 22744 13228 22784
rect 13268 22744 13420 22784
rect 13460 22744 13469 22784
rect 0 22724 80 22744
rect 14755 22700 14813 22701
rect 18595 22700 18653 22701
rect 3679 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 4065 22700
rect 4771 22660 4780 22700
rect 4820 22660 5452 22700
rect 5492 22660 5501 22700
rect 5635 22660 5644 22700
rect 5684 22660 6508 22700
rect 6548 22660 6557 22700
rect 7459 22660 7468 22700
rect 7508 22660 14764 22700
rect 14804 22660 14813 22700
rect 16003 22660 16012 22700
rect 16052 22660 16396 22700
rect 16436 22660 16445 22700
rect 18403 22660 18412 22700
rect 18452 22660 18604 22700
rect 18644 22660 18653 22700
rect 18799 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 19185 22700
rect 14755 22659 14813 22660
rect 18595 22659 18653 22660
rect 9571 22616 9629 22617
rect 21424 22616 21504 22636
rect 2659 22576 2668 22616
rect 2708 22576 4300 22616
rect 4340 22576 4349 22616
rect 8899 22576 8908 22616
rect 8948 22576 9580 22616
rect 9620 22576 10156 22616
rect 10196 22576 10205 22616
rect 12739 22576 12748 22616
rect 12788 22576 13132 22616
rect 13172 22576 13181 22616
rect 20803 22576 20812 22616
rect 20852 22576 21504 22616
rect 9571 22575 9629 22576
rect 21424 22556 21504 22576
rect 15811 22532 15869 22533
rect 3043 22492 3052 22532
rect 3092 22492 3956 22532
rect 4003 22492 4012 22532
rect 4052 22492 5356 22532
rect 5396 22492 5405 22532
rect 9187 22492 9196 22532
rect 9236 22492 9772 22532
rect 9812 22492 9821 22532
rect 10243 22492 10252 22532
rect 10292 22492 12556 22532
rect 12596 22492 12605 22532
rect 12931 22492 12940 22532
rect 12980 22492 12989 22532
rect 14467 22492 14476 22532
rect 14516 22492 15148 22532
rect 15188 22492 15197 22532
rect 15715 22492 15724 22532
rect 15764 22492 15820 22532
rect 15860 22492 15869 22532
rect 3916 22448 3956 22492
rect 12940 22448 12980 22492
rect 15811 22491 15869 22492
rect 2500 22408 2860 22448
rect 2900 22408 2909 22448
rect 3907 22408 3916 22448
rect 3956 22408 3965 22448
rect 5443 22408 5452 22448
rect 5492 22408 7276 22448
rect 7316 22408 7325 22448
rect 12355 22408 12364 22448
rect 12404 22408 12692 22448
rect 12940 22408 17932 22448
rect 17972 22408 19852 22448
rect 19892 22408 19901 22448
rect 2500 22364 2540 22408
rect 7363 22364 7421 22365
rect 12652 22364 12692 22408
rect 16387 22364 16445 22365
rect 16867 22364 16925 22365
rect 2467 22324 2476 22364
rect 2516 22324 2668 22364
rect 2708 22324 2717 22364
rect 3331 22324 3340 22364
rect 3380 22324 4588 22364
rect 4628 22324 4637 22364
rect 7278 22324 7372 22364
rect 7412 22324 7421 22364
rect 12643 22324 12652 22364
rect 12692 22324 12701 22364
rect 15715 22324 15724 22364
rect 15764 22324 16108 22364
rect 16148 22324 16157 22364
rect 16387 22324 16396 22364
rect 16436 22324 16684 22364
rect 16724 22324 16876 22364
rect 16916 22324 16925 22364
rect 7363 22323 7421 22324
rect 16387 22323 16445 22324
rect 16867 22323 16925 22324
rect 2371 22280 2429 22281
rect 1315 22240 1324 22280
rect 1364 22240 2380 22280
rect 2420 22240 2429 22280
rect 2371 22239 2429 22240
rect 2659 22280 2717 22281
rect 14083 22280 14141 22281
rect 21424 22280 21504 22300
rect 2659 22240 2668 22280
rect 2708 22240 3628 22280
rect 3668 22240 3677 22280
rect 3811 22240 3820 22280
rect 3860 22240 4108 22280
rect 4148 22240 6604 22280
rect 6644 22240 6653 22280
rect 7171 22240 7180 22280
rect 7220 22240 7852 22280
rect 7892 22240 7901 22280
rect 9475 22240 9484 22280
rect 9524 22240 9868 22280
rect 9908 22240 9917 22280
rect 14083 22240 14092 22280
rect 14132 22240 14380 22280
rect 14420 22240 14572 22280
rect 14612 22240 14621 22280
rect 14755 22240 14764 22280
rect 14804 22240 15052 22280
rect 15092 22240 15101 22280
rect 15427 22240 15436 22280
rect 15476 22240 21504 22280
rect 2659 22239 2717 22240
rect 14083 22239 14141 22240
rect 21424 22220 21504 22240
rect 16867 22196 16925 22197
rect 3523 22156 3532 22196
rect 3572 22156 6892 22196
rect 6932 22156 16876 22196
rect 16916 22156 16925 22196
rect 16867 22155 16925 22156
rect 0 22112 80 22132
rect 7075 22112 7133 22113
rect 7363 22112 7421 22113
rect 13123 22112 13181 22113
rect 0 22072 2540 22112
rect 5251 22072 5260 22112
rect 5300 22072 6796 22112
rect 6836 22072 6845 22112
rect 7075 22072 7084 22112
rect 7124 22072 7372 22112
rect 7412 22072 8140 22112
rect 8180 22072 10924 22112
rect 10964 22072 10973 22112
rect 13038 22072 13132 22112
rect 13172 22072 13181 22112
rect 15331 22072 15340 22112
rect 15380 22072 15389 22112
rect 15619 22072 15628 22112
rect 15668 22072 16012 22112
rect 16052 22072 16061 22112
rect 0 22052 80 22072
rect 2500 21860 2540 22072
rect 7075 22071 7133 22072
rect 7363 22071 7421 22072
rect 13123 22071 13181 22072
rect 3235 22028 3293 22029
rect 6979 22028 7037 22029
rect 15340 22028 15380 22072
rect 3139 21988 3148 22028
rect 3188 21988 3244 22028
rect 3284 21988 3293 22028
rect 4387 21988 4396 22028
rect 4436 21988 5932 22028
rect 5972 21988 5981 22028
rect 6979 21988 6988 22028
rect 7028 21988 7276 22028
rect 7316 21988 7325 22028
rect 14764 21988 15380 22028
rect 3235 21987 3293 21988
rect 6979 21987 7037 21988
rect 4919 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 5305 21944
rect 7651 21904 7660 21944
rect 7700 21904 8332 21944
rect 8372 21904 8381 21944
rect 13699 21904 13708 21944
rect 13748 21904 14284 21944
rect 14324 21904 14668 21944
rect 14708 21904 14717 21944
rect 6691 21860 6749 21861
rect 14764 21860 14804 21988
rect 16963 21944 17021 21945
rect 21424 21944 21504 21964
rect 16878 21904 16972 21944
rect 17012 21904 17021 21944
rect 20039 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20425 21944
rect 20611 21904 20620 21944
rect 20660 21904 21504 21944
rect 16963 21903 17021 21904
rect 21424 21884 21504 21904
rect 2500 21820 6700 21860
rect 6740 21820 6749 21860
rect 7171 21820 7180 21860
rect 7220 21820 7372 21860
rect 7412 21820 7421 21860
rect 7555 21820 7564 21860
rect 7604 21820 8812 21860
rect 8852 21820 10924 21860
rect 10964 21820 11116 21860
rect 11156 21820 11165 21860
rect 14083 21820 14092 21860
rect 14132 21820 14324 21860
rect 14563 21820 14572 21860
rect 14612 21820 14804 21860
rect 6691 21819 6749 21820
rect 2947 21776 3005 21777
rect 14284 21776 14324 21820
rect 2862 21736 2956 21776
rect 2996 21736 3005 21776
rect 4195 21736 4204 21776
rect 4244 21736 4684 21776
rect 4724 21736 4733 21776
rect 5827 21736 5836 21776
rect 5876 21736 6892 21776
rect 6932 21736 7948 21776
rect 7988 21736 7997 21776
rect 8044 21736 11360 21776
rect 14275 21736 14284 21776
rect 14324 21736 14333 21776
rect 19555 21736 19564 21776
rect 19604 21736 19644 21776
rect 2947 21735 3005 21736
rect 3523 21652 3532 21692
rect 3572 21652 3724 21692
rect 3764 21652 5356 21692
rect 5396 21652 7508 21692
rect 7468 21609 7508 21652
rect 5635 21608 5693 21609
rect 7459 21608 7517 21609
rect 8044 21608 8084 21736
rect 9571 21692 9629 21693
rect 9571 21652 9580 21692
rect 9620 21652 9676 21692
rect 9716 21652 9725 21692
rect 9571 21651 9629 21652
rect 11320 21608 11360 21736
rect 15331 21692 15389 21693
rect 19564 21692 19604 21736
rect 15246 21652 15340 21692
rect 15380 21652 15389 21692
rect 16483 21652 16492 21692
rect 16532 21652 17068 21692
rect 17108 21652 17117 21692
rect 18691 21652 18700 21692
rect 18740 21652 19852 21692
rect 19892 21652 19901 21692
rect 15331 21651 15389 21652
rect 17635 21608 17693 21609
rect 20611 21608 20669 21609
rect 21424 21608 21504 21628
rect 1507 21568 1516 21608
rect 1556 21568 2540 21608
rect 0 21440 80 21460
rect 1219 21440 1277 21441
rect 0 21400 1228 21440
rect 1268 21400 1277 21440
rect 2500 21440 2540 21568
rect 2668 21568 3340 21608
rect 3380 21568 3628 21608
rect 3668 21568 3677 21608
rect 5443 21568 5452 21608
rect 5492 21568 5644 21608
rect 5684 21568 6220 21608
rect 6260 21568 6269 21608
rect 6499 21568 6508 21608
rect 6548 21568 6700 21608
rect 6740 21568 6749 21608
rect 7374 21568 7468 21608
rect 7508 21568 7517 21608
rect 8035 21568 8044 21608
rect 8084 21568 8093 21608
rect 9763 21568 9772 21608
rect 9812 21568 10732 21608
rect 10772 21568 10781 21608
rect 11320 21568 12556 21608
rect 12596 21568 12605 21608
rect 14851 21568 14860 21608
rect 14900 21568 15244 21608
rect 15284 21568 15293 21608
rect 16387 21568 16396 21608
rect 16436 21568 16876 21608
rect 16916 21568 17164 21608
rect 17204 21568 17213 21608
rect 17550 21568 17644 21608
rect 17684 21568 17693 21608
rect 19171 21568 19180 21608
rect 19220 21568 19564 21608
rect 19604 21568 19948 21608
rect 19988 21568 19997 21608
rect 20131 21568 20140 21608
rect 20180 21568 20189 21608
rect 20611 21568 20620 21608
rect 20660 21568 21504 21608
rect 2668 21524 2708 21568
rect 5635 21567 5693 21568
rect 7459 21567 7517 21568
rect 8044 21524 8084 21568
rect 17635 21567 17693 21568
rect 14371 21524 14429 21525
rect 20140 21524 20180 21568
rect 20611 21567 20669 21568
rect 21424 21548 21504 21568
rect 20995 21524 21053 21525
rect 2659 21484 2668 21524
rect 2708 21484 2717 21524
rect 2851 21484 2860 21524
rect 2900 21484 4396 21524
rect 4436 21484 4445 21524
rect 6115 21484 6124 21524
rect 6164 21484 6892 21524
rect 6932 21484 8084 21524
rect 10339 21484 10348 21524
rect 10388 21484 14380 21524
rect 14420 21484 14429 21524
rect 15427 21484 15436 21524
rect 15476 21484 15724 21524
rect 15764 21484 17260 21524
rect 17300 21484 17309 21524
rect 20140 21484 21004 21524
rect 21044 21484 21053 21524
rect 14371 21483 14429 21484
rect 2500 21400 5548 21440
rect 5588 21400 5597 21440
rect 6979 21400 6988 21440
rect 7028 21400 7468 21440
rect 7508 21400 7517 21440
rect 12163 21400 12172 21440
rect 12212 21400 13844 21440
rect 16003 21400 16012 21440
rect 16052 21400 16916 21440
rect 0 21380 80 21400
rect 1219 21399 1277 21400
rect 7555 21356 7613 21357
rect 13804 21356 13844 21400
rect 7470 21316 7564 21356
rect 7604 21316 7613 21356
rect 13795 21316 13804 21356
rect 13844 21316 13853 21356
rect 7555 21315 7613 21316
rect 16876 21272 16916 21400
rect 16972 21356 17012 21484
rect 20995 21483 21053 21484
rect 16963 21316 16972 21356
rect 17012 21316 17021 21356
rect 21424 21272 21504 21292
rect 2500 21232 16052 21272
rect 16876 21232 17164 21272
rect 17204 21232 17213 21272
rect 21187 21232 21196 21272
rect 21236 21232 21504 21272
rect 2500 21104 2540 21232
rect 15811 21188 15869 21189
rect 3679 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 4065 21188
rect 7843 21148 7852 21188
rect 7892 21148 8716 21188
rect 8756 21148 8765 21188
rect 9187 21148 9196 21188
rect 9236 21148 9772 21188
rect 9812 21148 9821 21188
rect 11395 21148 11404 21188
rect 11444 21148 15628 21188
rect 15668 21148 15820 21188
rect 15860 21148 15869 21188
rect 16012 21188 16052 21232
rect 21424 21212 21504 21232
rect 18499 21188 18557 21189
rect 16012 21148 18508 21188
rect 18548 21148 18557 21188
rect 18799 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 19185 21188
rect 15811 21147 15869 21148
rect 18499 21147 18557 21148
rect 20 21064 2540 21104
rect 10339 21064 10348 21104
rect 10388 21064 10924 21104
rect 10964 21064 12076 21104
rect 12116 21064 12125 21104
rect 20 20936 60 21064
rect 14179 21020 14237 21021
rect 19267 21020 19325 21021
rect 2500 20980 14188 21020
rect 14228 20980 14237 21020
rect 17443 20980 17452 21020
rect 17492 20980 19276 21020
rect 19316 20980 19325 21020
rect 2500 20936 2540 20980
rect 14179 20979 14237 20980
rect 19267 20979 19325 20980
rect 20 20896 212 20936
rect 1507 20896 1516 20936
rect 1556 20896 2540 20936
rect 4099 20936 4157 20937
rect 21424 20936 21504 20956
rect 4099 20896 4108 20936
rect 4148 20896 8332 20936
rect 8372 20896 8524 20936
rect 8564 20896 8573 20936
rect 11011 20896 11020 20936
rect 11060 20896 11596 20936
rect 11636 20896 11980 20936
rect 12020 20896 12029 20936
rect 12931 20896 12940 20936
rect 12980 20896 13324 20936
rect 13364 20896 13373 20936
rect 15331 20896 15340 20936
rect 15380 20896 19468 20936
rect 19508 20896 19517 20936
rect 21091 20896 21100 20936
rect 21140 20896 21504 20936
rect 0 20768 80 20788
rect 172 20768 212 20896
rect 4099 20895 4157 20896
rect 21424 20876 21504 20896
rect 6892 20812 11404 20852
rect 11444 20812 11453 20852
rect 16675 20812 16684 20852
rect 16724 20812 17260 20852
rect 17300 20812 17309 20852
rect 6892 20768 6932 20812
rect 9667 20768 9725 20769
rect 10723 20768 10781 20769
rect 0 20728 212 20768
rect 2179 20728 2188 20768
rect 2228 20728 6932 20768
rect 9571 20728 9580 20768
rect 9620 20728 9676 20768
rect 9716 20728 9725 20768
rect 10638 20728 10732 20768
rect 10772 20728 10781 20768
rect 0 20708 80 20728
rect 9667 20727 9725 20728
rect 10723 20727 10781 20728
rect 11299 20768 11357 20769
rect 11299 20728 11308 20768
rect 11348 20728 11753 20768
rect 11793 20728 11802 20768
rect 13123 20728 13132 20768
rect 13172 20728 13420 20768
rect 13460 20728 17492 20768
rect 18014 20728 18023 20768
rect 18063 20728 19180 20768
rect 19220 20728 19229 20768
rect 11299 20727 11357 20728
rect 9676 20684 9716 20727
rect 4675 20644 4684 20684
rect 4724 20644 6412 20684
rect 6452 20644 6461 20684
rect 9676 20644 14476 20684
rect 14516 20644 14525 20684
rect 9955 20600 10013 20601
rect 17452 20600 17492 20728
rect 21424 20600 21504 20620
rect 2851 20560 2860 20600
rect 2900 20560 5452 20600
rect 5492 20560 8620 20600
rect 8660 20560 8669 20600
rect 9571 20560 9580 20600
rect 9620 20560 9964 20600
rect 10004 20560 10013 20600
rect 15139 20560 15148 20600
rect 15188 20560 16204 20600
rect 16244 20560 16253 20600
rect 16867 20560 16876 20600
rect 16916 20560 17356 20600
rect 17396 20560 17405 20600
rect 17452 20560 17548 20600
rect 17588 20560 18604 20600
rect 18644 20560 18653 20600
rect 21283 20560 21292 20600
rect 21332 20560 21504 20600
rect 9955 20559 10013 20560
rect 21424 20540 21504 20560
rect 2563 20516 2621 20517
rect 2563 20476 2572 20516
rect 2612 20476 2706 20516
rect 15331 20476 15340 20516
rect 15380 20476 15628 20516
rect 15668 20476 15677 20516
rect 2563 20475 2621 20476
rect 4099 20432 4157 20433
rect 16291 20432 16349 20433
rect 4014 20392 4108 20432
rect 4148 20392 4157 20432
rect 4919 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 5305 20432
rect 8611 20392 8620 20432
rect 8660 20392 8840 20432
rect 13123 20392 13132 20432
rect 13172 20392 13804 20432
rect 13844 20392 13853 20432
rect 16291 20392 16300 20432
rect 16340 20392 18796 20432
rect 18836 20392 18845 20432
rect 20039 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20425 20432
rect 4099 20391 4157 20392
rect 1699 20308 1708 20348
rect 1748 20308 5452 20348
rect 5492 20308 5501 20348
rect 6019 20264 6077 20265
rect 8800 20264 8840 20392
rect 16291 20391 16349 20392
rect 17251 20348 17309 20349
rect 11203 20308 11212 20348
rect 11252 20308 11500 20348
rect 11540 20308 11549 20348
rect 11971 20308 11980 20348
rect 12020 20308 12364 20348
rect 12404 20308 12413 20348
rect 16195 20308 16204 20348
rect 16244 20308 17260 20348
rect 17300 20308 17309 20348
rect 17251 20307 17309 20308
rect 19555 20348 19613 20349
rect 19555 20308 19564 20348
rect 19604 20308 19948 20348
rect 19988 20308 19997 20348
rect 19555 20307 19613 20308
rect 13027 20264 13085 20265
rect 2668 20224 4300 20264
rect 4340 20224 4349 20264
rect 6019 20224 6028 20264
rect 6068 20224 6124 20264
rect 6164 20224 6173 20264
rect 7939 20224 7948 20264
rect 7988 20224 8524 20264
rect 8564 20224 8573 20264
rect 8800 20224 11788 20264
rect 11828 20224 11837 20264
rect 12942 20224 13036 20264
rect 13076 20224 13085 20264
rect 2668 20180 2708 20224
rect 6019 20223 6077 20224
rect 13027 20223 13085 20224
rect 17059 20264 17117 20265
rect 19267 20264 19325 20265
rect 21424 20264 21504 20284
rect 17059 20224 17068 20264
rect 17108 20224 17300 20264
rect 17059 20223 17117 20224
rect 17260 20181 17300 20224
rect 19267 20224 19276 20264
rect 19316 20224 21504 20264
rect 19267 20223 19325 20224
rect 21424 20204 21504 20224
rect 10435 20180 10493 20181
rect 17251 20180 17309 20181
rect 2659 20140 2668 20180
rect 2708 20140 2717 20180
rect 3043 20140 3052 20180
rect 3092 20140 4684 20180
rect 4724 20140 7372 20180
rect 7412 20140 7421 20180
rect 10435 20140 10444 20180
rect 10484 20140 10676 20180
rect 10980 20140 11020 20180
rect 11060 20140 11069 20180
rect 17251 20140 17260 20180
rect 17300 20140 17309 20180
rect 18468 20140 18508 20180
rect 18548 20140 18557 20180
rect 21091 20140 21100 20180
rect 21140 20140 21149 20180
rect 10435 20139 10493 20140
rect 0 20096 80 20116
rect 2083 20096 2141 20097
rect 9667 20096 9725 20097
rect 10636 20096 10676 20140
rect 11020 20096 11060 20140
rect 17251 20139 17309 20140
rect 16579 20096 16637 20097
rect 18508 20096 18548 20140
rect 21100 20096 21140 20140
rect 0 20056 268 20096
rect 308 20056 317 20096
rect 1411 20056 1420 20096
rect 1460 20056 2092 20096
rect 2132 20056 2141 20096
rect 8035 20056 8044 20096
rect 8084 20056 9100 20096
rect 9140 20056 9149 20096
rect 9582 20056 9676 20096
rect 9716 20056 10540 20096
rect 10580 20056 10589 20096
rect 10636 20056 10924 20096
rect 10964 20056 10973 20096
rect 11020 20056 11404 20096
rect 11444 20056 11453 20096
rect 12835 20056 12844 20096
rect 12884 20056 13228 20096
rect 13268 20056 13748 20096
rect 0 20036 80 20056
rect 2083 20055 2141 20056
rect 8620 20012 8660 20056
rect 9667 20055 9725 20056
rect 10819 20012 10877 20013
rect 11299 20012 11357 20013
rect 13708 20012 13748 20056
rect 16579 20056 16588 20096
rect 16628 20056 17452 20096
rect 17492 20056 17501 20096
rect 18508 20056 20044 20096
rect 20084 20056 20093 20096
rect 21100 20056 21388 20096
rect 21428 20056 21437 20096
rect 16579 20055 16637 20056
rect 8323 19972 8332 20012
rect 8372 19972 8381 20012
rect 8620 19972 8668 20012
rect 8708 19972 8717 20012
rect 10627 19972 10636 20012
rect 10676 19972 10828 20012
rect 10868 19972 10877 20012
rect 11107 19972 11116 20012
rect 11156 19972 11308 20012
rect 11348 19972 11357 20012
rect 13699 19972 13708 20012
rect 13748 19972 13757 20012
rect 16963 19972 16972 20012
rect 17012 19972 18220 20012
rect 18260 19972 18269 20012
rect 8332 19928 8372 19972
rect 10819 19971 10877 19972
rect 11299 19971 11357 19972
rect 16387 19928 16445 19929
rect 21424 19928 21504 19948
rect 4291 19888 4300 19928
rect 4340 19888 4492 19928
rect 4532 19888 4541 19928
rect 5059 19888 5068 19928
rect 5108 19888 5740 19928
rect 5780 19888 5789 19928
rect 8131 19888 8140 19928
rect 8180 19888 8372 19928
rect 8563 19888 8572 19928
rect 8612 19888 9388 19928
rect 9428 19888 9437 19928
rect 10723 19888 10732 19928
rect 10772 19888 11500 19928
rect 11540 19888 11549 19928
rect 13507 19888 13516 19928
rect 13556 19888 16396 19928
rect 16436 19888 16445 19928
rect 17251 19888 17260 19928
rect 17300 19888 18412 19928
rect 18452 19888 19852 19928
rect 19892 19888 19901 19928
rect 20899 19888 20908 19928
rect 20948 19888 21504 19928
rect 16387 19887 16445 19888
rect 21424 19868 21504 19888
rect 16291 19844 16349 19845
rect 19939 19844 19997 19845
rect 3523 19804 3532 19844
rect 3572 19804 4012 19844
rect 4052 19804 5644 19844
rect 5684 19804 5693 19844
rect 10531 19804 10540 19844
rect 10580 19804 16300 19844
rect 16340 19804 16349 19844
rect 19651 19804 19660 19844
rect 19700 19804 19948 19844
rect 19988 19804 19997 19844
rect 16291 19803 16349 19804
rect 19939 19803 19997 19804
rect 1699 19720 1708 19760
rect 1748 19720 6412 19760
rect 6452 19720 8812 19760
rect 8852 19720 8861 19760
rect 9676 19720 10252 19760
rect 10292 19720 10301 19760
rect 12835 19720 12844 19760
rect 12884 19720 13036 19760
rect 13076 19720 17068 19760
rect 17108 19720 17117 19760
rect 17260 19720 18124 19760
rect 18164 19720 19948 19760
rect 19988 19720 19997 19760
rect 9676 19676 9716 19720
rect 10339 19676 10397 19677
rect 16579 19676 16637 19677
rect 17260 19676 17300 19720
rect 3679 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 4065 19676
rect 6115 19636 6124 19676
rect 6164 19636 8908 19676
rect 8948 19636 9676 19676
rect 9716 19636 9725 19676
rect 10254 19636 10348 19676
rect 10388 19636 10397 19676
rect 10723 19636 10732 19676
rect 10772 19636 12692 19676
rect 15907 19636 15916 19676
rect 15956 19636 16588 19676
rect 16628 19636 16637 19676
rect 17251 19636 17260 19676
rect 17300 19636 17309 19676
rect 18799 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 19185 19676
rect 10339 19635 10397 19636
rect 12652 19592 12692 19636
rect 16579 19635 16637 19636
rect 21424 19592 21504 19612
rect 451 19552 460 19592
rect 500 19552 9292 19592
rect 9332 19552 9341 19592
rect 10435 19552 10444 19592
rect 10484 19552 11212 19592
rect 11252 19552 11261 19592
rect 12652 19552 17932 19592
rect 17972 19552 17981 19592
rect 20803 19552 20812 19592
rect 20852 19552 21504 19592
rect 6019 19508 6077 19509
rect 9292 19508 9332 19552
rect 21424 19532 21504 19552
rect 20803 19508 20861 19509
rect 6019 19468 6028 19508
rect 6068 19468 6220 19508
rect 6260 19468 6269 19508
rect 9292 19468 11596 19508
rect 11636 19468 11645 19508
rect 14179 19468 14188 19508
rect 14228 19468 14860 19508
rect 14900 19468 14909 19508
rect 18115 19468 18124 19508
rect 18164 19468 20812 19508
rect 20852 19468 20861 19508
rect 6019 19467 6077 19468
rect 20803 19467 20861 19468
rect 0 19424 80 19444
rect 11203 19424 11261 19425
rect 0 19384 11212 19424
rect 11252 19384 11261 19424
rect 11683 19384 11692 19424
rect 11732 19384 12364 19424
rect 12404 19384 12413 19424
rect 13219 19384 13228 19424
rect 13268 19384 15340 19424
rect 15380 19384 15389 19424
rect 17827 19384 17836 19424
rect 17876 19384 17885 19424
rect 0 19364 80 19384
rect 11203 19383 11261 19384
rect 2563 19340 2621 19341
rect 17836 19340 17876 19384
rect 2563 19300 2572 19340
rect 2612 19300 2706 19340
rect 4291 19300 4300 19340
rect 4340 19300 6028 19340
rect 6068 19300 6077 19340
rect 6691 19300 6700 19340
rect 6740 19300 8044 19340
rect 8084 19300 9908 19340
rect 9955 19300 9964 19340
rect 10004 19300 10060 19340
rect 10100 19300 12844 19340
rect 12884 19300 12893 19340
rect 13699 19300 13708 19340
rect 13748 19300 14092 19340
rect 14132 19300 14141 19340
rect 14755 19300 14764 19340
rect 14804 19300 19948 19340
rect 19988 19300 19997 19340
rect 2563 19299 2621 19300
rect 7555 19256 7613 19257
rect 4771 19216 4780 19256
rect 4820 19216 7564 19256
rect 7604 19216 7613 19256
rect 9868 19256 9908 19300
rect 10435 19256 10493 19257
rect 21424 19256 21504 19276
rect 9868 19216 10444 19256
rect 10484 19216 12556 19256
rect 12596 19216 12605 19256
rect 15811 19216 15820 19256
rect 15860 19216 16204 19256
rect 16244 19216 16253 19256
rect 17539 19216 17548 19256
rect 17588 19216 21504 19256
rect 7555 19215 7613 19216
rect 10435 19215 10493 19216
rect 21424 19196 21504 19216
rect 5443 19172 5501 19173
rect 7459 19172 7517 19173
rect 2500 19132 5452 19172
rect 5492 19132 6796 19172
rect 6836 19132 7468 19172
rect 7508 19132 7517 19172
rect 9091 19132 9100 19172
rect 9140 19132 14188 19172
rect 14228 19132 14237 19172
rect 17059 19132 17068 19172
rect 17108 19132 18604 19172
rect 18644 19132 18653 19172
rect 19267 19132 19276 19172
rect 19316 19132 19660 19172
rect 19700 19132 19709 19172
rect 2500 19088 2540 19132
rect 5443 19131 5501 19132
rect 7459 19131 7517 19132
rect 1315 19048 1324 19088
rect 1364 19048 2540 19088
rect 6019 19048 6028 19088
rect 6068 19048 7276 19088
rect 7316 19048 7325 19088
rect 7555 19048 7564 19088
rect 7604 19048 8332 19088
rect 8372 19048 8381 19088
rect 12643 19048 12652 19088
rect 12692 19048 12940 19088
rect 12980 19048 12989 19088
rect 13603 19048 13612 19088
rect 13652 19048 14380 19088
rect 14420 19048 14429 19088
rect 17635 19048 17644 19088
rect 17684 19048 17836 19088
rect 17876 19048 17885 19088
rect 9667 18964 9676 19004
rect 9716 18964 13364 19004
rect 13324 18920 13364 18964
rect 14467 18920 14525 18921
rect 15907 18920 15965 18921
rect 16291 18920 16349 18921
rect 21091 18920 21149 18921
rect 21424 18920 21504 18940
rect 4919 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 5305 18920
rect 9475 18880 9484 18920
rect 9524 18880 9964 18920
rect 10004 18880 10013 18920
rect 11203 18880 11212 18920
rect 11252 18880 12268 18920
rect 12308 18880 12317 18920
rect 13315 18880 13324 18920
rect 13364 18880 13804 18920
rect 13844 18880 13853 18920
rect 14467 18880 14476 18920
rect 14516 18880 14668 18920
rect 14708 18880 14717 18920
rect 15907 18880 15916 18920
rect 15956 18880 16300 18920
rect 16340 18880 16349 18920
rect 20039 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20425 18920
rect 21091 18880 21100 18920
rect 21140 18880 21504 18920
rect 14467 18879 14525 18880
rect 15907 18879 15965 18880
rect 16291 18879 16349 18880
rect 21091 18879 21149 18880
rect 21424 18860 21504 18880
rect 12259 18836 12317 18837
rect 12259 18796 12268 18836
rect 12308 18796 20084 18836
rect 12259 18795 12317 18796
rect 0 18752 80 18772
rect 1219 18752 1277 18753
rect 11107 18752 11165 18753
rect 20044 18752 20084 18796
rect 20515 18752 20573 18753
rect 0 18712 1228 18752
rect 1268 18712 1277 18752
rect 0 18692 80 18712
rect 1219 18711 1277 18712
rect 4108 18712 6220 18752
rect 6260 18712 6269 18752
rect 6691 18712 6700 18752
rect 6740 18712 7564 18752
rect 7604 18712 7613 18752
rect 11107 18712 11116 18752
rect 11156 18712 11212 18752
rect 11252 18712 11261 18752
rect 14659 18712 14668 18752
rect 14708 18712 14956 18752
rect 14996 18712 15005 18752
rect 20035 18712 20044 18752
rect 20084 18712 20093 18752
rect 20227 18712 20236 18752
rect 20276 18712 20524 18752
rect 20564 18712 20573 18752
rect 4108 18668 4148 18712
rect 11107 18711 11165 18712
rect 20515 18711 20573 18712
rect 20995 18752 21053 18753
rect 20995 18712 21004 18752
rect 21044 18712 21053 18752
rect 20995 18711 21053 18712
rect 14083 18668 14141 18669
rect 21004 18668 21044 18711
rect 2467 18628 2476 18668
rect 2516 18628 4108 18668
rect 4148 18628 4157 18668
rect 5059 18628 5068 18668
rect 5108 18628 5644 18668
rect 5684 18628 5836 18668
rect 5876 18628 5885 18668
rect 7939 18628 7948 18668
rect 7988 18628 8620 18668
rect 8660 18628 8669 18668
rect 9772 18628 14092 18668
rect 14132 18628 15052 18668
rect 15092 18628 15101 18668
rect 16195 18628 16204 18668
rect 16244 18628 16684 18668
rect 16724 18628 16733 18668
rect 19075 18628 19084 18668
rect 19124 18628 19756 18668
rect 19796 18628 19805 18668
rect 20524 18628 21044 18668
rect 3715 18584 3773 18585
rect 6403 18584 6461 18585
rect 3331 18544 3340 18584
rect 3380 18544 3724 18584
rect 3764 18544 3773 18584
rect 4195 18544 4204 18584
rect 4244 18544 4972 18584
rect 5012 18544 5021 18584
rect 6318 18544 6412 18584
rect 6452 18544 6461 18584
rect 3715 18543 3773 18544
rect 6403 18543 6461 18544
rect 6595 18584 6653 18585
rect 8035 18584 8093 18585
rect 6595 18544 6604 18584
rect 6644 18544 6796 18584
rect 6836 18544 6845 18584
rect 6979 18544 6988 18584
rect 7028 18544 8044 18584
rect 8084 18544 8716 18584
rect 8756 18544 8765 18584
rect 6595 18543 6653 18544
rect 8035 18543 8093 18544
rect 7939 18500 7997 18501
rect 9772 18500 9812 18628
rect 14083 18627 14141 18628
rect 20524 18585 20564 18628
rect 13699 18584 13757 18585
rect 20515 18584 20573 18585
rect 10147 18544 10156 18584
rect 10196 18544 10348 18584
rect 10388 18544 10540 18584
rect 10580 18544 10924 18584
rect 10964 18544 10973 18584
rect 13219 18544 13228 18584
rect 13268 18544 13708 18584
rect 13748 18544 15916 18584
rect 15956 18544 15965 18584
rect 20515 18544 20524 18584
rect 20564 18544 20573 18584
rect 13699 18543 13757 18544
rect 20515 18543 20573 18544
rect 20995 18584 21053 18585
rect 21424 18584 21504 18604
rect 20995 18544 21004 18584
rect 21044 18544 21504 18584
rect 20995 18543 21053 18544
rect 21424 18524 21504 18544
rect 2083 18460 2092 18500
rect 2132 18460 5356 18500
rect 5396 18460 5932 18500
rect 5972 18460 5981 18500
rect 7939 18460 7948 18500
rect 7988 18460 9812 18500
rect 9859 18460 9868 18500
rect 9908 18460 16972 18500
rect 17012 18460 17021 18500
rect 7939 18459 7997 18460
rect 2563 18416 2621 18417
rect 10339 18416 10397 18417
rect 17059 18416 17117 18417
rect 2563 18376 2572 18416
rect 2612 18376 4204 18416
rect 4244 18376 4253 18416
rect 5635 18376 5644 18416
rect 5684 18376 7660 18416
rect 7700 18376 7948 18416
rect 7988 18376 7997 18416
rect 9763 18376 9772 18416
rect 9812 18376 10348 18416
rect 10388 18376 10636 18416
rect 10676 18376 10685 18416
rect 12547 18376 12556 18416
rect 12596 18376 14572 18416
rect 14612 18376 15052 18416
rect 15092 18376 15101 18416
rect 17059 18376 17068 18416
rect 17108 18376 17164 18416
rect 17204 18376 19180 18416
rect 19220 18376 19852 18416
rect 19892 18376 19901 18416
rect 2563 18375 2621 18376
rect 10339 18375 10397 18376
rect 17059 18375 17117 18376
rect 14467 18332 14525 18333
rect 20515 18332 20573 18333
rect 1123 18292 1132 18332
rect 1172 18292 1612 18332
rect 1652 18292 1661 18332
rect 1795 18292 1804 18332
rect 1844 18292 6412 18332
rect 6452 18292 6461 18332
rect 12835 18292 12844 18332
rect 12884 18292 13900 18332
rect 13940 18292 13949 18332
rect 14382 18292 14476 18332
rect 14516 18292 14525 18332
rect 16003 18292 16012 18332
rect 16052 18292 20524 18332
rect 20564 18292 20573 18332
rect 14467 18291 14525 18292
rect 20515 18291 20573 18292
rect 15139 18248 15197 18249
rect 21424 18248 21504 18268
rect 3436 18208 7852 18248
rect 7892 18208 7901 18248
rect 8800 18208 13228 18248
rect 13268 18208 13277 18248
rect 14371 18208 14380 18248
rect 14420 18208 15148 18248
rect 15188 18208 15197 18248
rect 16771 18208 16780 18248
rect 16820 18208 21504 18248
rect 3235 18164 3293 18165
rect 3043 18124 3052 18164
rect 3092 18124 3244 18164
rect 3284 18124 3293 18164
rect 3235 18123 3293 18124
rect 0 18080 80 18100
rect 1219 18080 1277 18081
rect 0 18040 1228 18080
rect 1268 18040 1277 18080
rect 0 18020 80 18040
rect 1219 18039 1277 18040
rect 1507 18080 1565 18081
rect 3436 18080 3476 18208
rect 8800 18164 8840 18208
rect 15139 18207 15197 18208
rect 21424 18188 21504 18208
rect 16387 18164 16445 18165
rect 3679 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 4065 18164
rect 5443 18124 5452 18164
rect 5492 18124 5836 18164
rect 5876 18124 5885 18164
rect 6211 18124 6220 18164
rect 6260 18124 6604 18164
rect 6644 18124 6653 18164
rect 8419 18124 8428 18164
rect 8468 18124 8840 18164
rect 9187 18124 9196 18164
rect 9236 18124 10156 18164
rect 10196 18124 15436 18164
rect 15476 18124 15485 18164
rect 16387 18124 16396 18164
rect 16436 18124 17260 18164
rect 17300 18124 17309 18164
rect 18799 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 19185 18164
rect 16387 18123 16445 18124
rect 13699 18080 13757 18081
rect 19459 18080 19517 18081
rect 1507 18040 1516 18080
rect 1556 18040 3436 18080
rect 3476 18040 3485 18080
rect 5548 18040 13556 18080
rect 13614 18040 13708 18080
rect 13748 18040 13757 18080
rect 1507 18039 1565 18040
rect 1507 17956 1516 17996
rect 1556 17956 2188 17996
rect 2228 17956 2237 17996
rect 2467 17956 2476 17996
rect 2516 17956 3340 17996
rect 3380 17956 4396 17996
rect 4436 17956 4445 17996
rect 67 17912 125 17913
rect 5548 17912 5588 18040
rect 6403 17996 6461 17997
rect 6318 17956 6412 17996
rect 6452 17956 6461 17996
rect 6403 17955 6461 17956
rect 8227 17996 8285 17997
rect 13516 17996 13556 18040
rect 13699 18039 13757 18040
rect 15532 18040 18220 18080
rect 18260 18040 19468 18080
rect 19508 18040 19948 18080
rect 19988 18040 19997 18080
rect 15532 17996 15572 18040
rect 19459 18039 19517 18040
rect 17443 17996 17501 17997
rect 8227 17956 8236 17996
rect 8276 17956 9196 17996
rect 9236 17956 9245 17996
rect 13516 17956 15572 17996
rect 15619 17956 15628 17996
rect 15668 17956 15916 17996
rect 15956 17956 15965 17996
rect 17155 17956 17164 17996
rect 17204 17956 17452 17996
rect 17492 17956 17501 17996
rect 18787 17956 18796 17996
rect 18836 17956 19468 17996
rect 19508 17956 19517 17996
rect 8227 17955 8285 17956
rect 17443 17955 17501 17956
rect 15331 17912 15389 17913
rect 16483 17912 16541 17913
rect 21424 17912 21504 17932
rect 67 17872 76 17912
rect 116 17872 2860 17912
rect 2900 17872 5588 17912
rect 5827 17872 5836 17912
rect 5876 17872 6452 17912
rect 7747 17872 7756 17912
rect 7796 17872 8140 17912
rect 8180 17872 8524 17912
rect 8564 17872 8573 17912
rect 9475 17872 9484 17912
rect 9524 17872 10828 17912
rect 10868 17872 10877 17912
rect 12835 17872 12844 17912
rect 12884 17872 13516 17912
rect 13556 17872 13565 17912
rect 15331 17872 15340 17912
rect 15380 17872 16012 17912
rect 16052 17872 16061 17912
rect 16483 17872 16492 17912
rect 16532 17872 17260 17912
rect 17300 17872 17309 17912
rect 17443 17872 17452 17912
rect 17492 17872 21504 17912
rect 67 17871 125 17872
rect 2563 17828 2621 17829
rect 2755 17828 2813 17829
rect 6412 17828 6452 17872
rect 15331 17871 15389 17872
rect 16483 17871 16541 17872
rect 21424 17852 21504 17872
rect 9571 17828 9629 17829
rect 17251 17828 17309 17829
rect 2179 17788 2188 17828
rect 2228 17788 2572 17828
rect 2612 17788 2621 17828
rect 2669 17788 2764 17828
rect 2804 17788 2956 17828
rect 2996 17788 3005 17828
rect 5155 17788 5164 17828
rect 5204 17788 5452 17828
rect 5492 17788 6316 17828
rect 6356 17788 6365 17828
rect 6412 17788 9580 17828
rect 9620 17788 9629 17828
rect 2563 17787 2621 17788
rect 2755 17787 2813 17788
rect 9571 17787 9629 17788
rect 9676 17788 11020 17828
rect 11060 17788 11069 17828
rect 13132 17788 16588 17828
rect 16628 17788 16637 17828
rect 17251 17788 17260 17828
rect 17300 17788 17356 17828
rect 17396 17788 17405 17828
rect 1891 17746 1900 17786
rect 1940 17746 2132 17786
rect 2092 17744 2132 17746
rect 5059 17744 5117 17745
rect 6403 17744 6461 17745
rect 9676 17744 9716 17788
rect 2092 17704 4876 17744
rect 4916 17704 4925 17744
rect 5059 17704 5068 17744
rect 5108 17704 5202 17744
rect 5347 17704 5356 17744
rect 5396 17704 6412 17744
rect 6452 17704 6461 17744
rect 6883 17704 6892 17744
rect 6932 17704 7084 17744
rect 7124 17704 7133 17744
rect 9379 17704 9388 17744
rect 9428 17704 9676 17744
rect 9716 17704 9725 17744
rect 9955 17704 9964 17744
rect 10004 17704 10924 17744
rect 10964 17704 10973 17744
rect 5059 17703 5117 17704
rect 6403 17703 6461 17704
rect 7651 17660 7709 17661
rect 11779 17660 11837 17661
rect 1804 17620 2476 17660
rect 2516 17620 2525 17660
rect 3052 17620 3820 17660
rect 3860 17620 3869 17660
rect 5539 17620 5548 17660
rect 5588 17620 7660 17660
rect 7700 17620 8428 17660
rect 8468 17620 8477 17660
rect 8995 17620 9004 17660
rect 9044 17620 9053 17660
rect 9283 17620 9292 17660
rect 9332 17620 10636 17660
rect 10676 17620 10685 17660
rect 11683 17620 11692 17660
rect 11732 17620 11788 17660
rect 11828 17620 11837 17660
rect 0 17408 80 17428
rect 1804 17408 1844 17620
rect 3052 17576 3092 17620
rect 7651 17619 7709 17620
rect 7171 17576 7229 17577
rect 9004 17576 9044 17620
rect 11779 17619 11837 17620
rect 13132 17576 13172 17788
rect 17251 17787 17309 17788
rect 13228 17704 13900 17744
rect 13940 17704 13949 17744
rect 15235 17704 15244 17744
rect 15284 17704 18892 17744
rect 18932 17704 18941 17744
rect 19267 17704 19276 17744
rect 19316 17704 20044 17744
rect 20084 17704 20093 17744
rect 13228 17660 13268 17704
rect 13219 17620 13228 17660
rect 13268 17620 13277 17660
rect 18019 17620 18028 17660
rect 18068 17620 19948 17660
rect 19988 17620 19997 17660
rect 21424 17576 21504 17596
rect 3043 17536 3052 17576
rect 3092 17536 3101 17576
rect 3427 17536 3436 17576
rect 3476 17536 4684 17576
rect 4724 17536 4733 17576
rect 6019 17536 6028 17576
rect 6068 17536 6604 17576
rect 6644 17536 6653 17576
rect 7086 17536 7180 17576
rect 7220 17536 7229 17576
rect 7555 17536 7564 17576
rect 7604 17536 8044 17576
rect 8084 17536 8093 17576
rect 9004 17536 12404 17576
rect 13123 17536 13132 17576
rect 13172 17536 13181 17576
rect 17827 17536 17836 17576
rect 17876 17536 21504 17576
rect 7171 17535 7229 17536
rect 7939 17492 7997 17493
rect 2500 17452 7948 17492
rect 7988 17452 7997 17492
rect 2500 17408 2540 17452
rect 7939 17451 7997 17452
rect 10819 17492 10877 17493
rect 12364 17492 12404 17536
rect 21424 17516 21504 17536
rect 10819 17452 10828 17492
rect 10868 17452 10924 17492
rect 10964 17452 10973 17492
rect 12364 17452 16972 17492
rect 17012 17452 17021 17492
rect 19171 17452 19180 17492
rect 19220 17452 19660 17492
rect 19700 17452 19709 17492
rect 10819 17451 10877 17452
rect 4195 17408 4253 17409
rect 4771 17408 4829 17409
rect 8707 17408 8765 17409
rect 0 17368 172 17408
rect 212 17368 221 17408
rect 1795 17368 1804 17408
rect 1844 17368 1853 17408
rect 2179 17368 2188 17408
rect 2228 17368 2540 17408
rect 2947 17368 2956 17408
rect 2996 17368 4204 17408
rect 4244 17368 4780 17408
rect 4820 17368 4829 17408
rect 4919 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 5305 17408
rect 7459 17368 7468 17408
rect 7508 17368 8140 17408
rect 8180 17368 8189 17408
rect 8622 17368 8716 17408
rect 8756 17368 8765 17408
rect 0 17348 80 17368
rect 4195 17367 4253 17368
rect 4771 17367 4829 17368
rect 8707 17367 8765 17368
rect 9571 17408 9629 17409
rect 9571 17368 9580 17408
rect 9620 17368 12076 17408
rect 12116 17368 12125 17408
rect 12931 17368 12940 17408
rect 12980 17368 13516 17408
rect 13556 17368 14092 17408
rect 14132 17368 14141 17408
rect 14188 17368 18412 17408
rect 18452 17368 18461 17408
rect 20039 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20425 17408
rect 9571 17367 9629 17368
rect 2563 17324 2621 17325
rect 6403 17324 6461 17325
rect 7363 17324 7421 17325
rect 14188 17324 14228 17368
rect 20611 17324 20669 17325
rect 2563 17284 2572 17324
rect 2612 17284 4108 17324
rect 4148 17284 4300 17324
rect 4340 17284 4349 17324
rect 6403 17284 6412 17324
rect 6452 17284 7372 17324
rect 7412 17284 8852 17324
rect 2563 17283 2621 17284
rect 6403 17283 6461 17284
rect 7363 17283 7421 17284
rect 8812 17240 8852 17284
rect 8908 17284 14228 17324
rect 17155 17284 17164 17324
rect 17204 17284 17548 17324
rect 17588 17284 17597 17324
rect 19843 17284 19852 17324
rect 19892 17284 20620 17324
rect 20660 17284 20669 17324
rect 8908 17240 8948 17284
rect 20611 17283 20669 17284
rect 9859 17240 9917 17241
rect 13699 17240 13757 17241
rect 21424 17240 21504 17260
rect 1315 17200 1324 17240
rect 1364 17200 2092 17240
rect 2132 17200 2141 17240
rect 2476 17200 2668 17240
rect 2708 17200 2717 17240
rect 3907 17200 3916 17240
rect 3956 17200 4204 17240
rect 4244 17200 4253 17240
rect 8812 17200 8948 17240
rect 8995 17200 9004 17240
rect 9044 17200 9868 17240
rect 9908 17200 9917 17240
rect 11875 17200 11884 17240
rect 11924 17200 12460 17240
rect 12500 17200 12509 17240
rect 13614 17200 13708 17240
rect 13748 17200 13757 17240
rect 14083 17200 14092 17240
rect 14132 17200 14668 17240
rect 14708 17200 14717 17240
rect 16387 17200 16396 17240
rect 16436 17200 21504 17240
rect 2476 17072 2516 17200
rect 9859 17199 9917 17200
rect 13699 17199 13757 17200
rect 21424 17180 21504 17200
rect 2563 17156 2621 17157
rect 7555 17156 7613 17157
rect 13219 17156 13277 17157
rect 2563 17116 2572 17156
rect 2612 17116 2621 17156
rect 2563 17115 2621 17116
rect 2668 17116 3239 17156
rect 3279 17116 4588 17156
rect 4628 17116 4637 17156
rect 7555 17116 7564 17156
rect 7604 17116 9524 17156
rect 13123 17116 13132 17156
rect 13172 17116 13228 17156
rect 13268 17116 13804 17156
rect 13844 17116 13853 17156
rect 14755 17116 14764 17156
rect 14804 17116 19276 17156
rect 19316 17116 19325 17156
rect 2572 17072 2612 17115
rect 2668 17072 2708 17116
rect 7555 17115 7613 17116
rect 6211 17072 6269 17073
rect 7171 17072 7229 17073
rect 9484 17072 9524 17116
rect 13219 17115 13277 17116
rect 16675 17072 16733 17073
rect 2467 17032 2476 17072
rect 2516 17032 2612 17072
rect 2659 17032 2668 17072
rect 2708 17032 2717 17072
rect 3715 17032 3724 17072
rect 3764 17032 4492 17072
rect 4532 17032 4541 17072
rect 6211 17032 6220 17072
rect 6260 17032 7180 17072
rect 7220 17032 7660 17072
rect 7700 17032 7709 17072
rect 9475 17032 9484 17072
rect 9524 17032 9533 17072
rect 9667 17032 9676 17072
rect 9716 17032 9868 17072
rect 9908 17032 9917 17072
rect 12067 17032 12076 17072
rect 12116 17032 15148 17072
rect 15188 17032 15820 17072
rect 15860 17032 15869 17072
rect 16675 17032 16684 17072
rect 16724 17032 17644 17072
rect 17684 17032 17693 17072
rect 6211 17031 6269 17032
rect 7171 17031 7229 17032
rect 16675 17031 16733 17032
rect 19651 16988 19709 16989
rect 2500 16948 13516 16988
rect 13556 16948 13565 16988
rect 15043 16948 15052 16988
rect 15092 16948 16396 16988
rect 16436 16948 18700 16988
rect 18740 16948 18749 16988
rect 19566 16948 19660 16988
rect 19700 16948 19709 16988
rect 0 16736 80 16756
rect 931 16736 989 16737
rect 0 16696 940 16736
rect 980 16696 989 16736
rect 0 16676 80 16696
rect 931 16695 989 16696
rect 2500 16568 2540 16948
rect 19651 16947 19709 16948
rect 21424 16904 21504 16924
rect 2851 16864 2860 16904
rect 2900 16864 3244 16904
rect 3284 16864 3293 16904
rect 3427 16864 3436 16904
rect 3476 16864 4012 16904
rect 4052 16864 4061 16904
rect 4108 16864 21504 16904
rect 3235 16736 3293 16737
rect 3235 16696 3244 16736
rect 3284 16696 3340 16736
rect 3380 16696 3389 16736
rect 3235 16695 3293 16696
rect 3679 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 4065 16652
rect 355 16528 364 16568
rect 404 16528 2540 16568
rect 4108 16484 4148 16864
rect 21424 16844 21504 16864
rect 15715 16820 15773 16821
rect 4195 16780 4204 16820
rect 4244 16780 7852 16820
rect 7892 16780 7901 16820
rect 8131 16780 8140 16820
rect 8180 16780 15724 16820
rect 15764 16780 15773 16820
rect 15715 16779 15773 16780
rect 18499 16820 18557 16821
rect 18499 16780 18508 16820
rect 18548 16780 18604 16820
rect 18644 16780 18892 16820
rect 18932 16780 18941 16820
rect 18499 16779 18557 16780
rect 7651 16736 7709 16737
rect 11395 16736 11453 16737
rect 6883 16696 6892 16736
rect 6932 16696 7084 16736
rect 7124 16696 7133 16736
rect 7566 16696 7660 16736
rect 7700 16696 7709 16736
rect 10915 16696 10924 16736
rect 10964 16696 11404 16736
rect 11444 16696 11453 16736
rect 7651 16695 7709 16696
rect 11395 16695 11453 16696
rect 13315 16736 13373 16737
rect 18691 16736 18749 16737
rect 13315 16696 13324 16736
rect 13364 16696 13612 16736
rect 13652 16696 14764 16736
rect 14804 16696 14813 16736
rect 15523 16696 15532 16736
rect 15572 16696 15820 16736
rect 15860 16696 15869 16736
rect 18115 16696 18124 16736
rect 18164 16696 18700 16736
rect 18740 16696 18749 16736
rect 13315 16695 13373 16696
rect 18691 16695 18749 16696
rect 13795 16652 13853 16653
rect 4291 16612 4300 16652
rect 4340 16612 5356 16652
rect 5396 16612 11212 16652
rect 11252 16612 11261 16652
rect 13795 16612 13804 16652
rect 13844 16612 16436 16652
rect 18211 16612 18220 16652
rect 18260 16612 18604 16652
rect 18644 16612 18653 16652
rect 18799 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 19185 16652
rect 13795 16611 13853 16612
rect 4195 16568 4253 16569
rect 16291 16568 16349 16569
rect 4195 16528 4204 16568
rect 4244 16528 7564 16568
rect 7604 16528 7613 16568
rect 9475 16528 9484 16568
rect 9524 16528 11308 16568
rect 11348 16528 11357 16568
rect 15331 16528 15340 16568
rect 15380 16528 16300 16568
rect 16340 16528 16349 16568
rect 16396 16568 16436 16612
rect 21424 16568 21504 16588
rect 16396 16528 21504 16568
rect 4195 16527 4253 16528
rect 16291 16527 16349 16528
rect 21424 16508 21504 16528
rect 3619 16444 3628 16484
rect 3668 16444 4148 16484
rect 9571 16444 9580 16484
rect 9620 16444 9772 16484
rect 9812 16444 9821 16484
rect 10051 16444 10060 16484
rect 10100 16444 20044 16484
rect 20084 16444 20093 16484
rect 4867 16400 4925 16401
rect 9379 16400 9437 16401
rect 19267 16400 19325 16401
rect 3523 16360 3532 16400
rect 3572 16360 3916 16400
rect 3956 16360 3965 16400
rect 4195 16360 4204 16400
rect 4244 16360 4588 16400
rect 4628 16360 4637 16400
rect 4782 16360 4876 16400
rect 4916 16360 4925 16400
rect 6979 16360 6988 16400
rect 7028 16360 7276 16400
rect 7316 16360 8908 16400
rect 8948 16360 8957 16400
rect 9379 16360 9388 16400
rect 9428 16360 10732 16400
rect 10772 16360 10781 16400
rect 11203 16360 11212 16400
rect 11252 16360 13708 16400
rect 13748 16360 13757 16400
rect 14659 16360 14668 16400
rect 14708 16360 15052 16400
rect 15092 16360 15101 16400
rect 15427 16360 15436 16400
rect 15476 16360 19276 16400
rect 19316 16360 19325 16400
rect 19459 16360 19468 16400
rect 19508 16360 21236 16400
rect 4867 16359 4925 16360
rect 9379 16359 9437 16360
rect 19267 16359 19325 16360
rect 21091 16316 21149 16317
rect 2500 16276 10964 16316
rect 11107 16276 11116 16316
rect 11156 16276 17260 16316
rect 17300 16276 17309 16316
rect 17635 16276 17644 16316
rect 17684 16276 19180 16316
rect 19220 16276 19229 16316
rect 21006 16276 21100 16316
rect 21140 16276 21149 16316
rect 2500 16232 2540 16276
rect 10924 16232 10964 16276
rect 21091 16275 21149 16276
rect 11011 16232 11069 16233
rect 15907 16232 15965 16233
rect 20995 16232 21053 16233
rect 1699 16192 1708 16232
rect 1748 16192 2284 16232
rect 2324 16192 2540 16232
rect 2755 16192 2764 16232
rect 2804 16192 4108 16232
rect 4148 16192 4157 16232
rect 4579 16192 4588 16232
rect 4628 16192 5452 16232
rect 5492 16192 5501 16232
rect 8323 16192 8332 16232
rect 8372 16192 10828 16232
rect 10868 16192 10877 16232
rect 10924 16192 11020 16232
rect 11060 16192 11596 16232
rect 11636 16192 11645 16232
rect 15619 16192 15628 16232
rect 15668 16192 15916 16232
rect 15956 16192 15965 16232
rect 16579 16192 16588 16232
rect 16628 16192 16876 16232
rect 16916 16192 16925 16232
rect 18787 16192 18796 16232
rect 18836 16192 19084 16232
rect 19124 16192 19133 16232
rect 19363 16192 19372 16232
rect 19412 16192 19756 16232
rect 19796 16192 19805 16232
rect 20910 16192 21004 16232
rect 21044 16192 21053 16232
rect 21196 16232 21236 16360
rect 21424 16232 21504 16252
rect 21196 16192 21504 16232
rect 4588 16148 4628 16192
rect 11011 16191 11069 16192
rect 15907 16191 15965 16192
rect 19372 16148 19412 16192
rect 20995 16191 21053 16192
rect 21424 16172 21504 16192
rect 3715 16108 3724 16148
rect 3764 16108 4628 16148
rect 9091 16108 9100 16148
rect 9140 16108 12940 16148
rect 12980 16108 12989 16148
rect 18691 16108 18700 16148
rect 18740 16108 19412 16148
rect 0 16064 80 16084
rect 4099 16064 4157 16065
rect 13027 16064 13085 16065
rect 0 16024 4108 16064
rect 4148 16024 4157 16064
rect 9571 16024 9580 16064
rect 9620 16024 9868 16064
rect 9908 16024 9917 16064
rect 11779 16024 11788 16064
rect 11828 16024 13036 16064
rect 13076 16024 13085 16064
rect 14659 16024 14668 16064
rect 14708 16024 14956 16064
rect 14996 16024 15005 16064
rect 19267 16024 19276 16064
rect 19316 16024 20044 16064
rect 20084 16024 20093 16064
rect 0 16004 80 16024
rect 4099 16023 4157 16024
rect 13027 16023 13085 16024
rect 1891 15980 1949 15981
rect 4483 15980 4541 15981
rect 18019 15980 18077 15981
rect 1891 15940 1900 15980
rect 1940 15940 1996 15980
rect 2036 15940 2045 15980
rect 3523 15940 3532 15980
rect 3572 15940 4012 15980
rect 4052 15940 4061 15980
rect 4398 15940 4492 15980
rect 4532 15940 18028 15980
rect 18068 15940 18077 15980
rect 18691 15940 18700 15980
rect 18740 15940 18988 15980
rect 19028 15940 19037 15980
rect 19468 15940 21292 15980
rect 21332 15940 21341 15980
rect 1891 15939 1949 15940
rect 4483 15939 4541 15940
rect 18019 15939 18077 15940
rect 19468 15896 19508 15940
rect 21424 15896 21504 15916
rect 4919 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 5305 15896
rect 6019 15856 6028 15896
rect 6068 15856 10156 15896
rect 10196 15856 11212 15896
rect 11252 15856 11261 15896
rect 16675 15856 16684 15896
rect 16724 15856 16972 15896
rect 17012 15856 17021 15896
rect 17923 15856 17932 15896
rect 17972 15856 19276 15896
rect 19316 15856 19325 15896
rect 19459 15856 19468 15896
rect 19508 15856 19517 15896
rect 20039 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20425 15896
rect 21292 15856 21504 15896
rect 20 15772 1612 15812
rect 1652 15772 1661 15812
rect 1891 15772 1900 15812
rect 1940 15772 1949 15812
rect 2851 15772 2860 15812
rect 2900 15772 8236 15812
rect 8276 15772 9580 15812
rect 9620 15772 9629 15812
rect 9763 15772 9772 15812
rect 9812 15772 10060 15812
rect 10100 15772 17644 15812
rect 17684 15772 17693 15812
rect 19843 15772 19852 15812
rect 19892 15772 21196 15812
rect 21236 15772 21245 15812
rect 20 15560 60 15772
rect 1900 15728 1940 15772
rect 16291 15728 16349 15729
rect 16771 15728 16829 15729
rect 21292 15728 21332 15856
rect 21424 15836 21504 15856
rect 1900 15688 1996 15728
rect 2036 15688 2045 15728
rect 2500 15688 14092 15728
rect 14132 15688 14141 15728
rect 16291 15688 16300 15728
rect 16340 15688 16780 15728
rect 16820 15688 16829 15728
rect 16963 15688 16972 15728
rect 17012 15688 17548 15728
rect 17588 15688 18220 15728
rect 18260 15688 18269 15728
rect 20140 15688 21332 15728
rect 1219 15644 1277 15645
rect 2500 15644 2540 15688
rect 16291 15687 16349 15688
rect 16771 15687 16829 15688
rect 20140 15644 20180 15688
rect 1219 15604 1228 15644
rect 1268 15604 2540 15644
rect 5539 15604 5548 15644
rect 5588 15604 8908 15644
rect 8948 15604 8957 15644
rect 13027 15604 13036 15644
rect 13076 15604 20180 15644
rect 1219 15603 1277 15604
rect 1891 15560 1949 15561
rect 20131 15560 20189 15561
rect 21424 15560 21504 15580
rect 20 15520 212 15560
rect 1806 15520 1900 15560
rect 1940 15520 1949 15560
rect 4003 15520 4012 15560
rect 4052 15520 6988 15560
rect 7028 15520 7037 15560
rect 8515 15520 8524 15560
rect 8564 15520 10540 15560
rect 10580 15520 10589 15560
rect 12835 15520 12844 15560
rect 12884 15520 14956 15560
rect 14996 15520 15820 15560
rect 15860 15520 16588 15560
rect 16628 15520 16780 15560
rect 16820 15520 16829 15560
rect 17443 15520 17452 15560
rect 17492 15520 18124 15560
rect 18164 15520 18173 15560
rect 20131 15520 20140 15560
rect 20180 15520 21504 15560
rect 0 15392 80 15412
rect 172 15392 212 15520
rect 1891 15519 1949 15520
rect 20131 15519 20189 15520
rect 21424 15500 21504 15520
rect 931 15436 940 15476
rect 980 15436 5644 15476
rect 5684 15436 5693 15476
rect 5827 15436 5836 15476
rect 5876 15436 7468 15476
rect 7508 15436 11360 15476
rect 16099 15436 16108 15476
rect 16148 15436 19660 15476
rect 19700 15436 19709 15476
rect 11320 15392 11360 15436
rect 16387 15392 16445 15393
rect 18211 15392 18269 15393
rect 0 15352 212 15392
rect 4963 15352 4972 15392
rect 5012 15352 7948 15392
rect 7988 15352 7997 15392
rect 11320 15352 16396 15392
rect 16436 15352 16445 15392
rect 17731 15352 17740 15392
rect 17780 15352 18220 15392
rect 18260 15352 18269 15392
rect 0 15332 80 15352
rect 16387 15351 16445 15352
rect 18211 15351 18269 15352
rect 20140 15352 21388 15392
rect 21428 15352 21437 15392
rect 16483 15308 16541 15309
rect 20140 15308 20180 15352
rect 4387 15268 4396 15308
rect 4436 15268 7372 15308
rect 7412 15268 7421 15308
rect 8899 15268 8908 15308
rect 8948 15268 15764 15308
rect 15724 15224 15764 15268
rect 16483 15268 16492 15308
rect 16532 15268 17452 15308
rect 17492 15268 17501 15308
rect 17635 15268 17644 15308
rect 17684 15268 19564 15308
rect 19604 15268 19613 15308
rect 20035 15268 20044 15308
rect 20084 15268 20180 15308
rect 16483 15267 16541 15268
rect 18499 15224 18557 15225
rect 3244 15184 3476 15224
rect 6979 15184 6988 15224
rect 7028 15184 12748 15224
rect 12788 15184 12797 15224
rect 15724 15184 17740 15224
rect 17780 15184 17789 15224
rect 18211 15184 18220 15224
rect 18260 15184 18508 15224
rect 18548 15184 18557 15224
rect 2467 15100 2476 15140
rect 2516 15100 2860 15140
rect 2900 15100 2909 15140
rect 3244 15056 3284 15184
rect 3331 15100 3340 15140
rect 3380 15100 3389 15140
rect 835 15016 844 15056
rect 884 15016 3284 15056
rect 3340 14972 3380 15100
rect 3436 15056 3476 15184
rect 18499 15183 18557 15184
rect 20803 15224 20861 15225
rect 21424 15224 21504 15244
rect 20803 15184 20812 15224
rect 20852 15184 21504 15224
rect 20803 15183 20861 15184
rect 21424 15164 21504 15184
rect 3679 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 4065 15140
rect 8035 15100 8044 15140
rect 8084 15100 8716 15140
rect 8756 15100 8765 15140
rect 8812 15100 12844 15140
rect 12884 15100 12893 15140
rect 17251 15100 17260 15140
rect 17300 15100 17932 15140
rect 17972 15100 17981 15140
rect 18799 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 19185 15140
rect 8812 15056 8852 15100
rect 3436 15016 5932 15056
rect 5972 15016 7564 15056
rect 7604 15016 7613 15056
rect 7939 15016 7948 15056
rect 7988 15016 8852 15056
rect 12163 15016 12172 15056
rect 12212 15016 12364 15056
rect 12404 15016 12413 15056
rect 13411 15016 13420 15056
rect 13460 15016 17836 15056
rect 17876 15016 17885 15056
rect 13420 14972 13460 15016
rect 3340 14932 6604 14972
rect 6644 14932 6653 14972
rect 8131 14932 8140 14972
rect 8180 14932 8428 14972
rect 8468 14932 8477 14972
rect 11587 14932 11596 14972
rect 11636 14932 13460 14972
rect 13507 14932 13516 14972
rect 13556 14932 14092 14972
rect 14132 14932 20180 14972
rect 3235 14888 3293 14889
rect 7939 14888 7997 14889
rect 8803 14888 8861 14889
rect 3235 14848 3244 14888
rect 3284 14848 4012 14888
rect 4052 14848 4300 14888
rect 4340 14848 4349 14888
rect 7939 14848 7948 14888
rect 7988 14848 8812 14888
rect 8852 14848 8947 14888
rect 9571 14848 9580 14888
rect 9620 14848 9964 14888
rect 10004 14848 10013 14888
rect 13987 14848 13996 14888
rect 14036 14848 14284 14888
rect 14324 14848 14333 14888
rect 16771 14848 16780 14888
rect 16820 14848 17356 14888
rect 17396 14848 17405 14888
rect 3235 14847 3293 14848
rect 7939 14847 7997 14848
rect 8803 14847 8861 14848
rect 5731 14804 5789 14805
rect 1228 14764 5740 14804
rect 5780 14764 5789 14804
rect 0 14720 80 14740
rect 1228 14720 1268 14764
rect 5731 14763 5789 14764
rect 6988 14764 10868 14804
rect 11299 14764 11308 14804
rect 11348 14764 13556 14804
rect 13603 14764 13612 14804
rect 13652 14764 19852 14804
rect 19892 14764 19901 14804
rect 3235 14720 3293 14721
rect 4195 14720 4253 14721
rect 0 14680 1268 14720
rect 1315 14680 1324 14720
rect 1364 14680 3244 14720
rect 3284 14680 3293 14720
rect 3523 14680 3532 14720
rect 3572 14680 3581 14720
rect 3715 14680 3724 14720
rect 3764 14680 4204 14720
rect 4244 14680 4253 14720
rect 5251 14680 5260 14720
rect 5300 14680 6028 14720
rect 6068 14680 6077 14720
rect 0 14660 80 14680
rect 3235 14679 3293 14680
rect 3532 14636 3572 14680
rect 4195 14679 4253 14680
rect 6988 14636 7028 14764
rect 7267 14680 7276 14720
rect 7316 14680 7948 14720
rect 7988 14680 7997 14720
rect 9187 14680 9196 14720
rect 9236 14680 9580 14720
rect 9620 14680 9629 14720
rect 10828 14636 10868 14764
rect 13516 14720 13556 14764
rect 18499 14720 18557 14721
rect 10915 14680 10924 14720
rect 10964 14680 11444 14720
rect 11491 14680 11500 14720
rect 11540 14680 12212 14720
rect 13516 14680 16780 14720
rect 16820 14680 17660 14720
rect 11404 14636 11444 14680
rect 11491 14636 11549 14637
rect 12067 14636 12125 14637
rect 3235 14596 3244 14636
rect 3284 14596 3436 14636
rect 3476 14596 3485 14636
rect 3532 14596 7028 14636
rect 10819 14596 10828 14636
rect 10868 14596 11116 14636
rect 11156 14596 11165 14636
rect 11404 14596 11500 14636
rect 11540 14596 11549 14636
rect 11982 14596 12076 14636
rect 12116 14596 12125 14636
rect 12172 14636 12212 14680
rect 17620 14636 17660 14680
rect 18499 14680 18508 14720
rect 18548 14680 19372 14720
rect 19412 14680 19421 14720
rect 19651 14680 19660 14720
rect 19700 14680 19948 14720
rect 19988 14680 19997 14720
rect 18499 14679 18557 14680
rect 12172 14596 15916 14636
rect 15956 14596 15965 14636
rect 17620 14596 18700 14636
rect 18740 14596 18749 14636
rect 3532 14552 3572 14596
rect 11491 14595 11549 14596
rect 12067 14595 12125 14596
rect 15139 14552 15197 14553
rect 20140 14552 20180 14932
rect 21424 14888 21504 14908
rect 20803 14848 20812 14888
rect 20852 14848 21504 14888
rect 21424 14828 21504 14848
rect 21424 14552 21504 14572
rect 1219 14512 1228 14552
rect 1268 14512 3572 14552
rect 4003 14512 4012 14552
rect 4052 14512 4396 14552
rect 4436 14512 4445 14552
rect 4492 14512 5260 14552
rect 5300 14512 5309 14552
rect 9955 14512 9964 14552
rect 10004 14512 14476 14552
rect 14516 14512 14525 14552
rect 15054 14512 15148 14552
rect 15188 14512 15197 14552
rect 17059 14512 17068 14552
rect 17108 14512 17548 14552
rect 17588 14512 17597 14552
rect 20140 14512 21504 14552
rect 4492 14384 4532 14512
rect 15139 14511 15197 14512
rect 21424 14492 21504 14512
rect 6115 14468 6173 14469
rect 19555 14468 19613 14469
rect 4579 14428 4588 14468
rect 4628 14428 6124 14468
rect 6164 14428 6173 14468
rect 8035 14428 8044 14468
rect 8084 14428 8524 14468
rect 8564 14428 8573 14468
rect 8707 14428 8716 14468
rect 8756 14428 18164 14468
rect 18595 14428 18604 14468
rect 18644 14428 19564 14468
rect 19604 14428 19660 14468
rect 19700 14428 19709 14468
rect 6115 14427 6173 14428
rect 15715 14384 15773 14385
rect 17059 14384 17117 14385
rect 18124 14384 18164 14428
rect 19555 14427 19613 14428
rect 19843 14384 19901 14385
rect 2947 14344 2956 14384
rect 2996 14344 4532 14384
rect 4919 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 5305 14384
rect 5827 14344 5836 14384
rect 5876 14344 6028 14384
rect 6068 14344 6077 14384
rect 6787 14344 6796 14384
rect 6836 14344 12172 14384
rect 12212 14344 12221 14384
rect 15715 14344 15724 14384
rect 15764 14344 16012 14384
rect 16052 14344 16061 14384
rect 17059 14344 17068 14384
rect 17108 14344 17164 14384
rect 17204 14344 17213 14384
rect 17539 14344 17548 14384
rect 17588 14344 18028 14384
rect 18068 14344 18077 14384
rect 18124 14344 19852 14384
rect 19892 14344 19901 14384
rect 20039 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20425 14384
rect 5836 14300 5876 14344
rect 15715 14343 15773 14344
rect 17059 14343 17117 14344
rect 19843 14343 19901 14344
rect 3811 14260 3820 14300
rect 3860 14260 5876 14300
rect 6115 14260 6124 14300
rect 6164 14260 6412 14300
rect 6452 14260 6461 14300
rect 7747 14260 7756 14300
rect 7796 14260 9524 14300
rect 11395 14260 11404 14300
rect 11444 14260 11884 14300
rect 11924 14260 11933 14300
rect 15907 14260 15916 14300
rect 15956 14260 16588 14300
rect 16628 14260 16637 14300
rect 17443 14260 17452 14300
rect 17492 14260 17836 14300
rect 17876 14260 17885 14300
rect 9484 14216 9524 14260
rect 21424 14216 21504 14236
rect 1795 14176 1804 14216
rect 1844 14176 2188 14216
rect 2228 14176 2237 14216
rect 3139 14176 3148 14216
rect 3188 14176 4108 14216
rect 4148 14176 4157 14216
rect 4579 14176 4588 14216
rect 4628 14176 4637 14216
rect 5155 14176 5164 14216
rect 5204 14176 7180 14216
rect 7220 14176 7229 14216
rect 8227 14176 8236 14216
rect 8276 14176 9388 14216
rect 9428 14176 9437 14216
rect 9484 14176 21504 14216
rect 4588 14132 4628 14176
rect 21424 14156 21504 14176
rect 2500 14092 4628 14132
rect 5243 14092 5252 14132
rect 5292 14092 6796 14132
rect 6836 14092 6845 14132
rect 7939 14092 7948 14132
rect 7988 14092 9580 14132
rect 9620 14092 9629 14132
rect 15523 14092 15532 14132
rect 15572 14092 16300 14132
rect 16340 14092 16349 14132
rect 0 14048 80 14068
rect 0 13988 116 14048
rect 76 13964 116 13988
rect 2500 13964 2540 14092
rect 3523 14048 3581 14049
rect 6115 14048 6173 14049
rect 3438 14008 3532 14048
rect 3572 14008 3581 14048
rect 3811 14008 3820 14048
rect 3860 14008 5740 14048
rect 5780 14008 5789 14048
rect 6030 14008 6124 14048
rect 6164 14008 6173 14048
rect 6691 14008 6700 14048
rect 6740 14008 9964 14048
rect 10004 14008 10156 14048
rect 10196 14008 10205 14048
rect 11203 14008 11212 14048
rect 11252 14008 12844 14048
rect 12884 14008 15436 14048
rect 15476 14008 15485 14048
rect 17347 14008 17356 14048
rect 17396 14008 17740 14048
rect 17780 14008 17789 14048
rect 3523 14007 3581 14008
rect 6115 14007 6173 14008
rect 4099 13964 4157 13965
rect 76 13924 2540 13964
rect 4003 13924 4012 13964
rect 4052 13924 4108 13964
rect 4148 13924 4157 13964
rect 4291 13924 4300 13964
rect 4340 13924 5644 13964
rect 5684 13924 6316 13964
rect 6356 13924 6365 13964
rect 7843 13924 7852 13964
rect 7892 13924 8428 13964
rect 8468 13924 8477 13964
rect 11320 13924 11596 13964
rect 11636 13924 11645 13964
rect 12355 13924 12364 13964
rect 12404 13924 20044 13964
rect 20084 13924 20093 13964
rect 4099 13923 4157 13924
rect 11320 13880 11360 13924
rect 4099 13840 4108 13880
rect 4148 13840 5836 13880
rect 5876 13840 5885 13880
rect 6595 13840 6604 13880
rect 6644 13840 6988 13880
rect 7028 13840 11360 13880
rect 11491 13880 11549 13881
rect 15715 13880 15773 13881
rect 18019 13880 18077 13881
rect 21424 13880 21504 13900
rect 11491 13840 11500 13880
rect 11540 13840 15724 13880
rect 15764 13840 15773 13880
rect 15907 13840 15916 13880
rect 15956 13840 17836 13880
rect 17876 13840 17885 13880
rect 18019 13840 18028 13880
rect 18068 13840 21504 13880
rect 11491 13839 11549 13840
rect 15715 13839 15773 13840
rect 18019 13839 18077 13840
rect 21424 13820 21504 13840
rect 4195 13796 4253 13797
rect 19267 13796 19325 13797
rect 4195 13756 4204 13796
rect 4244 13756 4972 13796
rect 5012 13756 6412 13796
rect 6452 13756 6461 13796
rect 13123 13756 13132 13796
rect 13172 13756 16012 13796
rect 16052 13756 16300 13796
rect 16340 13756 16349 13796
rect 18979 13756 18988 13796
rect 19028 13756 19276 13796
rect 19316 13756 19325 13796
rect 4195 13755 4253 13756
rect 19267 13755 19325 13756
rect 13987 13712 14045 13713
rect 1027 13672 1036 13712
rect 1076 13672 4684 13712
rect 4724 13672 4733 13712
rect 13891 13672 13900 13712
rect 13940 13672 13996 13712
rect 14036 13672 14045 13712
rect 14659 13672 14668 13712
rect 14708 13672 20716 13712
rect 20756 13672 20765 13712
rect 13987 13671 14045 13672
rect 5443 13628 5501 13629
rect 3679 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 4065 13628
rect 5155 13588 5164 13628
rect 5204 13588 5452 13628
rect 5492 13588 6028 13628
rect 6068 13588 6077 13628
rect 18799 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 19185 13628
rect 5443 13587 5501 13588
rect 8803 13544 8861 13545
rect 17251 13544 17309 13545
rect 21424 13544 21504 13564
rect 6115 13504 6124 13544
rect 6164 13504 6700 13544
rect 6740 13504 6749 13544
rect 7651 13504 7660 13544
rect 7700 13504 8044 13544
rect 8084 13504 8093 13544
rect 8803 13504 8812 13544
rect 8852 13504 8908 13544
rect 8948 13504 8957 13544
rect 9955 13504 9964 13544
rect 10004 13504 17260 13544
rect 17300 13504 17309 13544
rect 19267 13504 19276 13544
rect 19316 13504 21504 13544
rect 8803 13503 8861 13504
rect 17251 13503 17309 13504
rect 21424 13484 21504 13504
rect 163 13460 221 13461
rect 14851 13460 14909 13461
rect 163 13420 172 13460
rect 212 13420 11360 13460
rect 163 13419 221 13420
rect 0 13376 80 13396
rect 7747 13376 7805 13377
rect 0 13336 7756 13376
rect 7796 13336 7805 13376
rect 11320 13376 11360 13420
rect 14851 13420 14860 13460
rect 14900 13420 21196 13460
rect 21236 13420 21245 13460
rect 14851 13419 14909 13420
rect 11320 13336 19084 13376
rect 19124 13336 19133 13376
rect 0 13316 80 13336
rect 7747 13335 7805 13336
rect 4291 13292 4349 13293
rect 19939 13292 19997 13293
rect 1507 13252 1516 13292
rect 1556 13252 2956 13292
rect 2996 13252 3005 13292
rect 4003 13252 4012 13292
rect 4052 13252 4300 13292
rect 4340 13252 8716 13292
rect 8756 13252 8765 13292
rect 13516 13252 16396 13292
rect 16436 13252 19276 13292
rect 19316 13252 19325 13292
rect 19939 13252 19948 13292
rect 19988 13252 20044 13292
rect 20084 13252 20093 13292
rect 4291 13251 4349 13252
rect 4387 13208 4445 13209
rect 5635 13208 5693 13209
rect 6595 13208 6653 13209
rect 13516 13208 13556 13252
rect 19939 13251 19997 13252
rect 21424 13208 21504 13228
rect 1699 13168 1708 13208
rect 1748 13168 1996 13208
rect 2036 13168 2045 13208
rect 3907 13168 3916 13208
rect 3956 13168 4396 13208
rect 4436 13168 4588 13208
rect 4628 13168 4637 13208
rect 5550 13168 5644 13208
rect 5684 13168 5693 13208
rect 6499 13168 6508 13208
rect 6548 13168 6604 13208
rect 6644 13168 6653 13208
rect 7843 13168 7852 13208
rect 7892 13168 10636 13208
rect 10676 13168 10685 13208
rect 12067 13168 12076 13208
rect 12116 13168 13516 13208
rect 13556 13168 13565 13208
rect 13987 13168 13996 13208
rect 14036 13168 14380 13208
rect 14420 13168 14429 13208
rect 15235 13168 15244 13208
rect 15284 13168 15820 13208
rect 15860 13168 16204 13208
rect 16244 13168 16253 13208
rect 16483 13168 16492 13208
rect 16532 13168 17260 13208
rect 17300 13168 17309 13208
rect 20140 13168 21504 13208
rect 4387 13167 4445 13168
rect 5635 13167 5693 13168
rect 6595 13167 6653 13168
rect 14563 13124 14621 13125
rect 6883 13084 6892 13124
rect 6932 13084 7084 13124
rect 7124 13084 7133 13124
rect 11395 13084 11404 13124
rect 11444 13084 12940 13124
rect 12980 13084 12989 13124
rect 14563 13084 14572 13124
rect 14612 13084 14668 13124
rect 14708 13084 14717 13124
rect 15523 13084 15532 13124
rect 15572 13084 16108 13124
rect 16148 13084 16157 13124
rect 14563 13083 14621 13084
rect 20140 13040 20180 13168
rect 21424 13148 21504 13168
rect 3139 13000 3148 13040
rect 3188 13000 4108 13040
rect 4148 13000 4157 13040
rect 7363 13000 7372 13040
rect 7412 13000 7948 13040
rect 7988 13000 7997 13040
rect 9763 13000 9772 13040
rect 9812 13000 10828 13040
rect 10868 13000 10877 13040
rect 15715 13000 15724 13040
rect 15764 13000 20180 13040
rect 1699 12916 1708 12956
rect 1748 12916 7180 12956
rect 7220 12916 7229 12956
rect 8131 12916 8140 12956
rect 8180 12916 9868 12956
rect 9908 12916 10348 12956
rect 10388 12916 10397 12956
rect 11320 12916 20852 12956
rect 11320 12872 11360 12916
rect 20812 12872 20852 12916
rect 21424 12872 21504 12892
rect 4919 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 5305 12872
rect 5635 12832 5644 12872
rect 5684 12832 6124 12872
rect 6164 12832 6173 12872
rect 6403 12832 6412 12872
rect 6452 12832 7084 12872
rect 7124 12832 7133 12872
rect 7459 12832 7468 12872
rect 7508 12832 7852 12872
rect 7892 12832 11360 12872
rect 20039 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20425 12872
rect 20812 12832 21504 12872
rect 21424 12812 21504 12832
rect 1795 12748 1804 12788
rect 1844 12748 9964 12788
rect 10004 12748 10013 12788
rect 11395 12748 11404 12788
rect 11444 12748 11788 12788
rect 11828 12748 11837 12788
rect 12643 12748 12652 12788
rect 12692 12748 13708 12788
rect 13748 12748 13757 12788
rect 19459 12748 19468 12788
rect 19508 12748 19517 12788
rect 0 12704 80 12724
rect 3043 12704 3101 12705
rect 7363 12704 7421 12705
rect 0 12664 3052 12704
rect 3092 12664 3101 12704
rect 3331 12664 3340 12704
rect 3380 12664 3389 12704
rect 4291 12664 4300 12704
rect 4340 12664 5644 12704
rect 5684 12664 5693 12704
rect 5923 12664 5932 12704
rect 5972 12664 5981 12704
rect 7278 12664 7372 12704
rect 7412 12664 7421 12704
rect 0 12644 80 12664
rect 3043 12663 3101 12664
rect 3340 12620 3380 12664
rect 2851 12580 2860 12620
rect 2900 12580 3380 12620
rect 3523 12620 3581 12621
rect 5443 12620 5501 12621
rect 3523 12580 3532 12620
rect 3572 12580 3916 12620
rect 3956 12580 3965 12620
rect 4675 12580 4684 12620
rect 4724 12580 4876 12620
rect 4916 12580 4925 12620
rect 5251 12580 5260 12620
rect 5300 12580 5452 12620
rect 5492 12580 5501 12620
rect 5932 12620 5972 12664
rect 7363 12663 7421 12664
rect 8800 12664 9100 12704
rect 9140 12664 9149 12704
rect 13987 12664 13996 12704
rect 14036 12664 14284 12704
rect 14324 12664 14333 12704
rect 15139 12664 15148 12704
rect 15188 12664 15820 12704
rect 15860 12664 15869 12704
rect 16291 12664 16300 12704
rect 16340 12664 16972 12704
rect 17012 12664 17548 12704
rect 17588 12664 17597 12704
rect 8800 12620 8840 12664
rect 10147 12620 10205 12621
rect 19468 12620 19508 12748
rect 19555 12664 19564 12704
rect 19604 12664 19852 12704
rect 19892 12664 19901 12704
rect 5932 12580 6356 12620
rect 8323 12580 8332 12620
rect 8372 12580 8840 12620
rect 8995 12580 9004 12620
rect 9044 12580 10156 12620
rect 10196 12580 10205 12620
rect 10627 12580 10636 12620
rect 10676 12580 12940 12620
rect 12980 12580 12989 12620
rect 16579 12580 16588 12620
rect 16628 12580 18604 12620
rect 18644 12580 18653 12620
rect 19468 12580 20236 12620
rect 20276 12580 20285 12620
rect 3523 12579 3581 12580
rect 5443 12579 5501 12580
rect 3235 12536 3293 12537
rect 3811 12536 3869 12537
rect 6211 12536 6269 12537
rect 1411 12496 1420 12536
rect 1460 12496 1996 12536
rect 2036 12496 2045 12536
rect 3235 12496 3244 12536
rect 3284 12496 3340 12536
rect 3380 12496 3389 12536
rect 3523 12496 3532 12536
rect 3572 12496 3581 12536
rect 3726 12496 3820 12536
rect 3860 12496 3869 12536
rect 4003 12496 4012 12536
rect 4052 12496 5548 12536
rect 5588 12496 5597 12536
rect 5731 12496 5740 12536
rect 5780 12496 6220 12536
rect 6260 12496 6269 12536
rect 6316 12536 6356 12580
rect 10147 12579 10205 12580
rect 8419 12536 8477 12537
rect 21424 12536 21504 12556
rect 6316 12496 8140 12536
rect 8180 12496 8189 12536
rect 8419 12496 8428 12536
rect 8468 12496 13036 12536
rect 13076 12496 13085 12536
rect 14947 12496 14956 12536
rect 14996 12496 17932 12536
rect 17972 12496 17981 12536
rect 18499 12496 18508 12536
rect 18548 12496 18796 12536
rect 18836 12496 18845 12536
rect 19555 12496 19564 12536
rect 19604 12496 20812 12536
rect 20852 12496 20861 12536
rect 20908 12496 21504 12536
rect 3235 12495 3293 12496
rect 3532 12452 3572 12496
rect 3811 12495 3869 12496
rect 6211 12495 6269 12496
rect 8419 12495 8477 12496
rect 4771 12452 4829 12453
rect 20908 12452 20948 12496
rect 21424 12476 21504 12496
rect 2659 12412 2668 12452
rect 2708 12412 4396 12452
rect 4436 12412 4445 12452
rect 4771 12412 4780 12452
rect 4820 12412 4972 12452
rect 5012 12412 11308 12452
rect 11348 12412 11357 12452
rect 12259 12412 12268 12452
rect 12308 12412 12556 12452
rect 12596 12412 12605 12452
rect 12835 12412 12844 12452
rect 12884 12412 14284 12452
rect 14324 12412 14333 12452
rect 16003 12412 16012 12452
rect 16052 12412 16396 12452
rect 16436 12412 16780 12452
rect 16820 12412 16829 12452
rect 17059 12412 17068 12452
rect 17108 12412 17644 12452
rect 17684 12412 17693 12452
rect 20140 12412 20948 12452
rect 4771 12411 4829 12412
rect 16195 12368 16253 12369
rect 3427 12328 3436 12368
rect 3476 12328 4588 12368
rect 4628 12328 4637 12368
rect 5443 12328 5452 12368
rect 5492 12328 5932 12368
rect 5972 12328 5981 12368
rect 15139 12328 15148 12368
rect 15188 12328 16204 12368
rect 16244 12328 16253 12368
rect 16579 12328 16588 12368
rect 16628 12328 19564 12368
rect 19604 12328 19613 12368
rect 16195 12327 16253 12328
rect 3139 12244 3148 12284
rect 3188 12244 3340 12284
rect 3380 12244 5260 12284
rect 5300 12244 5309 12284
rect 9571 12244 9580 12284
rect 9620 12244 12076 12284
rect 12116 12244 12125 12284
rect 15619 12244 15628 12284
rect 15668 12244 16012 12284
rect 16052 12244 16061 12284
rect 16483 12244 16492 12284
rect 16532 12244 17164 12284
rect 17204 12244 17213 12284
rect 7267 12200 7325 12201
rect 20140 12200 20180 12412
rect 21424 12200 21504 12220
rect 2851 12160 2860 12200
rect 2900 12160 4340 12200
rect 4300 12116 4340 12160
rect 7267 12160 7276 12200
rect 7316 12160 7468 12200
rect 7508 12160 20180 12200
rect 20812 12160 21504 12200
rect 7267 12159 7325 12160
rect 16675 12116 16733 12117
rect 20812 12116 20852 12160
rect 21424 12140 21504 12160
rect 3679 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 4065 12116
rect 4291 12076 4300 12116
rect 4340 12076 4349 12116
rect 6220 12076 7220 12116
rect 7555 12076 7564 12116
rect 7604 12076 7948 12116
rect 7988 12076 7997 12116
rect 11299 12076 11308 12116
rect 11348 12076 11788 12116
rect 11828 12076 11837 12116
rect 13027 12076 13036 12116
rect 13076 12076 16684 12116
rect 16724 12076 16733 12116
rect 18799 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 19185 12116
rect 19363 12076 19372 12116
rect 19412 12076 20852 12116
rect 0 12032 80 12052
rect 1219 12032 1277 12033
rect 0 11992 1228 12032
rect 1268 11992 1277 12032
rect 0 11972 80 11992
rect 1219 11991 1277 11992
rect 3235 11948 3293 11949
rect 4195 11948 4253 11949
rect 6220 11948 6260 12076
rect 7180 12032 7220 12076
rect 16675 12075 16733 12076
rect 12163 12032 12221 12033
rect 7180 11992 8840 12032
rect 10051 11992 10060 12032
rect 10100 11992 11500 12032
rect 11540 11992 12172 12032
rect 12212 11992 12221 12032
rect 12931 11992 12940 12032
rect 12980 11992 16780 12032
rect 16820 11992 16829 12032
rect 3139 11908 3148 11948
rect 3188 11908 3244 11948
rect 3284 11908 3916 11948
rect 3956 11908 4204 11948
rect 4244 11908 4253 11948
rect 6211 11908 6220 11948
rect 6260 11908 6269 11948
rect 6403 11908 6412 11948
rect 6452 11908 7276 11948
rect 7316 11908 7325 11948
rect 3235 11907 3293 11908
rect 4195 11907 4253 11908
rect 8800 11864 8840 11992
rect 12163 11991 12221 11992
rect 10627 11908 10636 11948
rect 10676 11908 11884 11948
rect 11924 11908 11933 11948
rect 14851 11908 14860 11948
rect 14900 11908 17932 11948
rect 17972 11908 17981 11948
rect 1507 11824 1516 11864
rect 1556 11824 3052 11864
rect 3092 11824 3101 11864
rect 3427 11824 3436 11864
rect 3476 11824 3485 11864
rect 3715 11824 3724 11864
rect 3764 11824 4780 11864
rect 4820 11824 4829 11864
rect 4963 11824 4972 11864
rect 5012 11824 8236 11864
rect 8276 11824 8285 11864
rect 8800 11824 8812 11864
rect 8852 11824 11212 11864
rect 11252 11824 11261 11864
rect 3436 11780 3476 11824
rect 11884 11780 11924 11908
rect 21187 11864 21245 11865
rect 21424 11864 21504 11884
rect 12163 11824 12172 11864
rect 12212 11824 13268 11864
rect 15139 11824 15148 11864
rect 15188 11824 19372 11864
rect 19412 11824 19421 11864
rect 21187 11824 21196 11864
rect 21236 11824 21504 11864
rect 13228 11781 13268 11824
rect 21187 11823 21245 11824
rect 21424 11804 21504 11824
rect 13219 11780 13277 11781
rect 3436 11740 4492 11780
rect 4532 11740 6932 11780
rect 8323 11740 8332 11780
rect 8372 11740 8908 11780
rect 8948 11740 8957 11780
rect 11884 11740 12364 11780
rect 12404 11740 12413 11780
rect 13219 11740 13228 11780
rect 13268 11740 17012 11780
rect 6892 11696 6932 11740
rect 13219 11739 13277 11740
rect 16195 11696 16253 11697
rect 16972 11696 17012 11740
rect 17251 11696 17309 11697
rect 3235 11656 3244 11696
rect 3284 11656 4108 11696
rect 4148 11656 4157 11696
rect 4675 11656 4684 11696
rect 4724 11656 6604 11696
rect 6644 11656 6653 11696
rect 6883 11656 6892 11696
rect 6932 11656 6941 11696
rect 7555 11656 7564 11696
rect 7604 11656 10828 11696
rect 10868 11656 11020 11696
rect 11060 11656 11069 11696
rect 11587 11656 11596 11696
rect 11636 11656 12172 11696
rect 12212 11656 12221 11696
rect 14275 11656 14284 11696
rect 14324 11656 15148 11696
rect 15188 11656 15724 11696
rect 15764 11656 16204 11696
rect 16244 11656 16253 11696
rect 16963 11656 16972 11696
rect 17012 11656 17021 11696
rect 17166 11656 17260 11696
rect 17300 11656 17309 11696
rect 6604 11612 6644 11656
rect 16195 11655 16253 11656
rect 17251 11655 17309 11656
rect 6604 11572 9004 11612
rect 9044 11572 9196 11612
rect 9236 11572 9245 11612
rect 12067 11572 12076 11612
rect 12116 11572 14572 11612
rect 14612 11572 14621 11612
rect 15331 11572 15340 11612
rect 15380 11572 17068 11612
rect 17108 11572 17356 11612
rect 17396 11572 17405 11612
rect 18316 11572 20180 11612
rect 1315 11488 1324 11528
rect 1364 11488 3340 11528
rect 3380 11488 3389 11528
rect 4483 11488 4492 11528
rect 4532 11488 6124 11528
rect 6164 11488 7756 11528
rect 7796 11488 7805 11528
rect 9571 11488 9580 11528
rect 9620 11488 10060 11528
rect 10100 11488 10109 11528
rect 15523 11488 15532 11528
rect 15572 11488 18220 11528
rect 18260 11488 18269 11528
rect 6307 11444 6365 11445
rect 7939 11444 7997 11445
rect 1507 11404 1516 11444
rect 1556 11404 3476 11444
rect 6211 11404 6220 11444
rect 6260 11404 6316 11444
rect 6356 11404 6365 11444
rect 6595 11404 6604 11444
rect 6644 11404 7180 11444
rect 7220 11404 7229 11444
rect 7843 11404 7852 11444
rect 7892 11404 7948 11444
rect 7988 11404 7997 11444
rect 0 11360 80 11380
rect 3436 11360 3476 11404
rect 6307 11403 6365 11404
rect 7939 11403 7997 11404
rect 13795 11444 13853 11445
rect 16387 11444 16445 11445
rect 16867 11444 16925 11445
rect 18316 11444 18356 11572
rect 20140 11528 20180 11572
rect 21424 11528 21504 11548
rect 20140 11488 21504 11528
rect 21424 11468 21504 11488
rect 13795 11404 13804 11444
rect 13844 11404 13900 11444
rect 13940 11404 13949 11444
rect 16387 11404 16396 11444
rect 16436 11404 16588 11444
rect 16628 11404 16637 11444
rect 16867 11404 16876 11444
rect 16916 11404 18356 11444
rect 13795 11403 13853 11404
rect 16387 11403 16445 11404
rect 16867 11403 16925 11404
rect 13219 11360 13277 11361
rect 0 11320 460 11360
rect 500 11320 509 11360
rect 3396 11320 3436 11360
rect 3476 11320 3485 11360
rect 4919 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 5305 11360
rect 12931 11320 12940 11360
rect 12980 11320 13228 11360
rect 13268 11320 13277 11360
rect 13411 11320 13420 11360
rect 13460 11320 13469 11360
rect 17731 11320 17740 11360
rect 17780 11320 17789 11360
rect 20039 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20425 11360
rect 0 11300 80 11320
rect 13219 11319 13277 11320
rect 9379 11276 9437 11277
rect 12835 11276 12893 11277
rect 2083 11236 2092 11276
rect 2132 11236 2860 11276
rect 2900 11236 3724 11276
rect 3764 11236 3773 11276
rect 6595 11236 6604 11276
rect 6644 11236 7084 11276
rect 7124 11236 7133 11276
rect 9283 11236 9292 11276
rect 9332 11236 9388 11276
rect 9428 11236 9437 11276
rect 12739 11236 12748 11276
rect 12788 11236 12844 11276
rect 12884 11236 12893 11276
rect 9379 11235 9437 11236
rect 12835 11235 12893 11236
rect 13027 11276 13085 11277
rect 13027 11236 13036 11276
rect 13076 11236 13170 11276
rect 13027 11235 13085 11236
rect 1219 11152 1228 11192
rect 1268 11152 4204 11192
rect 4244 11152 5452 11192
rect 5492 11152 5932 11192
rect 5972 11152 5981 11192
rect 6499 11152 6508 11192
rect 6548 11152 10252 11192
rect 10292 11152 10301 11192
rect 10819 11152 10828 11192
rect 10868 11152 11212 11192
rect 11252 11152 12788 11192
rect 4099 11108 4157 11109
rect 8419 11108 8477 11109
rect 12067 11108 12125 11109
rect 12748 11108 12788 11152
rect 13420 11108 13460 11320
rect 16387 11276 16445 11277
rect 17740 11276 17780 11320
rect 13795 11236 13804 11276
rect 13844 11236 16396 11276
rect 16436 11236 16445 11276
rect 16579 11236 16588 11276
rect 16628 11236 17780 11276
rect 18019 11236 18028 11276
rect 18068 11236 18220 11276
rect 18260 11236 18269 11276
rect 18412 11236 18892 11276
rect 18932 11236 18941 11276
rect 16387 11235 16445 11236
rect 13795 11192 13853 11193
rect 13795 11152 13804 11192
rect 13844 11152 13996 11192
rect 14036 11152 14045 11192
rect 15907 11152 15916 11192
rect 15956 11152 15965 11192
rect 16963 11152 16972 11192
rect 17012 11152 17932 11192
rect 17972 11152 17981 11192
rect 13795 11151 13853 11152
rect 15916 11108 15956 11152
rect 18412 11108 18452 11236
rect 20131 11192 20189 11193
rect 21424 11192 21504 11212
rect 20131 11152 20140 11192
rect 20180 11152 21504 11192
rect 20131 11151 20189 11152
rect 21424 11132 21504 11152
rect 2467 11068 2476 11108
rect 2516 11068 2996 11108
rect 3523 11068 3532 11108
rect 3572 11068 4108 11108
rect 4148 11068 4157 11108
rect 2956 11024 2996 11068
rect 4099 11067 4157 11068
rect 5452 11068 8428 11108
rect 8468 11068 8477 11108
rect 8611 11068 8620 11108
rect 8660 11068 9388 11108
rect 9428 11068 10156 11108
rect 10196 11068 10205 11108
rect 11011 11068 11020 11108
rect 11060 11068 11308 11108
rect 11348 11068 11357 11108
rect 11683 11068 11692 11108
rect 11732 11068 12076 11108
rect 12116 11068 12125 11108
rect 12739 11068 12748 11108
rect 12788 11068 12797 11108
rect 13420 11068 13900 11108
rect 13940 11068 13949 11108
rect 14083 11068 14092 11108
rect 14132 11068 15052 11108
rect 15092 11068 15101 11108
rect 15916 11068 18452 11108
rect 4675 11024 4733 11025
rect 1315 10984 1324 11024
rect 1364 10984 2900 11024
rect 2947 10984 2956 11024
rect 2996 10984 4108 11024
rect 4148 10984 4157 11024
rect 4675 10984 4684 11024
rect 4724 10984 5164 11024
rect 5204 10984 5356 11024
rect 5396 10984 5405 11024
rect 2860 10940 2900 10984
rect 4675 10983 4733 10984
rect 5452 10940 5492 11068
rect 8419 11067 8477 11068
rect 12067 11067 12125 11068
rect 9571 11024 9629 11025
rect 5731 10984 5740 11024
rect 5780 10984 6316 11024
rect 6356 10984 6365 11024
rect 7171 10984 7180 11024
rect 7220 10984 9580 11024
rect 9620 10984 9629 11024
rect 10915 10984 10924 11024
rect 10964 10984 11404 11024
rect 11444 10984 11596 11024
rect 11636 10984 11645 11024
rect 15715 10984 15724 11024
rect 15764 10984 15916 11024
rect 15956 10984 16876 11024
rect 16916 10984 16925 11024
rect 17635 10984 17644 11024
rect 17684 10984 18508 11024
rect 18548 10984 18557 11024
rect 9571 10983 9629 10984
rect 1987 10900 1996 10940
rect 2036 10900 2540 10940
rect 2860 10900 5492 10940
rect 5827 10900 5836 10940
rect 5876 10900 6836 10940
rect 8419 10900 8428 10940
rect 8468 10900 8812 10940
rect 8852 10900 14668 10940
rect 14708 10900 14717 10940
rect 16003 10900 16012 10940
rect 16052 10900 16300 10940
rect 16340 10900 18260 10940
rect 259 10772 317 10773
rect 2500 10772 2540 10900
rect 6796 10856 6836 10900
rect 17251 10856 17309 10857
rect 18220 10856 18260 10900
rect 21424 10856 21504 10876
rect 3715 10816 3724 10856
rect 3764 10816 6740 10856
rect 6796 10816 13228 10856
rect 13268 10816 13277 10856
rect 13891 10816 13900 10856
rect 13940 10816 17068 10856
rect 17108 10816 17260 10856
rect 17300 10816 17309 10856
rect 17539 10816 17548 10856
rect 17588 10816 17740 10856
rect 17780 10816 17789 10856
rect 18211 10816 18220 10856
rect 18260 10816 18269 10856
rect 18883 10816 18892 10856
rect 18932 10816 21504 10856
rect 4099 10772 4157 10773
rect 6700 10772 6740 10816
rect 17251 10815 17309 10816
rect 21424 10796 21504 10816
rect 11779 10772 11837 10773
rect 259 10732 268 10772
rect 308 10732 1652 10772
rect 2500 10732 4108 10772
rect 4148 10732 4300 10772
rect 4340 10732 4349 10772
rect 4771 10732 4780 10772
rect 4820 10732 6604 10772
rect 6644 10732 6653 10772
rect 6700 10732 11788 10772
rect 11828 10732 13324 10772
rect 13364 10732 13373 10772
rect 259 10731 317 10732
rect 0 10688 80 10708
rect 1507 10688 1565 10689
rect 0 10648 1516 10688
rect 1556 10648 1565 10688
rect 1612 10688 1652 10732
rect 4099 10731 4157 10732
rect 11779 10731 11837 10732
rect 1612 10648 2540 10688
rect 6403 10648 6412 10688
rect 6452 10648 8140 10688
rect 8180 10648 8189 10688
rect 11587 10648 11596 10688
rect 11636 10648 11980 10688
rect 12020 10648 12029 10688
rect 17155 10648 17164 10688
rect 17204 10648 18028 10688
rect 18068 10648 18077 10688
rect 0 10628 80 10648
rect 1507 10647 1565 10648
rect 2500 10520 2540 10648
rect 3679 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 4065 10604
rect 5347 10564 5356 10604
rect 5396 10564 10540 10604
rect 10580 10564 10589 10604
rect 18799 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 19185 10604
rect 18019 10520 18077 10521
rect 18499 10520 18557 10521
rect 21424 10520 21504 10540
rect 2500 10480 17260 10520
rect 17300 10480 17309 10520
rect 17443 10480 17452 10520
rect 17492 10480 17740 10520
rect 17780 10480 17789 10520
rect 18019 10480 18028 10520
rect 18068 10480 18124 10520
rect 18164 10480 18173 10520
rect 18307 10480 18316 10520
rect 18356 10480 18508 10520
rect 18548 10480 18557 10520
rect 21187 10480 21196 10520
rect 21236 10480 21504 10520
rect 18019 10479 18077 10480
rect 18499 10479 18557 10480
rect 21424 10460 21504 10480
rect 6115 10436 6173 10437
rect 18211 10436 18269 10437
rect 4012 10396 6124 10436
rect 6164 10396 6173 10436
rect 10243 10396 10252 10436
rect 10292 10396 11596 10436
rect 11636 10396 11645 10436
rect 18211 10396 18220 10436
rect 18260 10396 18604 10436
rect 18644 10396 18653 10436
rect 67 10312 76 10352
rect 116 10312 3820 10352
rect 3860 10312 3869 10352
rect 4012 10184 4052 10396
rect 6115 10395 6173 10396
rect 18211 10395 18269 10396
rect 17923 10352 17981 10353
rect 5635 10312 5644 10352
rect 5684 10312 6988 10352
rect 7028 10312 7037 10352
rect 9772 10312 11212 10352
rect 11252 10312 11261 10352
rect 11875 10312 11884 10352
rect 11924 10312 12652 10352
rect 12692 10312 12701 10352
rect 17827 10312 17836 10352
rect 17876 10312 17932 10352
rect 17972 10312 17981 10352
rect 4099 10268 4157 10269
rect 9772 10268 9812 10312
rect 17923 10311 17981 10312
rect 9955 10268 10013 10269
rect 4099 10228 4108 10268
rect 4148 10228 7276 10268
rect 7316 10228 7325 10268
rect 8995 10228 9004 10268
rect 9044 10228 9772 10268
rect 9812 10228 9821 10268
rect 9955 10228 9964 10268
rect 10004 10228 10444 10268
rect 10484 10228 10493 10268
rect 16099 10228 16108 10268
rect 16148 10228 16972 10268
rect 17012 10228 18892 10268
rect 18932 10228 19948 10268
rect 19988 10228 19997 10268
rect 4099 10227 4157 10228
rect 9955 10227 10013 10228
rect 21424 10184 21504 10204
rect 2467 10144 2476 10184
rect 2516 10144 2525 10184
rect 3427 10144 3436 10184
rect 3476 10144 4052 10184
rect 4867 10144 4876 10184
rect 4916 10144 5260 10184
rect 5300 10144 5452 10184
rect 5492 10144 5501 10184
rect 7555 10144 7564 10184
rect 7604 10144 11404 10184
rect 11444 10144 11453 10184
rect 12547 10144 12556 10184
rect 12596 10144 15724 10184
rect 15764 10144 15773 10184
rect 16195 10144 16204 10184
rect 16244 10144 17932 10184
rect 17972 10144 17981 10184
rect 18028 10144 20140 10184
rect 20180 10144 20189 10184
rect 20707 10144 20716 10184
rect 20756 10144 21504 10184
rect 2476 10100 2516 10144
rect 3427 10100 3485 10101
rect 76 10060 212 10100
rect 2476 10060 2764 10100
rect 2804 10060 2813 10100
rect 2947 10060 2956 10100
rect 2996 10060 3436 10100
rect 3476 10060 3628 10100
rect 3668 10060 3677 10100
rect 6019 10060 6028 10100
rect 6068 10060 6356 10100
rect 76 10036 116 10060
rect 0 9976 116 10036
rect 0 9956 80 9976
rect 172 9848 212 10060
rect 3427 10059 3485 10060
rect 4195 10016 4253 10017
rect 6316 10016 6356 10060
rect 9772 10060 10348 10100
rect 10388 10060 10868 10100
rect 9772 10016 9812 10060
rect 10828 10016 10868 10060
rect 18028 10016 18068 10144
rect 21424 10124 21504 10144
rect 18691 10016 18749 10017
rect 3907 9976 3916 10016
rect 3956 9976 4204 10016
rect 4244 9976 4253 10016
rect 5150 9976 5159 10016
rect 5199 9976 5932 10016
rect 5972 9976 5981 10016
rect 6307 9976 6316 10016
rect 6356 9976 6365 10016
rect 9763 9976 9772 10016
rect 9812 9976 9821 10016
rect 10819 9976 10828 10016
rect 10868 9976 10877 10016
rect 13027 9976 13036 10016
rect 13076 9976 13516 10016
rect 13556 9976 13565 10016
rect 14371 9976 14380 10016
rect 14420 9976 15244 10016
rect 15284 9976 15293 10016
rect 16963 9976 16972 10016
rect 17012 9976 18028 10016
rect 18068 9976 18077 10016
rect 18595 9976 18604 10016
rect 18644 9976 18700 10016
rect 18740 9976 18749 10016
rect 4195 9975 4253 9976
rect 18691 9975 18749 9976
rect 20515 9932 20573 9933
rect 2500 9892 20524 9932
rect 20564 9892 20573 9932
rect 2500 9848 2540 9892
rect 20515 9891 20573 9892
rect 8803 9848 8861 9849
rect 13987 9848 14045 9849
rect 17923 9848 17981 9849
rect 19459 9848 19517 9849
rect 20803 9848 20861 9849
rect 21424 9848 21504 9868
rect 172 9808 2540 9848
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 5827 9808 5836 9848
rect 5876 9808 7084 9848
rect 7124 9808 7133 9848
rect 8803 9808 8812 9848
rect 8852 9808 9004 9848
rect 9044 9808 9053 9848
rect 13603 9808 13612 9848
rect 13652 9808 13661 9848
rect 13987 9808 13996 9848
rect 14036 9808 14956 9848
rect 14996 9808 15005 9848
rect 16675 9808 16684 9848
rect 16724 9808 17356 9848
rect 17396 9808 17405 9848
rect 17838 9808 17932 9848
rect 17972 9808 17981 9848
rect 19374 9808 19468 9848
rect 19508 9808 19517 9848
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 20803 9808 20812 9848
rect 20852 9808 21504 9848
rect 8803 9807 8861 9808
rect 8515 9764 8573 9765
rect 1795 9724 1804 9764
rect 1844 9724 2540 9764
rect 4675 9724 4684 9764
rect 4724 9724 6988 9764
rect 7028 9724 7037 9764
rect 8515 9724 8524 9764
rect 8564 9724 8716 9764
rect 8756 9724 8765 9764
rect 2500 9680 2540 9724
rect 8515 9723 8573 9724
rect 13612 9680 13652 9808
rect 13987 9807 14045 9808
rect 17923 9807 17981 9808
rect 19459 9807 19517 9808
rect 20803 9807 20861 9808
rect 21424 9788 21504 9808
rect 18019 9764 18077 9765
rect 13795 9724 13804 9764
rect 13844 9724 14860 9764
rect 14900 9724 14909 9764
rect 17934 9724 18028 9764
rect 18068 9724 18077 9764
rect 19267 9724 19276 9764
rect 19316 9724 21100 9764
rect 21140 9724 21149 9764
rect 18019 9723 18077 9724
rect 2500 9640 13652 9680
rect 14659 9640 14668 9680
rect 14708 9640 14900 9680
rect 18115 9640 18124 9680
rect 18164 9640 19084 9680
rect 19124 9640 19133 9680
rect 19363 9640 19372 9680
rect 19412 9640 21332 9680
rect 3907 9556 3916 9596
rect 3956 9556 5204 9596
rect 10915 9556 10924 9596
rect 10964 9556 12940 9596
rect 12980 9556 12989 9596
rect 1603 9512 1661 9513
rect 4387 9512 4445 9513
rect 5164 9512 5204 9556
rect 1518 9472 1612 9512
rect 1652 9472 1661 9512
rect 2851 9472 2860 9512
rect 2900 9472 3244 9512
rect 3284 9472 3293 9512
rect 3427 9472 3436 9512
rect 3476 9472 3628 9512
rect 3668 9472 3677 9512
rect 4302 9472 4396 9512
rect 4436 9472 4445 9512
rect 5155 9472 5164 9512
rect 5204 9472 5213 9512
rect 6403 9472 6412 9512
rect 6452 9472 6988 9512
rect 7028 9472 7037 9512
rect 8035 9472 8044 9512
rect 8084 9472 9964 9512
rect 10004 9472 10013 9512
rect 11320 9472 11692 9512
rect 11732 9472 12460 9512
rect 12500 9472 12509 9512
rect 1603 9471 1661 9472
rect 4387 9471 4445 9472
rect 11320 9428 11360 9472
rect 13612 9428 13652 9640
rect 13699 9472 13708 9512
rect 13748 9472 14284 9512
rect 14324 9472 14333 9512
rect 1891 9388 1900 9428
rect 1940 9388 11360 9428
rect 13603 9388 13612 9428
rect 13652 9388 13661 9428
rect 0 9344 80 9364
rect 2563 9344 2621 9345
rect 4291 9344 4349 9345
rect 6211 9344 6269 9345
rect 14860 9344 14900 9640
rect 16387 9556 16396 9596
rect 16436 9556 20084 9596
rect 16195 9512 16253 9513
rect 17443 9512 17501 9513
rect 19363 9512 19421 9513
rect 19555 9512 19613 9513
rect 20044 9512 20084 9556
rect 16195 9472 16204 9512
rect 16244 9472 16588 9512
rect 16628 9472 16637 9512
rect 17443 9472 17452 9512
rect 17492 9472 17644 9512
rect 17684 9472 17693 9512
rect 19277 9472 19367 9512
rect 19412 9472 19421 9512
rect 19470 9472 19564 9512
rect 19604 9472 19613 9512
rect 20035 9472 20044 9512
rect 20084 9472 20093 9512
rect 16195 9471 16253 9472
rect 17443 9471 17501 9472
rect 19363 9471 19421 9472
rect 19555 9471 19613 9472
rect 21292 9428 21332 9640
rect 21424 9512 21504 9532
rect 21388 9452 21504 9512
rect 21388 9428 21428 9452
rect 19651 9388 19660 9428
rect 19700 9388 20140 9428
rect 20180 9388 20189 9428
rect 21292 9388 21428 9428
rect 0 9304 2572 9344
rect 2612 9304 2621 9344
rect 2851 9304 2860 9344
rect 2900 9304 4300 9344
rect 4340 9304 4349 9344
rect 6126 9304 6220 9344
rect 6260 9304 6269 9344
rect 6883 9304 6892 9344
rect 6932 9304 9676 9344
rect 9716 9304 9725 9344
rect 14563 9304 14572 9344
rect 14612 9304 14900 9344
rect 18499 9304 18508 9344
rect 18548 9304 20236 9344
rect 20276 9304 20285 9344
rect 0 9284 80 9304
rect 2563 9303 2621 9304
rect 4291 9303 4349 9304
rect 6211 9303 6269 9304
rect 2572 9260 2612 9303
rect 2851 9260 2909 9261
rect 3619 9260 3677 9261
rect 4483 9260 4541 9261
rect 2572 9220 2860 9260
rect 2900 9220 2909 9260
rect 3427 9220 3436 9260
rect 3476 9220 3485 9260
rect 3619 9220 3628 9260
rect 3675 9220 3763 9260
rect 4398 9220 4492 9260
rect 4532 9220 4541 9260
rect 2851 9219 2909 9220
rect 3436 9176 3476 9220
rect 3619 9219 3677 9220
rect 4483 9219 4541 9220
rect 7363 9260 7421 9261
rect 7363 9220 7372 9260
rect 7412 9220 7468 9260
rect 7508 9220 7517 9260
rect 7363 9219 7421 9220
rect 9676 9176 9716 9304
rect 19075 9220 19084 9260
rect 19124 9220 19468 9260
rect 19508 9220 19517 9260
rect 20515 9176 20573 9177
rect 3436 9136 6988 9176
rect 7028 9136 7037 9176
rect 9676 9136 12556 9176
rect 12596 9136 12605 9176
rect 20430 9136 20524 9176
rect 20564 9136 20573 9176
rect 20515 9135 20573 9136
rect 20899 9176 20957 9177
rect 21424 9176 21504 9196
rect 20899 9136 20908 9176
rect 20948 9136 21504 9176
rect 20899 9135 20957 9136
rect 21424 9116 21504 9136
rect 6595 9092 6653 9093
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 6595 9052 6604 9092
rect 6644 9052 7372 9092
rect 7412 9052 7421 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 6595 9051 6653 9052
rect 3427 9008 3485 9009
rect 3427 8968 3436 9008
rect 3476 8968 3860 9008
rect 4483 8968 4492 9008
rect 4532 8968 4876 9008
rect 4916 8968 4925 9008
rect 11011 8968 11020 9008
rect 11060 8968 19372 9008
rect 19412 8968 19852 9008
rect 19892 8968 19901 9008
rect 3427 8967 3485 8968
rect 3523 8924 3581 8925
rect 3523 8884 3532 8924
rect 3572 8884 3628 8924
rect 3668 8884 3677 8924
rect 3523 8883 3581 8884
rect 3715 8840 3773 8841
rect 3820 8840 3860 8968
rect 3907 8884 3916 8924
rect 3956 8884 4972 8924
rect 5012 8884 5021 8924
rect 19075 8884 19084 8924
rect 19124 8884 19756 8924
rect 19796 8884 19805 8924
rect 20227 8884 20236 8924
rect 20276 8884 21196 8924
rect 21236 8884 21245 8924
rect 6307 8840 6365 8841
rect 9379 8840 9437 8841
rect 20131 8840 20189 8841
rect 21424 8840 21504 8860
rect 3630 8800 3724 8840
rect 3764 8800 3773 8840
rect 3818 8800 3827 8840
rect 3867 8800 3876 8840
rect 4771 8800 4780 8840
rect 4820 8800 5548 8840
rect 5588 8800 5597 8840
rect 6115 8800 6124 8840
rect 6164 8800 6316 8840
rect 6356 8800 8140 8840
rect 8180 8800 8189 8840
rect 9294 8800 9388 8840
rect 9428 8800 9437 8840
rect 11299 8800 11308 8840
rect 11348 8800 11788 8840
rect 11828 8800 11837 8840
rect 14659 8800 14668 8840
rect 14708 8800 15340 8840
rect 15380 8800 15389 8840
rect 17155 8800 17164 8840
rect 17204 8800 17836 8840
rect 17876 8800 17885 8840
rect 20131 8800 20140 8840
rect 20180 8800 21504 8840
rect 3715 8799 3773 8800
rect 6307 8799 6365 8800
rect 9379 8799 9437 8800
rect 20131 8799 20189 8800
rect 21424 8780 21504 8800
rect 5635 8756 5693 8757
rect 4675 8716 4684 8756
rect 4724 8716 5644 8756
rect 5684 8716 6316 8756
rect 6356 8716 6365 8756
rect 7075 8716 7084 8756
rect 7124 8716 9292 8756
rect 9332 8716 9580 8756
rect 9620 8716 9629 8756
rect 5635 8715 5693 8716
rect 0 8672 80 8692
rect 19459 8672 19517 8673
rect 0 8632 364 8672
rect 404 8632 413 8672
rect 3331 8632 3340 8672
rect 3380 8632 4012 8672
rect 4052 8632 4396 8672
rect 4436 8632 4445 8672
rect 4867 8632 4876 8672
rect 4916 8632 11212 8672
rect 11252 8632 11692 8672
rect 11732 8632 11741 8672
rect 12451 8632 12460 8672
rect 12500 8632 12940 8672
rect 12980 8632 12989 8672
rect 15427 8632 15436 8672
rect 15476 8632 16012 8672
rect 16052 8632 16061 8672
rect 17635 8632 17644 8672
rect 17684 8632 17693 8672
rect 19459 8632 19468 8672
rect 19508 8632 19564 8672
rect 19604 8632 19613 8672
rect 0 8612 80 8632
rect 4099 8588 4157 8589
rect 9187 8588 9245 8589
rect 17644 8588 17684 8632
rect 19459 8631 19517 8632
rect 3043 8548 3052 8588
rect 3092 8548 3916 8588
rect 3956 8548 4108 8588
rect 4148 8548 4780 8588
rect 4820 8548 4829 8588
rect 9187 8548 9196 8588
rect 9236 8548 11360 8588
rect 13603 8548 13612 8588
rect 13652 8548 13996 8588
rect 14036 8548 17684 8588
rect 4099 8547 4157 8548
rect 9187 8547 9245 8548
rect 4483 8504 4541 8505
rect 11320 8504 11360 8548
rect 21424 8504 21504 8524
rect 4195 8464 4204 8504
rect 4244 8464 4492 8504
rect 4532 8464 4541 8504
rect 8899 8464 8908 8504
rect 8948 8464 9292 8504
rect 9332 8464 9341 8504
rect 11320 8464 13324 8504
rect 13364 8464 15532 8504
rect 15572 8464 17644 8504
rect 17684 8464 17693 8504
rect 20140 8464 21504 8504
rect 4483 8463 4541 8464
rect 12835 8420 12893 8421
rect 20140 8420 20180 8464
rect 21424 8444 21504 8464
rect 2947 8380 2956 8420
rect 2996 8380 3148 8420
rect 3188 8380 4492 8420
rect 4532 8380 4684 8420
rect 4724 8380 5836 8420
rect 5876 8380 5885 8420
rect 6307 8380 6316 8420
rect 6356 8380 7276 8420
rect 7316 8380 9196 8420
rect 9236 8380 9245 8420
rect 12067 8380 12076 8420
rect 12116 8380 12460 8420
rect 12500 8380 12509 8420
rect 12835 8380 12844 8420
rect 12884 8380 12940 8420
rect 12980 8380 12989 8420
rect 15724 8380 20180 8420
rect 4108 8336 4148 8380
rect 12835 8379 12893 8380
rect 3235 8296 3244 8336
rect 3284 8296 3628 8336
rect 3668 8296 3677 8336
rect 4099 8296 4108 8336
rect 4148 8296 4157 8336
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 7171 8296 7180 8336
rect 7220 8296 8812 8336
rect 8852 8296 9484 8336
rect 9524 8296 9533 8336
rect 2371 8212 2380 8252
rect 2420 8212 5836 8252
rect 5876 8212 5885 8252
rect 3523 8128 3532 8168
rect 3572 8128 3916 8168
rect 3956 8128 3965 8168
rect 4099 8128 4108 8168
rect 4148 8128 6028 8168
rect 6068 8128 6077 8168
rect 7171 8128 7180 8168
rect 7220 8128 10196 8168
rect 11107 8128 11116 8168
rect 11156 8128 13420 8168
rect 13460 8128 13469 8168
rect 13891 8128 13900 8168
rect 13940 8128 14476 8168
rect 14516 8128 14860 8168
rect 14900 8128 14909 8168
rect 0 8000 80 8020
rect 4771 8000 4829 8001
rect 7555 8000 7613 8001
rect 8227 8000 8285 8001
rect 9187 8000 9245 8001
rect 0 7960 2516 8000
rect 2947 7960 2956 8000
rect 2996 7960 3532 8000
rect 3572 7960 3581 8000
rect 4771 7960 4780 8000
rect 4820 7960 4972 8000
rect 5012 7960 5021 8000
rect 7555 7960 7564 8000
rect 7604 7960 8236 8000
rect 8276 7960 8285 8000
rect 8899 7960 8908 8000
rect 8948 7960 9196 8000
rect 9236 7960 9245 8000
rect 0 7940 80 7960
rect 2476 7664 2516 7960
rect 4771 7959 4829 7960
rect 7555 7959 7613 7960
rect 8227 7959 8285 7960
rect 9187 7959 9245 7960
rect 8035 7876 8044 7916
rect 8084 7876 9964 7916
rect 10004 7876 10013 7916
rect 10156 7832 10196 8128
rect 11683 8044 11692 8084
rect 11732 8044 12748 8084
rect 12788 8044 12797 8084
rect 13411 7960 13420 8000
rect 13460 7960 13612 8000
rect 13652 7960 13661 8000
rect 11491 7876 11500 7916
rect 11540 7876 11788 7916
rect 11828 7876 11837 7916
rect 13420 7832 13460 7960
rect 2563 7792 2572 7832
rect 2612 7792 8852 7832
rect 10156 7792 13460 7832
rect 7555 7748 7613 7749
rect 8812 7748 8852 7792
rect 15724 7748 15764 8380
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 21424 8168 21504 8188
rect 17251 8128 17260 8168
rect 17300 8128 19756 8168
rect 19796 8128 19805 8168
rect 19939 8128 19948 8168
rect 19988 8128 20140 8168
rect 20180 8128 20189 8168
rect 20707 8128 20716 8168
rect 20756 8128 20765 8168
rect 21091 8128 21100 8168
rect 21140 8128 21504 8168
rect 20716 8084 20756 8128
rect 21424 8108 21504 8128
rect 19564 8044 20756 8084
rect 19267 8000 19325 8001
rect 19564 8000 19604 8044
rect 18883 7960 18892 8000
rect 18932 7960 19276 8000
rect 19316 7960 19325 8000
rect 19555 7960 19564 8000
rect 19604 7960 19613 8000
rect 19939 7960 19948 8000
rect 19988 7960 19997 8000
rect 19267 7959 19325 7960
rect 19948 7916 19988 7960
rect 19171 7876 19180 7916
rect 19220 7876 19988 7916
rect 20035 7876 20044 7916
rect 20084 7876 20093 7916
rect 20044 7832 20084 7876
rect 21424 7832 21504 7852
rect 19372 7792 19756 7832
rect 19796 7792 20084 7832
rect 21292 7792 21504 7832
rect 19372 7749 19412 7792
rect 19363 7748 19421 7749
rect 5452 7708 7564 7748
rect 7604 7708 7613 7748
rect 7747 7708 7756 7748
rect 7796 7708 8716 7748
rect 8756 7708 8765 7748
rect 8812 7708 15764 7748
rect 19075 7708 19084 7748
rect 19124 7708 19372 7748
rect 19412 7708 19421 7748
rect 5452 7664 5492 7708
rect 7555 7707 7613 7708
rect 19363 7707 19421 7708
rect 13411 7664 13469 7665
rect 21292 7664 21332 7792
rect 21424 7772 21504 7792
rect 2476 7624 5492 7664
rect 6307 7624 6316 7664
rect 6356 7624 6604 7664
rect 6644 7624 11360 7664
rect 11320 7580 11360 7624
rect 13411 7624 13420 7664
rect 13460 7624 21332 7664
rect 13411 7623 13469 7624
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 4195 7540 4204 7580
rect 4244 7540 4780 7580
rect 4820 7540 4829 7580
rect 7459 7540 7468 7580
rect 7508 7540 8812 7580
rect 8852 7540 8861 7580
rect 11320 7540 15052 7580
rect 15092 7540 15101 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 4675 7496 4733 7497
rect 4590 7456 4684 7496
rect 4724 7456 4733 7496
rect 4675 7455 4733 7456
rect 5347 7496 5405 7497
rect 21424 7496 21504 7516
rect 5347 7456 5356 7496
rect 5396 7456 5876 7496
rect 7747 7456 7756 7496
rect 7796 7456 8428 7496
rect 8468 7456 9676 7496
rect 9716 7456 10156 7496
rect 10196 7456 10924 7496
rect 10964 7456 10973 7496
rect 11020 7456 21504 7496
rect 5347 7455 5405 7456
rect 5836 7412 5876 7456
rect 11020 7412 11060 7456
rect 21424 7436 21504 7456
rect 4483 7372 4492 7412
rect 4532 7372 5740 7412
rect 5780 7372 5789 7412
rect 5836 7372 11060 7412
rect 11320 7372 18988 7412
rect 19028 7372 19037 7412
rect 0 7329 80 7348
rect 0 7328 125 7329
rect 0 7288 76 7328
rect 116 7288 125 7328
rect 0 7287 125 7288
rect 2563 7328 2621 7329
rect 11320 7328 11360 7372
rect 2563 7288 2572 7328
rect 2612 7288 11360 7328
rect 12355 7288 12364 7328
rect 12404 7288 12652 7328
rect 12692 7288 12701 7328
rect 13699 7288 13708 7328
rect 13748 7288 16492 7328
rect 16532 7288 16541 7328
rect 18787 7288 18796 7328
rect 18836 7288 19372 7328
rect 19412 7288 19421 7328
rect 2563 7287 2621 7288
rect 0 7268 80 7287
rect 13123 7204 13132 7244
rect 13172 7204 15916 7244
rect 15956 7204 15965 7244
rect 7459 7160 7517 7161
rect 20131 7160 20189 7161
rect 21424 7160 21504 7180
rect 7459 7120 7468 7160
rect 7508 7120 10924 7160
rect 10964 7120 10973 7160
rect 12739 7120 12748 7160
rect 12788 7120 13516 7160
rect 13556 7120 13565 7160
rect 14851 7120 14860 7160
rect 14900 7120 15436 7160
rect 15476 7120 15485 7160
rect 18691 7120 18700 7160
rect 18740 7120 19412 7160
rect 7459 7119 7517 7120
rect 17155 7076 17213 7077
rect 13219 7036 13228 7076
rect 13268 7036 15532 7076
rect 15572 7036 15581 7076
rect 17070 7036 17164 7076
rect 17204 7036 17213 7076
rect 19372 7076 19412 7120
rect 20131 7120 20140 7160
rect 20180 7120 21504 7160
rect 20131 7119 20189 7120
rect 21424 7100 21504 7120
rect 19372 7036 20180 7076
rect 17155 7035 17213 7036
rect 19267 6992 19325 6993
rect 19555 6992 19613 6993
rect 9955 6952 9964 6992
rect 10004 6952 10156 6992
rect 10196 6952 10205 6992
rect 13315 6952 13324 6992
rect 13364 6952 14380 6992
rect 14420 6952 14429 6992
rect 18595 6952 18604 6992
rect 18644 6952 19276 6992
rect 19316 6952 19325 6992
rect 19470 6952 19564 6992
rect 19604 6952 19613 6992
rect 19267 6951 19325 6952
rect 19555 6951 19613 6952
rect 20140 6908 20180 7036
rect 11320 6868 14092 6908
rect 14132 6868 14141 6908
rect 20140 6868 21332 6908
rect 11320 6824 11360 6868
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 9955 6784 9964 6824
rect 10004 6784 11360 6824
rect 12067 6784 12076 6824
rect 12116 6784 19756 6824
rect 19796 6784 19805 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 16387 6740 16445 6741
rect 17443 6740 17501 6741
rect 19564 6740 19604 6784
rect 21292 6740 21332 6868
rect 21424 6824 21504 6844
rect 21388 6764 21504 6824
rect 21388 6740 21428 6764
rect 15523 6700 15532 6740
rect 15572 6700 15820 6740
rect 15860 6700 15869 6740
rect 16387 6700 16396 6740
rect 16436 6700 17452 6740
rect 17492 6700 18700 6740
rect 18740 6700 18749 6740
rect 19555 6700 19564 6740
rect 19604 6700 19644 6740
rect 21292 6700 21428 6740
rect 16387 6699 16445 6700
rect 17443 6699 17501 6700
rect 14947 6616 14956 6656
rect 14996 6616 21332 6656
rect 16387 6572 16445 6573
rect 11320 6532 13420 6572
rect 13460 6532 16396 6572
rect 16436 6532 16445 6572
rect 16675 6532 16684 6572
rect 16724 6532 18028 6572
rect 18068 6532 18077 6572
rect 11320 6488 11360 6532
rect 16387 6531 16445 6532
rect 21292 6488 21332 6616
rect 21424 6488 21504 6508
rect 8419 6448 8428 6488
rect 8468 6448 11360 6488
rect 11491 6448 11500 6488
rect 11540 6448 11636 6488
rect 12163 6448 12172 6488
rect 12212 6448 13996 6488
rect 14036 6448 14045 6488
rect 16483 6448 16492 6488
rect 16532 6448 17932 6488
rect 17972 6448 17981 6488
rect 21292 6448 21504 6488
rect 11596 6320 11636 6448
rect 21424 6428 21504 6448
rect 16867 6364 16876 6404
rect 16916 6364 18604 6404
rect 18644 6364 19948 6404
rect 19988 6364 19997 6404
rect 10243 6280 10252 6320
rect 10292 6280 11500 6320
rect 11540 6280 11549 6320
rect 11596 6280 12076 6320
rect 12116 6280 12125 6320
rect 13987 6280 13996 6320
rect 14036 6280 16972 6320
rect 17012 6280 17021 6320
rect 14659 6196 14668 6236
rect 14708 6196 16396 6236
rect 16436 6196 17164 6236
rect 17204 6196 17213 6236
rect 19843 6152 19901 6153
rect 21424 6152 21504 6172
rect 19843 6112 19852 6152
rect 19892 6112 21504 6152
rect 19843 6111 19901 6112
rect 21424 6092 21504 6112
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 11491 6028 11500 6068
rect 11540 6028 11884 6068
rect 11924 6028 11933 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 21424 5816 21504 5836
rect 6979 5776 6988 5816
rect 7028 5776 21504 5816
rect 21424 5756 21504 5776
rect 12451 5524 12460 5564
rect 12500 5524 20180 5564
rect 19459 5480 19517 5481
rect 19374 5440 19468 5480
rect 19508 5440 19517 5480
rect 20140 5480 20180 5524
rect 21424 5480 21504 5500
rect 20140 5440 21504 5480
rect 19459 5439 19517 5440
rect 21424 5420 21504 5440
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 21424 5144 21504 5164
rect 12067 5104 12076 5144
rect 12116 5104 21504 5144
rect 21424 5084 21504 5104
rect 12355 5060 12413 5061
rect 20707 5060 20765 5061
rect 12355 5020 12364 5060
rect 12404 5020 12748 5060
rect 12788 5020 12797 5060
rect 14755 5020 14764 5060
rect 14804 5020 15532 5060
rect 15572 5020 15581 5060
rect 19939 5020 19948 5060
rect 19988 5020 20716 5060
rect 20756 5020 20765 5060
rect 12355 5019 12413 5020
rect 20707 5019 20765 5020
rect 21424 4808 21504 4828
rect 8707 4768 8716 4808
rect 8756 4768 21504 4808
rect 21424 4748 21504 4768
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 21424 4472 21504 4492
rect 9283 4432 9292 4472
rect 9332 4432 21504 4472
rect 21424 4412 21504 4432
rect 21424 4136 21504 4156
rect 9763 4096 9772 4136
rect 9812 4096 10444 4136
rect 10484 4096 10493 4136
rect 15907 4096 15916 4136
rect 15956 4096 21504 4136
rect 21424 4076 21504 4096
rect 13027 3844 13036 3884
rect 13076 3844 20852 3884
rect 20812 3800 20852 3844
rect 21424 3800 21504 3820
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 6403 3760 6412 3800
rect 6452 3760 7852 3800
rect 7892 3760 7901 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 20812 3760 21504 3800
rect 21424 3740 21504 3760
rect 9955 3716 10013 3717
rect 3139 3676 3148 3716
rect 3188 3676 9964 3716
rect 10004 3676 10013 3716
rect 9955 3675 10013 3676
rect 15139 3592 15148 3632
rect 15188 3592 17356 3632
rect 17396 3592 17405 3632
rect 6211 3464 6269 3465
rect 21424 3464 21504 3484
rect 6211 3424 6220 3464
rect 6260 3424 21504 3464
rect 6211 3423 6269 3424
rect 21424 3404 21504 3424
rect 3331 3172 3340 3212
rect 3380 3172 15916 3212
rect 15956 3172 15965 3212
rect 21424 3128 21504 3148
rect 12931 3088 12940 3128
rect 12980 3088 21504 3128
rect 21424 3068 21504 3088
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 931 2876 989 2877
rect 931 2836 940 2876
rect 980 2836 6892 2876
rect 6932 2836 6941 2876
rect 931 2835 989 2836
rect 21424 2792 21504 2812
rect 11971 2752 11980 2792
rect 12020 2752 21504 2792
rect 21424 2732 21504 2752
rect 13795 2708 13853 2709
rect 14371 2708 14429 2709
rect 13710 2668 13804 2708
rect 13844 2668 13853 2708
rect 14286 2668 14380 2708
rect 14420 2668 14429 2708
rect 13795 2667 13853 2668
rect 14371 2667 14429 2668
rect 9580 2584 11360 2624
rect 9580 2540 9620 2584
rect 9571 2500 9580 2540
rect 9620 2500 9629 2540
rect 11320 2456 11360 2584
rect 21424 2456 21504 2476
rect 11320 2416 14284 2456
rect 14324 2416 14333 2456
rect 14563 2416 14572 2456
rect 14612 2416 15148 2456
rect 15188 2416 15197 2456
rect 20140 2416 21504 2456
rect 451 2372 509 2373
rect 20140 2372 20180 2416
rect 21424 2396 21504 2416
rect 451 2332 460 2372
rect 500 2332 7660 2372
rect 7700 2332 7709 2372
rect 11875 2332 11884 2372
rect 11924 2332 20180 2372
rect 451 2331 509 2332
rect 17731 2288 17789 2289
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 17731 2248 17740 2288
rect 17780 2248 18796 2288
rect 18836 2248 18845 2288
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 17731 2247 17789 2248
rect 1027 2204 1085 2205
rect 1027 2164 1036 2204
rect 1076 2164 6124 2204
rect 6164 2164 6173 2204
rect 8803 2164 8812 2204
rect 8852 2164 20180 2204
rect 1027 2163 1085 2164
rect 5731 2120 5789 2121
rect 6499 2120 6557 2121
rect 6883 2120 6941 2121
rect 7267 2120 7325 2121
rect 13891 2120 13949 2121
rect 15427 2120 15485 2121
rect 5646 2080 5740 2120
rect 5780 2080 5789 2120
rect 6414 2080 6508 2120
rect 6548 2080 6557 2120
rect 6798 2080 6892 2120
rect 6932 2080 6941 2120
rect 7182 2080 7276 2120
rect 7316 2080 7325 2120
rect 13806 2080 13900 2120
rect 13940 2080 14572 2120
rect 14612 2080 14621 2120
rect 15235 2080 15244 2120
rect 15284 2080 15436 2120
rect 15476 2080 15485 2120
rect 5731 2079 5789 2080
rect 6499 2079 6557 2080
rect 6883 2079 6941 2080
rect 7267 2079 7325 2080
rect 13891 2079 13949 2080
rect 15427 2079 15485 2080
rect 16291 2120 16349 2121
rect 17539 2120 17597 2121
rect 18115 2120 18173 2121
rect 16291 2080 16300 2120
rect 16340 2080 17260 2120
rect 17300 2080 17309 2120
rect 17539 2080 17548 2120
rect 17588 2080 17644 2120
rect 17684 2080 17693 2120
rect 18019 2080 18028 2120
rect 18068 2080 18124 2120
rect 18164 2080 18173 2120
rect 16291 2079 16349 2080
rect 17539 2079 17597 2080
rect 18115 2079 18173 2080
rect 18307 2120 18365 2121
rect 18595 2120 18653 2121
rect 19555 2120 19613 2121
rect 18307 2080 18316 2120
rect 18356 2080 18412 2120
rect 18452 2080 18461 2120
rect 18595 2080 18604 2120
rect 18644 2080 19180 2120
rect 19220 2080 19229 2120
rect 19470 2080 19564 2120
rect 19604 2080 19613 2120
rect 20140 2120 20180 2164
rect 21424 2120 21504 2140
rect 20140 2080 21504 2120
rect 18307 2079 18365 2080
rect 18595 2079 18653 2080
rect 19555 2079 19613 2080
rect 21424 2060 21504 2080
rect 7075 1996 7084 2036
rect 7124 1996 7756 2036
rect 7796 1996 7805 2036
rect 8995 1996 9004 2036
rect 9044 1996 9053 2036
rect 9379 1996 9388 2036
rect 9428 1996 9437 2036
rect 9004 1952 9044 1996
rect 4099 1912 4108 1952
rect 4148 1912 9044 1952
rect 8131 1868 8189 1869
rect 6691 1828 6700 1868
rect 6740 1828 7948 1868
rect 7988 1828 7997 1868
rect 8046 1828 8140 1868
rect 8180 1828 8189 1868
rect 8131 1827 8189 1828
rect 9388 1784 9428 1996
rect 9667 1912 9676 1952
rect 9716 1912 21428 1952
rect 10531 1868 10589 1869
rect 10915 1868 10973 1869
rect 11683 1868 11741 1869
rect 10446 1828 10540 1868
rect 10580 1828 10589 1868
rect 10830 1828 10924 1868
rect 10964 1828 10973 1868
rect 11598 1828 11692 1868
rect 11732 1828 11741 1868
rect 10531 1827 10589 1828
rect 10915 1827 10973 1828
rect 11683 1827 11741 1828
rect 11971 1868 12029 1869
rect 14275 1868 14333 1869
rect 14659 1868 14717 1869
rect 11971 1828 11980 1868
rect 12020 1828 12076 1868
rect 12116 1828 12125 1868
rect 14190 1828 14284 1868
rect 14324 1828 14333 1868
rect 14574 1828 14668 1868
rect 14708 1828 14717 1868
rect 11971 1827 12029 1828
rect 14275 1827 14333 1828
rect 14659 1827 14717 1828
rect 15523 1868 15581 1869
rect 16003 1868 16061 1869
rect 16387 1868 16445 1869
rect 15523 1828 15532 1868
rect 15572 1828 15628 1868
rect 15668 1828 15677 1868
rect 15811 1828 15820 1868
rect 15860 1828 15869 1868
rect 15918 1828 16012 1868
rect 16052 1828 16061 1868
rect 16302 1828 16396 1868
rect 16436 1828 16445 1868
rect 15523 1827 15581 1828
rect 15427 1784 15485 1785
rect 9388 1744 9812 1784
rect 15342 1744 15436 1784
rect 15476 1744 15485 1784
rect 15820 1784 15860 1828
rect 16003 1827 16061 1828
rect 16387 1827 16445 1828
rect 16579 1868 16637 1869
rect 16579 1828 16588 1868
rect 16628 1828 16780 1868
rect 16820 1828 16829 1868
rect 17539 1828 17548 1868
rect 17588 1828 17836 1868
rect 17876 1828 17885 1868
rect 16579 1827 16637 1828
rect 21388 1804 21428 1912
rect 15820 1744 21292 1784
rect 21332 1744 21341 1784
rect 21388 1744 21504 1804
rect 9772 1700 9812 1744
rect 15427 1743 15485 1744
rect 21424 1724 21504 1744
rect 8323 1660 8332 1700
rect 8372 1660 8908 1700
rect 8948 1660 8957 1700
rect 9763 1660 9772 1700
rect 9812 1660 9821 1700
rect 10051 1660 10060 1700
rect 10100 1660 11308 1700
rect 11348 1660 11357 1700
rect 12739 1660 12748 1700
rect 12788 1660 14476 1700
rect 14516 1660 14525 1700
rect 14851 1660 14860 1700
rect 14900 1660 16204 1700
rect 16244 1660 16253 1700
rect 18499 1660 18508 1700
rect 18548 1660 18988 1700
rect 19028 1660 19037 1700
rect 11320 1576 19508 1616
rect 11320 1532 11360 1576
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 5923 1492 5932 1532
rect 5972 1492 7276 1532
rect 7316 1492 7325 1532
rect 8419 1492 8428 1532
rect 8468 1492 11360 1532
rect 13891 1492 13900 1532
rect 13940 1492 15820 1532
rect 15860 1492 15869 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 19363 1492 19372 1532
rect 19412 1492 19421 1532
rect 6307 1408 6316 1448
rect 6356 1408 7564 1448
rect 7604 1408 7613 1448
rect 10819 1408 10828 1448
rect 10868 1408 13132 1448
rect 13172 1408 13181 1448
rect 15427 1408 15436 1448
rect 15476 1408 16588 1448
rect 16628 1408 16637 1448
rect 7075 1324 7084 1364
rect 7124 1324 8140 1364
rect 8180 1324 8189 1364
rect 10723 1324 10732 1364
rect 10772 1324 10781 1364
rect 11875 1324 11884 1364
rect 11924 1324 14476 1364
rect 14516 1324 14525 1364
rect 15523 1324 15532 1364
rect 15572 1324 15820 1364
rect 15860 1324 15869 1364
rect 18499 1324 18508 1364
rect 18548 1324 18557 1364
rect 2947 1280 3005 1281
rect 2862 1240 2956 1280
rect 2996 1240 3005 1280
rect 2947 1239 3005 1240
rect 3139 1280 3197 1281
rect 6787 1280 6845 1281
rect 9763 1280 9821 1281
rect 10732 1280 10772 1324
rect 15427 1280 15485 1281
rect 15619 1280 15677 1281
rect 3139 1240 3148 1280
rect 3188 1240 6028 1280
rect 6068 1240 6077 1280
rect 6280 1240 6508 1280
rect 6548 1240 6557 1280
rect 6702 1240 6796 1280
rect 6836 1240 6845 1280
rect 7459 1240 7468 1280
rect 7508 1240 8332 1280
rect 8372 1240 8381 1280
rect 9763 1240 9772 1280
rect 9812 1240 10388 1280
rect 10732 1240 12172 1280
rect 12212 1240 12221 1280
rect 13699 1240 13708 1280
rect 13748 1240 15436 1280
rect 15476 1240 15485 1280
rect 15534 1240 15628 1280
rect 15668 1240 15677 1280
rect 3139 1239 3197 1240
rect 1795 1196 1853 1197
rect 6280 1196 6320 1240
rect 6787 1239 6845 1240
rect 9763 1239 9821 1240
rect 10348 1196 10388 1240
rect 15427 1239 15485 1240
rect 15619 1239 15677 1240
rect 17827 1280 17885 1281
rect 18403 1280 18461 1281
rect 17827 1240 17836 1280
rect 17876 1240 18028 1280
rect 18068 1240 18077 1280
rect 18318 1240 18412 1280
rect 18452 1240 18461 1280
rect 17827 1239 17885 1240
rect 18403 1239 18461 1240
rect 11587 1196 11645 1197
rect 13027 1196 13085 1197
rect 13411 1196 13469 1197
rect 14947 1196 15005 1197
rect 16099 1196 16157 1197
rect 1795 1156 1804 1196
rect 1844 1156 6320 1196
rect 6691 1156 6700 1196
rect 6740 1156 7372 1196
rect 7412 1156 7421 1196
rect 9379 1156 9388 1196
rect 9428 1156 9868 1196
rect 9908 1156 9917 1196
rect 10339 1156 10348 1196
rect 10388 1156 10397 1196
rect 11502 1156 11596 1196
rect 11636 1156 11645 1196
rect 12942 1156 13036 1196
rect 13076 1156 13085 1196
rect 13326 1156 13420 1196
rect 13460 1156 13469 1196
rect 13795 1156 13804 1196
rect 13844 1156 14804 1196
rect 14862 1156 14956 1196
rect 14996 1156 15005 1196
rect 16014 1156 16108 1196
rect 16148 1156 16157 1196
rect 1795 1155 1853 1156
rect 11587 1155 11645 1156
rect 13027 1155 13085 1156
rect 13411 1155 13469 1156
rect 3331 1112 3389 1113
rect 12739 1112 12797 1113
rect 3331 1072 3340 1112
rect 3380 1072 6604 1112
rect 6644 1072 6653 1112
rect 8227 1072 8236 1112
rect 8276 1072 10772 1112
rect 11203 1072 11212 1112
rect 11252 1072 11980 1112
rect 12020 1072 12029 1112
rect 12076 1072 12748 1112
rect 12788 1072 12797 1112
rect 14764 1112 14804 1156
rect 14947 1155 15005 1156
rect 16099 1155 16157 1156
rect 15523 1112 15581 1113
rect 14764 1072 15532 1112
rect 15572 1072 15581 1112
rect 3331 1071 3389 1072
rect 8995 1028 9053 1029
rect 10627 1028 10685 1029
rect 5347 988 5356 1028
rect 5396 988 9004 1028
rect 9044 988 9053 1028
rect 8995 987 9053 988
rect 9292 988 10636 1028
rect 10676 988 10685 1028
rect 10732 1028 10772 1072
rect 12076 1028 12116 1072
rect 12739 1071 12797 1072
rect 15523 1071 15581 1072
rect 18508 1028 18548 1324
rect 19372 1280 19412 1492
rect 19468 1364 19508 1576
rect 21424 1448 21504 1468
rect 21379 1408 21388 1448
rect 21428 1408 21504 1448
rect 21424 1388 21504 1408
rect 19468 1324 20524 1364
rect 20564 1324 20573 1364
rect 18700 1240 19412 1280
rect 18700 1112 18740 1240
rect 21424 1112 21504 1132
rect 18691 1072 18700 1112
rect 18740 1072 18749 1112
rect 21292 1072 21504 1112
rect 10732 988 12116 1028
rect 12547 988 12556 1028
rect 12596 988 14092 1028
rect 14132 988 14141 1028
rect 18403 988 18412 1028
rect 18452 988 18548 1028
rect 2563 904 2572 944
rect 2612 904 6412 944
rect 6452 904 6461 944
rect 7843 904 7852 944
rect 7892 904 8524 944
rect 8564 904 8573 944
rect 8707 904 8716 944
rect 8756 904 9196 944
rect 9236 904 9245 944
rect 8323 860 8381 861
rect 9292 860 9332 988
rect 10627 987 10685 988
rect 19171 944 19229 945
rect 10531 904 10540 944
rect 10580 904 11212 944
rect 11252 904 11261 944
rect 13603 904 13612 944
rect 13652 904 14284 944
rect 14324 904 14333 944
rect 14659 904 14668 944
rect 14708 904 15916 944
rect 15956 904 15965 944
rect 19086 904 19180 944
rect 19220 904 19229 944
rect 19171 903 19229 904
rect 3523 820 3532 860
rect 3572 820 8332 860
rect 8372 820 8381 860
rect 8323 819 8381 820
rect 8428 820 9332 860
rect 9955 820 9964 860
rect 10004 820 10636 860
rect 10676 820 10685 860
rect 12931 820 12940 860
rect 12980 820 15052 860
rect 15092 820 15101 860
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 5635 736 5644 776
rect 5684 736 8236 776
rect 8276 736 8285 776
rect 8428 692 8468 820
rect 8803 736 8812 776
rect 8852 736 9868 776
rect 9908 736 9917 776
rect 10243 736 10252 776
rect 10292 736 11020 776
rect 11060 736 11069 776
rect 12643 736 12652 776
rect 12692 736 15668 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 15628 692 15668 736
rect 21292 692 21332 1072
rect 21424 1052 21504 1072
rect 21424 776 21504 796
rect 6280 652 8468 692
rect 9475 652 9484 692
rect 9524 652 15532 692
rect 15572 652 15581 692
rect 15628 652 21332 692
rect 21388 716 21504 776
rect 739 608 797 609
rect 6280 608 6320 652
rect 9475 608 9533 609
rect 21388 608 21428 716
rect 739 568 748 608
rect 788 568 2764 608
rect 2804 568 2813 608
rect 5443 568 5452 608
rect 5492 568 6320 608
rect 6988 568 9484 608
rect 9524 568 9533 608
rect 739 567 797 568
rect 6988 524 7028 568
rect 9475 567 9533 568
rect 20140 568 21428 608
rect 4291 484 4300 524
rect 4340 484 7028 524
rect 7075 484 7084 524
rect 7124 484 9100 524
rect 9140 484 9149 524
rect 12931 484 12940 524
rect 12980 484 14764 524
rect 14804 484 14813 524
rect 11875 440 11933 441
rect 6403 400 6412 440
rect 6452 400 11884 440
rect 11924 400 11933 440
rect 13315 400 13324 440
rect 13364 400 15148 440
rect 15188 400 15197 440
rect 11875 399 11933 400
rect 10051 356 10109 357
rect 3907 316 3916 356
rect 3956 316 10060 356
rect 10100 316 10109 356
rect 13123 316 13132 356
rect 13172 316 14380 356
rect 14420 316 14429 356
rect 17923 316 17932 356
rect 17972 316 18316 356
rect 18356 316 18365 356
rect 10051 315 10109 316
rect 5059 272 5117 273
rect 20140 272 20180 568
rect 21424 440 21504 460
rect 20515 400 20524 440
rect 20564 400 21504 440
rect 21424 380 21504 400
rect 4974 232 5068 272
rect 5108 232 5117 272
rect 9763 232 9772 272
rect 9812 232 20180 272
rect 5059 231 5117 232
rect 4867 188 4925 189
rect 12931 188 12989 189
rect 4782 148 4876 188
rect 4916 148 4925 188
rect 6211 148 6220 188
rect 6260 148 12940 188
rect 12980 148 12989 188
rect 17635 148 17644 188
rect 17684 148 17693 188
rect 4867 147 4925 148
rect 12931 147 12989 148
rect 3331 104 3389 105
rect 13507 104 13565 105
rect 3246 64 3340 104
rect 3380 64 3389 104
rect 6979 64 6988 104
rect 7028 64 13516 104
rect 13556 64 13565 104
rect 17644 104 17684 148
rect 21424 104 21504 124
rect 17644 64 21504 104
rect 3331 63 3389 64
rect 13507 63 13565 64
rect 21424 44 21504 64
<< via3 >>
rect 19084 85912 19124 85952
rect 19276 85912 19316 85952
rect 6508 85576 6548 85616
rect 16012 85576 16052 85616
rect 16876 85576 16916 85616
rect 2380 85156 2420 85196
rect 17932 85072 17972 85112
rect 19852 85072 19892 85112
rect 16396 84904 16436 84944
rect 20620 84904 20660 84944
rect 3688 84652 3728 84692
rect 3770 84652 3810 84692
rect 3852 84652 3892 84692
rect 3934 84652 3974 84692
rect 4016 84652 4056 84692
rect 18808 84652 18848 84692
rect 18890 84652 18930 84692
rect 18972 84652 19012 84692
rect 19054 84652 19094 84692
rect 19136 84652 19176 84692
rect 13900 84568 13940 84608
rect 20716 84568 20756 84608
rect 6892 84484 6932 84524
rect 14284 84484 14324 84524
rect 14956 84484 14996 84524
rect 16780 84484 16820 84524
rect 17740 84484 17780 84524
rect 18604 84484 18644 84524
rect 5836 84400 5876 84440
rect 6220 84400 6260 84440
rect 6796 84400 6836 84440
rect 10636 84400 10676 84440
rect 12172 84400 12212 84440
rect 13324 84400 13364 84440
rect 13708 84400 13748 84440
rect 13996 84400 14036 84440
rect 14668 84400 14708 84440
rect 15052 84400 15092 84440
rect 15532 84400 15572 84440
rect 17260 84400 17300 84440
rect 17548 84400 17588 84440
rect 17836 84400 17876 84440
rect 18412 84400 18452 84440
rect 19660 84400 19700 84440
rect 8908 84316 8948 84356
rect 4928 83896 4968 83936
rect 5010 83896 5050 83936
rect 5092 83896 5132 83936
rect 5174 83896 5214 83936
rect 5256 83896 5296 83936
rect 20048 83896 20088 83936
rect 20130 83896 20170 83936
rect 20212 83896 20252 83936
rect 20294 83896 20334 83936
rect 20376 83896 20416 83936
rect 10924 83560 10964 83600
rect 1516 83476 1556 83516
rect 2092 83476 2132 83516
rect 2284 83476 2324 83516
rect 7180 83476 7220 83516
rect 7372 83476 7412 83516
rect 8140 83476 8180 83516
rect 13612 83476 13652 83516
rect 15340 83476 15380 83516
rect 16204 83476 16244 83516
rect 2668 83308 2708 83348
rect 3688 83140 3728 83180
rect 3770 83140 3810 83180
rect 3852 83140 3892 83180
rect 3934 83140 3974 83180
rect 4016 83140 4056 83180
rect 6988 83140 7028 83180
rect 8236 83140 8276 83180
rect 18808 83140 18848 83180
rect 18890 83140 18930 83180
rect 18972 83140 19012 83180
rect 19054 83140 19094 83180
rect 19136 83140 19176 83180
rect 2860 82804 2900 82844
rect 3244 82804 3284 82844
rect 3532 82804 3572 82844
rect 19276 82720 19316 82760
rect 4928 82384 4968 82424
rect 5010 82384 5050 82424
rect 5092 82384 5132 82424
rect 5174 82384 5214 82424
rect 5256 82384 5296 82424
rect 20048 82384 20088 82424
rect 20130 82384 20170 82424
rect 20212 82384 20252 82424
rect 20294 82384 20334 82424
rect 20376 82384 20416 82424
rect 21388 82048 21428 82088
rect 3688 81628 3728 81668
rect 3770 81628 3810 81668
rect 3852 81628 3892 81668
rect 3934 81628 3974 81668
rect 4016 81628 4056 81668
rect 18808 81628 18848 81668
rect 18890 81628 18930 81668
rect 18972 81628 19012 81668
rect 19054 81628 19094 81668
rect 19136 81628 19176 81668
rect 4928 80872 4968 80912
rect 5010 80872 5050 80912
rect 5092 80872 5132 80912
rect 5174 80872 5214 80912
rect 5256 80872 5296 80912
rect 20048 80872 20088 80912
rect 20130 80872 20170 80912
rect 20212 80872 20252 80912
rect 20294 80872 20334 80912
rect 20376 80872 20416 80912
rect 3688 80116 3728 80156
rect 3770 80116 3810 80156
rect 3852 80116 3892 80156
rect 3934 80116 3974 80156
rect 4016 80116 4056 80156
rect 18808 80116 18848 80156
rect 18890 80116 18930 80156
rect 18972 80116 19012 80156
rect 19054 80116 19094 80156
rect 19136 80116 19176 80156
rect 4928 79360 4968 79400
rect 5010 79360 5050 79400
rect 5092 79360 5132 79400
rect 5174 79360 5214 79400
rect 5256 79360 5296 79400
rect 20048 79360 20088 79400
rect 20130 79360 20170 79400
rect 20212 79360 20252 79400
rect 20294 79360 20334 79400
rect 20376 79360 20416 79400
rect 11116 79276 11156 79316
rect 11980 79024 12020 79064
rect 11116 78940 11156 78980
rect 20524 78772 20564 78812
rect 3688 78604 3728 78644
rect 3770 78604 3810 78644
rect 3852 78604 3892 78644
rect 3934 78604 3974 78644
rect 4016 78604 4056 78644
rect 18808 78604 18848 78644
rect 18890 78604 18930 78644
rect 18972 78604 19012 78644
rect 19054 78604 19094 78644
rect 19136 78604 19176 78644
rect 20812 78520 20852 78560
rect 19564 78352 19604 78392
rect 10252 78100 10292 78140
rect 16972 78100 17012 78140
rect 20812 77932 20852 77972
rect 76 77848 116 77888
rect 4928 77848 4968 77888
rect 5010 77848 5050 77888
rect 5092 77848 5132 77888
rect 5174 77848 5214 77888
rect 5256 77848 5296 77888
rect 20048 77848 20088 77888
rect 20130 77848 20170 77888
rect 20212 77848 20252 77888
rect 20294 77848 20334 77888
rect 20376 77848 20416 77888
rect 20524 77680 20564 77720
rect 17068 77596 17108 77636
rect 10444 77428 10484 77468
rect 16588 77428 16628 77468
rect 19756 77428 19796 77468
rect 1516 77176 1556 77216
rect 17068 77176 17108 77216
rect 3688 77092 3728 77132
rect 3770 77092 3810 77132
rect 3852 77092 3892 77132
rect 3934 77092 3974 77132
rect 4016 77092 4056 77132
rect 18808 77092 18848 77132
rect 18890 77092 18930 77132
rect 18972 77092 19012 77132
rect 19054 77092 19094 77132
rect 19136 77092 19176 77132
rect 13420 76924 13460 76964
rect 19948 76756 19988 76796
rect 8524 76672 8564 76712
rect 9004 76672 9044 76712
rect 13516 76672 13556 76712
rect 12940 76588 12980 76628
rect 652 76504 692 76544
rect 11020 76504 11060 76544
rect 19468 76504 19508 76544
rect 19564 76420 19604 76460
rect 4928 76336 4968 76376
rect 5010 76336 5050 76376
rect 5092 76336 5132 76376
rect 5174 76336 5214 76376
rect 5256 76336 5296 76376
rect 20048 76336 20088 76376
rect 20130 76336 20170 76376
rect 20212 76336 20252 76376
rect 20294 76336 20334 76376
rect 20376 76336 20416 76376
rect 10444 76252 10484 76292
rect 12940 76252 12980 76292
rect 15148 76000 15188 76040
rect 18892 75916 18932 75956
rect 268 75832 308 75872
rect 10348 75832 10388 75872
rect 12076 75664 12116 75704
rect 19756 75664 19796 75704
rect 3688 75580 3728 75620
rect 3770 75580 3810 75620
rect 3852 75580 3892 75620
rect 3934 75580 3974 75620
rect 4016 75580 4056 75620
rect 18808 75580 18848 75620
rect 18890 75580 18930 75620
rect 18972 75580 19012 75620
rect 19054 75580 19094 75620
rect 19136 75580 19176 75620
rect 13420 75496 13460 75536
rect 19468 75496 19508 75536
rect 1804 75160 1844 75200
rect 17068 75160 17108 75200
rect 4928 74824 4968 74864
rect 5010 74824 5050 74864
rect 5092 74824 5132 74864
rect 5174 74824 5214 74864
rect 5256 74824 5296 74864
rect 20048 74824 20088 74864
rect 20130 74824 20170 74864
rect 20212 74824 20252 74864
rect 20294 74824 20334 74864
rect 20376 74824 20416 74864
rect 8620 74488 8660 74528
rect 9388 74488 9428 74528
rect 13516 74488 13556 74528
rect 8812 74404 8852 74444
rect 11884 74404 11924 74444
rect 3688 74068 3728 74108
rect 3770 74068 3810 74108
rect 3852 74068 3892 74108
rect 3934 74068 3974 74108
rect 4016 74068 4056 74108
rect 18808 74068 18848 74108
rect 18890 74068 18930 74108
rect 18972 74068 19012 74108
rect 19054 74068 19094 74108
rect 19136 74068 19176 74108
rect 15148 73984 15188 74024
rect 16300 73984 16340 74024
rect 19948 73984 19988 74024
rect 19852 73900 19892 73940
rect 5356 73816 5396 73856
rect 6412 73816 6452 73856
rect 6028 73648 6068 73688
rect 8716 73648 8756 73688
rect 9100 73648 9140 73688
rect 18700 73648 18740 73688
rect 11884 73564 11924 73604
rect 4928 73312 4968 73352
rect 5010 73312 5050 73352
rect 5092 73312 5132 73352
rect 5174 73312 5214 73352
rect 5256 73312 5296 73352
rect 20048 73312 20088 73352
rect 20130 73312 20170 73352
rect 20212 73312 20252 73352
rect 20294 73312 20334 73352
rect 20376 73312 20416 73352
rect 18124 73228 18164 73268
rect 12268 73144 12308 73184
rect 17932 73060 17972 73100
rect 20140 73060 20180 73100
rect 12268 72976 12308 73016
rect 11596 72892 11636 72932
rect 20140 72892 20180 72932
rect 17164 72808 17204 72848
rect 18124 72808 18164 72848
rect 21388 72808 21428 72848
rect 3688 72556 3728 72596
rect 3770 72556 3810 72596
rect 3852 72556 3892 72596
rect 3934 72556 3974 72596
rect 4016 72556 4056 72596
rect 172 72472 212 72512
rect 11596 72640 11636 72680
rect 18808 72556 18848 72596
rect 18890 72556 18930 72596
rect 18972 72556 19012 72596
rect 19054 72556 19094 72596
rect 19136 72556 19176 72596
rect 18700 72388 18740 72428
rect 4300 72220 4340 72260
rect 19756 72220 19796 72260
rect 19948 72220 19988 72260
rect 16492 72136 16532 72176
rect 17164 71968 17204 72008
rect 1900 71800 1940 71840
rect 4928 71800 4968 71840
rect 5010 71800 5050 71840
rect 5092 71800 5132 71840
rect 5174 71800 5214 71840
rect 5256 71800 5296 71840
rect 14860 71800 14900 71840
rect 15436 71800 15476 71840
rect 20048 71800 20088 71840
rect 20130 71800 20170 71840
rect 20212 71800 20252 71840
rect 20294 71800 20334 71840
rect 20376 71800 20416 71840
rect 5356 71548 5396 71588
rect 19948 71632 19988 71672
rect 9292 71464 9332 71504
rect 15436 71464 15476 71504
rect 16300 71464 16340 71504
rect 11884 71296 11924 71336
rect 16492 71212 16532 71252
rect 364 71128 404 71168
rect 17932 71128 17972 71168
rect 3688 71044 3728 71084
rect 3770 71044 3810 71084
rect 3852 71044 3892 71084
rect 3934 71044 3974 71084
rect 4016 71044 4056 71084
rect 14860 71044 14900 71084
rect 18808 71044 18848 71084
rect 18890 71044 18930 71084
rect 18972 71044 19012 71084
rect 19054 71044 19094 71084
rect 19136 71044 19176 71084
rect 17068 70960 17108 71000
rect 17644 70792 17684 70832
rect 9868 70708 9908 70748
rect 13420 70708 13460 70748
rect 5548 70624 5588 70664
rect 4492 70456 4532 70496
rect 14092 70540 14132 70580
rect 14860 70540 14900 70580
rect 16108 70540 16148 70580
rect 4928 70288 4968 70328
rect 5010 70288 5050 70328
rect 5092 70288 5132 70328
rect 5174 70288 5214 70328
rect 5256 70288 5296 70328
rect 20048 70288 20088 70328
rect 20130 70288 20170 70328
rect 20212 70288 20252 70328
rect 20294 70288 20334 70328
rect 20376 70288 20416 70328
rect 16972 70036 17012 70076
rect 6604 69952 6644 69992
rect 8332 69952 8372 69992
rect 14956 69868 14996 69908
rect 15148 69868 15188 69908
rect 2188 69784 2228 69824
rect 15820 69784 15860 69824
rect 16492 69784 16532 69824
rect 17932 69700 17972 69740
rect 3688 69532 3728 69572
rect 3770 69532 3810 69572
rect 3852 69532 3892 69572
rect 3934 69532 3974 69572
rect 4016 69532 4056 69572
rect 18808 69532 18848 69572
rect 18890 69532 18930 69572
rect 18972 69532 19012 69572
rect 19054 69532 19094 69572
rect 19136 69532 19176 69572
rect 4108 69280 4148 69320
rect 9004 69280 9044 69320
rect 17452 69280 17492 69320
rect 15628 69196 15668 69236
rect 18028 69196 18068 69236
rect 556 69112 596 69152
rect 4492 69112 4532 69152
rect 5644 69112 5684 69152
rect 17644 68944 17684 68984
rect 4928 68776 4968 68816
rect 5010 68776 5050 68816
rect 5092 68776 5132 68816
rect 5174 68776 5214 68816
rect 5256 68776 5296 68816
rect 20048 68776 20088 68816
rect 20130 68776 20170 68816
rect 20212 68776 20252 68816
rect 20294 68776 20334 68816
rect 20376 68776 20416 68816
rect 10924 68692 10964 68732
rect 20716 68692 20756 68732
rect 15052 68608 15092 68648
rect 15436 68608 15476 68648
rect 17644 68608 17684 68648
rect 748 68440 788 68480
rect 4108 68356 4148 68396
rect 6796 68356 6836 68396
rect 11404 68272 11444 68312
rect 14092 68272 14132 68312
rect 14572 68188 14612 68228
rect 17644 68104 17684 68144
rect 3688 68020 3728 68060
rect 3770 68020 3810 68060
rect 3852 68020 3892 68060
rect 3934 68020 3974 68060
rect 4016 68020 4056 68060
rect 18124 68020 18164 68060
rect 18808 68020 18848 68060
rect 18890 68020 18930 68060
rect 18972 68020 19012 68060
rect 19054 68020 19094 68060
rect 19136 68020 19176 68060
rect 16588 67852 16628 67892
rect 5548 67516 5588 67556
rect 18124 67516 18164 67556
rect 6604 67348 6644 67388
rect 14956 67348 14996 67388
rect 16972 67348 17012 67388
rect 4928 67264 4968 67304
rect 5010 67264 5050 67304
rect 5092 67264 5132 67304
rect 5174 67264 5214 67304
rect 5256 67264 5296 67304
rect 20048 67264 20088 67304
rect 20130 67264 20170 67304
rect 20212 67264 20252 67304
rect 20294 67264 20334 67304
rect 20376 67264 20416 67304
rect 1036 67096 1076 67136
rect 6316 67096 6356 67136
rect 4396 67012 4436 67052
rect 6124 66928 6164 66968
rect 8428 66844 8468 66884
rect 11788 66760 11828 66800
rect 3688 66508 3728 66548
rect 3770 66508 3810 66548
rect 3852 66508 3892 66548
rect 3934 66508 3974 66548
rect 4016 66508 4056 66548
rect 18808 66508 18848 66548
rect 18890 66508 18930 66548
rect 18972 66508 19012 66548
rect 19054 66508 19094 66548
rect 19136 66508 19176 66548
rect 17932 66088 17972 66128
rect 4108 66004 4148 66044
rect 16972 65920 17012 65960
rect 18028 65920 18068 65960
rect 1228 65752 1268 65792
rect 4928 65752 4968 65792
rect 5010 65752 5050 65792
rect 5092 65752 5132 65792
rect 5174 65752 5214 65792
rect 5256 65752 5296 65792
rect 20048 65752 20088 65792
rect 20130 65752 20170 65792
rect 20212 65752 20252 65792
rect 20294 65752 20334 65792
rect 20376 65752 20416 65792
rect 13228 65584 13268 65624
rect 8524 65500 8564 65540
rect 2764 65416 2804 65456
rect 11404 65416 11444 65456
rect 17932 65416 17972 65456
rect 10540 65332 10580 65372
rect 4300 65248 4340 65288
rect 6124 65164 6164 65204
rect 3688 64996 3728 65036
rect 3770 64996 3810 65036
rect 3852 64996 3892 65036
rect 3934 64996 3974 65036
rect 4016 64996 4056 65036
rect 18808 64996 18848 65036
rect 18890 64996 18930 65036
rect 18972 64996 19012 65036
rect 19054 64996 19094 65036
rect 19136 64996 19176 65036
rect 10540 64828 10580 64868
rect 13804 64576 13844 64616
rect 14860 64576 14900 64616
rect 2956 64324 2996 64364
rect 3052 64240 3092 64280
rect 4928 64240 4968 64280
rect 5010 64240 5050 64280
rect 5092 64240 5132 64280
rect 5174 64240 5214 64280
rect 5256 64240 5296 64280
rect 7660 64240 7700 64280
rect 20048 64240 20088 64280
rect 20130 64240 20170 64280
rect 20212 64240 20252 64280
rect 20294 64240 20334 64280
rect 20376 64240 20416 64280
rect 8524 63988 8564 64028
rect 4204 63904 4244 63944
rect 9004 63904 9044 63944
rect 11308 63820 11348 63860
rect 15052 63820 15092 63860
rect 17932 63736 17972 63776
rect 18508 63736 18548 63776
rect 5548 63652 5588 63692
rect 3688 63484 3728 63524
rect 3770 63484 3810 63524
rect 3852 63484 3892 63524
rect 3934 63484 3974 63524
rect 4016 63484 4056 63524
rect 18808 63484 18848 63524
rect 18890 63484 18930 63524
rect 18972 63484 19012 63524
rect 19054 63484 19094 63524
rect 19136 63484 19176 63524
rect 5548 63316 5588 63356
rect 5836 63316 5876 63356
rect 9004 63148 9044 63188
rect 5548 63064 5588 63104
rect 6604 63064 6644 63104
rect 16108 63064 16148 63104
rect 18124 63064 18164 63104
rect 13804 62812 13844 62852
rect 14092 62812 14132 62852
rect 4928 62728 4968 62768
rect 5010 62728 5050 62768
rect 5092 62728 5132 62768
rect 5174 62728 5214 62768
rect 5256 62728 5296 62768
rect 6316 62728 6356 62768
rect 20048 62728 20088 62768
rect 20130 62728 20170 62768
rect 20212 62728 20252 62768
rect 20294 62728 20334 62768
rect 20376 62728 20416 62768
rect 14476 62560 14516 62600
rect 8332 62476 8372 62516
rect 1708 62392 1748 62432
rect 4204 62392 4244 62432
rect 7660 62392 7700 62432
rect 11212 62056 11252 62096
rect 3688 61972 3728 62012
rect 3770 61972 3810 62012
rect 3852 61972 3892 62012
rect 3934 61972 3974 62012
rect 4016 61972 4056 62012
rect 18808 61972 18848 62012
rect 18890 61972 18930 62012
rect 18972 61972 19012 62012
rect 19054 61972 19094 62012
rect 19136 61972 19176 62012
rect 16108 61888 16148 61928
rect 11980 61804 12020 61844
rect 17164 61804 17204 61844
rect 2764 61720 2804 61760
rect 7564 61720 7604 61760
rect 9772 61720 9812 61760
rect 15628 61720 15668 61760
rect 9004 61636 9044 61676
rect 3340 61552 3380 61592
rect 10444 61552 10484 61592
rect 18316 61552 18356 61592
rect 12460 61468 12500 61508
rect 16300 61468 16340 61508
rect 10924 61384 10964 61424
rect 16684 61384 16724 61424
rect 4928 61216 4968 61256
rect 5010 61216 5050 61256
rect 5092 61216 5132 61256
rect 5174 61216 5214 61256
rect 5256 61216 5296 61256
rect 20048 61216 20088 61256
rect 20130 61216 20170 61256
rect 20212 61216 20252 61256
rect 20294 61216 20334 61256
rect 20376 61216 20416 61256
rect 1132 61048 1172 61088
rect 11692 61048 11732 61088
rect 13804 60964 13844 61004
rect 2476 60880 2516 60920
rect 15628 60880 15668 60920
rect 9196 60796 9236 60836
rect 11212 60796 11252 60836
rect 3340 60712 3380 60752
rect 14380 60712 14420 60752
rect 18508 60712 18548 60752
rect 19372 60628 19412 60668
rect 3688 60460 3728 60500
rect 3770 60460 3810 60500
rect 3852 60460 3892 60500
rect 3934 60460 3974 60500
rect 4016 60460 4056 60500
rect 6796 60460 6836 60500
rect 18808 60460 18848 60500
rect 18890 60460 18930 60500
rect 18972 60460 19012 60500
rect 19054 60460 19094 60500
rect 19136 60460 19176 60500
rect 4396 60208 4436 60248
rect 15244 60124 15284 60164
rect 3148 60040 3188 60080
rect 6124 60040 6164 60080
rect 6700 60040 6740 60080
rect 8524 60040 8564 60080
rect 11980 59788 12020 59828
rect 4928 59704 4968 59744
rect 5010 59704 5050 59744
rect 5092 59704 5132 59744
rect 5174 59704 5214 59744
rect 5256 59704 5296 59744
rect 9484 59704 9524 59744
rect 14092 59704 14132 59744
rect 13420 59620 13460 59660
rect 3244 59536 3284 59576
rect 15244 59704 15284 59744
rect 20048 59704 20088 59744
rect 20130 59704 20170 59744
rect 20212 59704 20252 59744
rect 20294 59704 20334 59744
rect 20376 59704 20416 59744
rect 15916 59620 15956 59660
rect 16876 59536 16916 59576
rect 18700 59284 18740 59324
rect 4204 59200 4244 59240
rect 10060 59200 10100 59240
rect 11308 59200 11348 59240
rect 2956 59116 2996 59156
rect 3688 58948 3728 58988
rect 3770 58948 3810 58988
rect 3852 58948 3892 58988
rect 3934 58948 3974 58988
rect 4016 58948 4056 58988
rect 15916 58948 15956 58988
rect 18808 58948 18848 58988
rect 18890 58948 18930 58988
rect 18972 58948 19012 58988
rect 19054 58948 19094 58988
rect 19136 58948 19176 58988
rect 5644 58780 5684 58820
rect 13036 58780 13076 58820
rect 7852 58696 7892 58736
rect 2572 58528 2612 58568
rect 6316 58528 6356 58568
rect 7660 58528 7700 58568
rect 7948 58528 7988 58568
rect 11404 58528 11444 58568
rect 11788 58528 11828 58568
rect 12748 58528 12788 58568
rect 16684 58528 16724 58568
rect 18028 58528 18068 58568
rect 3244 58444 3284 58484
rect 2860 58276 2900 58316
rect 4928 58192 4968 58232
rect 5010 58192 5050 58232
rect 5092 58192 5132 58232
rect 5174 58192 5214 58232
rect 5256 58192 5296 58232
rect 20048 58192 20088 58232
rect 20130 58192 20170 58232
rect 20212 58192 20252 58232
rect 20294 58192 20334 58232
rect 20376 58192 20416 58232
rect 18220 58024 18260 58064
rect 16108 57940 16148 57980
rect 5356 57772 5396 57812
rect 9484 57688 9524 57728
rect 9964 57520 10004 57560
rect 3688 57436 3728 57476
rect 3770 57436 3810 57476
rect 3852 57436 3892 57476
rect 3934 57436 3974 57476
rect 4016 57436 4056 57476
rect 12268 57436 12308 57476
rect 18808 57436 18848 57476
rect 18890 57436 18930 57476
rect 18972 57436 19012 57476
rect 19054 57436 19094 57476
rect 19136 57436 19176 57476
rect 4492 57352 4532 57392
rect 8140 57268 8180 57308
rect 13132 57268 13172 57308
rect 20812 57184 20852 57224
rect 8140 57100 8180 57140
rect 10060 57100 10100 57140
rect 14188 57100 14228 57140
rect 17452 57100 17492 57140
rect 2476 57016 2516 57056
rect 16300 57016 16340 57056
rect 19372 56848 19412 56888
rect 19564 56848 19604 56888
rect 4928 56680 4968 56720
rect 5010 56680 5050 56720
rect 5092 56680 5132 56720
rect 5174 56680 5214 56720
rect 5256 56680 5296 56720
rect 8332 56680 8372 56720
rect 13420 56680 13460 56720
rect 17644 56680 17684 56720
rect 20048 56680 20088 56720
rect 20130 56680 20170 56720
rect 20212 56680 20252 56720
rect 20294 56680 20334 56720
rect 20376 56680 20416 56720
rect 17452 56596 17492 56636
rect 4396 56512 4436 56552
rect 2764 56344 2804 56384
rect 5836 56344 5876 56384
rect 10924 56428 10964 56468
rect 17260 56512 17300 56552
rect 19372 56512 19412 56552
rect 10540 56344 10580 56384
rect 7756 56260 7796 56300
rect 3532 56176 3572 56216
rect 8332 56176 8372 56216
rect 14188 56260 14228 56300
rect 17356 56260 17396 56300
rect 2668 56092 2708 56132
rect 7660 56092 7700 56132
rect 11596 56008 11636 56048
rect 12460 56008 12500 56048
rect 3052 55924 3092 55964
rect 3688 55924 3728 55964
rect 3770 55924 3810 55964
rect 3852 55924 3892 55964
rect 3934 55924 3974 55964
rect 4016 55924 4056 55964
rect 18808 55924 18848 55964
rect 18890 55924 18930 55964
rect 18972 55924 19012 55964
rect 19054 55924 19094 55964
rect 19136 55924 19176 55964
rect 4108 55756 4148 55796
rect 16684 55756 16724 55796
rect 7756 55588 7796 55628
rect 14860 55588 14900 55628
rect 7660 55420 7700 55460
rect 10156 55504 10196 55544
rect 13420 55504 13460 55544
rect 14860 55420 14900 55460
rect 18700 55420 18740 55460
rect 19468 55420 19508 55460
rect 4928 55168 4968 55208
rect 5010 55168 5050 55208
rect 5092 55168 5132 55208
rect 5174 55168 5214 55208
rect 5256 55168 5296 55208
rect 15916 55168 15956 55208
rect 20048 55168 20088 55208
rect 20130 55168 20170 55208
rect 20212 55168 20252 55208
rect 20294 55168 20334 55208
rect 20376 55168 20416 55208
rect 6604 55084 6644 55124
rect 19660 55084 19700 55124
rect 15820 55000 15860 55040
rect 14188 54916 14228 54956
rect 1996 54748 2036 54788
rect 4108 54748 4148 54788
rect 9004 54748 9044 54788
rect 18220 54748 18260 54788
rect 10060 54664 10100 54704
rect 10828 54580 10868 54620
rect 11692 54580 11732 54620
rect 16684 54580 16724 54620
rect 2764 54496 2804 54536
rect 3688 54412 3728 54452
rect 3770 54412 3810 54452
rect 3852 54412 3892 54452
rect 3934 54412 3974 54452
rect 4016 54412 4056 54452
rect 11404 54412 11444 54452
rect 15244 54412 15284 54452
rect 18808 54412 18848 54452
rect 18890 54412 18930 54452
rect 18972 54412 19012 54452
rect 19054 54412 19094 54452
rect 19136 54412 19176 54452
rect 3532 54328 3572 54368
rect 1036 54160 1076 54200
rect 3532 54160 3572 54200
rect 5740 54160 5780 54200
rect 9004 54244 9044 54284
rect 9484 54244 9524 54284
rect 10924 54160 10964 54200
rect 12940 54160 12980 54200
rect 21388 54160 21428 54200
rect 10156 54076 10196 54116
rect 14188 53908 14228 53948
rect 14572 53908 14612 53948
rect 17452 54076 17492 54116
rect 17644 53992 17684 54032
rect 19948 53992 19988 54032
rect 16876 53908 16916 53948
rect 8524 53824 8564 53864
rect 9772 53740 9812 53780
rect 13228 53740 13268 53780
rect 4928 53656 4968 53696
rect 5010 53656 5050 53696
rect 5092 53656 5132 53696
rect 5174 53656 5214 53696
rect 5256 53656 5296 53696
rect 5356 53656 5396 53696
rect 15916 53656 15956 53696
rect 9196 53572 9236 53612
rect 17260 53740 17300 53780
rect 17356 53656 17396 53696
rect 20048 53656 20088 53696
rect 20130 53656 20170 53696
rect 20212 53656 20252 53696
rect 20294 53656 20334 53696
rect 20376 53656 20416 53696
rect 10540 53572 10580 53612
rect 19372 53572 19412 53612
rect 19852 53572 19892 53612
rect 12940 53488 12980 53528
rect 21292 53404 21332 53444
rect 3244 53320 3284 53360
rect 18028 53320 18068 53360
rect 7276 53236 7316 53276
rect 10540 53236 10580 53276
rect 17452 53236 17492 53276
rect 16300 53152 16340 53192
rect 19948 53152 19988 53192
rect 20140 53152 20180 53192
rect 8140 53068 8180 53108
rect 11692 53068 11732 53108
rect 13036 52984 13076 53024
rect 18028 52984 18068 53024
rect 3688 52900 3728 52940
rect 3770 52900 3810 52940
rect 3852 52900 3892 52940
rect 3934 52900 3974 52940
rect 4016 52900 4056 52940
rect 10156 52900 10196 52940
rect 18700 52984 18740 53024
rect 10540 52900 10580 52940
rect 18808 52900 18848 52940
rect 18890 52900 18930 52940
rect 18972 52900 19012 52940
rect 19054 52900 19094 52940
rect 19136 52900 19176 52940
rect 2572 52816 2612 52856
rect 5932 52816 5972 52856
rect 16108 52816 16148 52856
rect 11404 52732 11444 52772
rect 19948 52816 19988 52856
rect 14188 52564 14228 52604
rect 5548 52480 5588 52520
rect 2284 52396 2324 52436
rect 9004 52312 9044 52352
rect 10924 52312 10964 52352
rect 11788 52396 11828 52436
rect 14572 52396 14612 52436
rect 19372 52396 19412 52436
rect 20812 52312 20852 52352
rect 4928 52144 4968 52184
rect 5010 52144 5050 52184
rect 5092 52144 5132 52184
rect 5174 52144 5214 52184
rect 5256 52144 5296 52184
rect 16876 52144 16916 52184
rect 3052 52060 3092 52100
rect 10540 52060 10580 52100
rect 16300 52060 16340 52100
rect 17932 52144 17972 52184
rect 19948 52144 19988 52184
rect 20048 52144 20088 52184
rect 20130 52144 20170 52184
rect 20212 52144 20252 52184
rect 20294 52144 20334 52184
rect 20376 52144 20416 52184
rect 13132 51976 13172 52016
rect 19660 51976 19700 52016
rect 3436 51808 3476 51848
rect 4300 51808 4340 51848
rect 17644 51808 17684 51848
rect 12844 51724 12884 51764
rect 14860 51724 14900 51764
rect 5452 51640 5492 51680
rect 16108 51640 16148 51680
rect 18028 51640 18068 51680
rect 19276 51640 19316 51680
rect 5548 51556 5588 51596
rect 10732 51556 10772 51596
rect 16300 51556 16340 51596
rect 17260 51556 17300 51596
rect 13036 51472 13076 51512
rect 3688 51388 3728 51428
rect 3770 51388 3810 51428
rect 3852 51388 3892 51428
rect 3934 51388 3974 51428
rect 4016 51388 4056 51428
rect 11596 51388 11636 51428
rect 18808 51388 18848 51428
rect 18890 51388 18930 51428
rect 18972 51388 19012 51428
rect 19054 51388 19094 51428
rect 19136 51388 19176 51428
rect 7276 51304 7316 51344
rect 3148 51220 3188 51260
rect 7660 51220 7700 51260
rect 8044 51220 8084 51260
rect 8332 51220 8372 51260
rect 7852 51136 7892 51176
rect 8524 51136 8564 51176
rect 16108 51052 16148 51092
rect 8044 50800 8084 50840
rect 9772 50800 9812 50840
rect 8332 50716 8372 50756
rect 12172 50716 12212 50756
rect 19276 50968 19316 51008
rect 19852 50884 19892 50924
rect 17068 50800 17108 50840
rect 19948 50800 19988 50840
rect 4928 50632 4968 50672
rect 5010 50632 5050 50672
rect 5092 50632 5132 50672
rect 5174 50632 5214 50672
rect 5256 50632 5296 50672
rect 15724 50632 15764 50672
rect 19852 50632 19892 50672
rect 20048 50632 20088 50672
rect 20130 50632 20170 50672
rect 20212 50632 20252 50672
rect 20294 50632 20334 50672
rect 20376 50632 20416 50672
rect 13228 50548 13268 50588
rect 9004 50380 9044 50420
rect 19948 50380 19988 50420
rect 4300 50296 4340 50336
rect 4492 50296 4532 50336
rect 3148 50212 3188 50252
rect 20812 50128 20852 50168
rect 12172 50044 12212 50084
rect 19660 50044 19700 50084
rect 3148 49960 3188 50000
rect 5836 49960 5876 50000
rect 3688 49876 3728 49916
rect 3770 49876 3810 49916
rect 3852 49876 3892 49916
rect 3934 49876 3974 49916
rect 4016 49876 4056 49916
rect 18808 49876 18848 49916
rect 18890 49876 18930 49916
rect 18972 49876 19012 49916
rect 19054 49876 19094 49916
rect 19136 49876 19176 49916
rect 7372 49792 7412 49832
rect 19564 49792 19604 49832
rect 5356 49708 5396 49748
rect 5836 49708 5876 49748
rect 15340 49708 15380 49748
rect 7660 49624 7700 49664
rect 8332 49624 8372 49664
rect 4588 49540 4628 49580
rect 18316 49456 18356 49496
rect 2092 49372 2132 49412
rect 4108 49372 4148 49412
rect 4780 49372 4820 49412
rect 11500 49372 11540 49412
rect 10156 49288 10196 49328
rect 19948 49288 19988 49328
rect 5932 49204 5972 49244
rect 4928 49120 4968 49160
rect 5010 49120 5050 49160
rect 5092 49120 5132 49160
rect 5174 49120 5214 49160
rect 5256 49120 5296 49160
rect 20048 49120 20088 49160
rect 20130 49120 20170 49160
rect 20212 49120 20252 49160
rect 20294 49120 20334 49160
rect 20376 49120 20416 49160
rect 2572 48700 2612 48740
rect 17932 48952 17972 48992
rect 11500 48868 11540 48908
rect 19372 48868 19412 48908
rect 20812 48868 20852 48908
rect 16492 48616 16532 48656
rect 12556 48532 12596 48572
rect 2860 48448 2900 48488
rect 6604 48448 6644 48488
rect 12844 48448 12884 48488
rect 16492 48448 16532 48488
rect 21292 48448 21332 48488
rect 3688 48364 3728 48404
rect 3770 48364 3810 48404
rect 3852 48364 3892 48404
rect 3934 48364 3974 48404
rect 4016 48364 4056 48404
rect 5932 48364 5972 48404
rect 8524 48364 8564 48404
rect 14860 48364 14900 48404
rect 18808 48364 18848 48404
rect 18890 48364 18930 48404
rect 18972 48364 19012 48404
rect 19054 48364 19094 48404
rect 19136 48364 19176 48404
rect 2860 48196 2900 48236
rect 19468 48028 19508 48068
rect 8236 47860 8276 47900
rect 8524 47860 8564 47900
rect 14284 47860 14324 47900
rect 1996 47608 2036 47648
rect 3148 47608 3188 47648
rect 4928 47608 4968 47648
rect 5010 47608 5050 47648
rect 5092 47608 5132 47648
rect 5174 47608 5214 47648
rect 5256 47608 5296 47648
rect 20048 47608 20088 47648
rect 20130 47608 20170 47648
rect 20212 47608 20252 47648
rect 20294 47608 20334 47648
rect 20376 47608 20416 47648
rect 9580 47524 9620 47564
rect 18316 47524 18356 47564
rect 9196 47440 9236 47480
rect 10828 47440 10868 47480
rect 15724 47356 15764 47396
rect 4588 47272 4628 47312
rect 8524 47272 8564 47312
rect 10636 47104 10676 47144
rect 13420 46936 13460 46976
rect 3688 46852 3728 46892
rect 3770 46852 3810 46892
rect 3852 46852 3892 46892
rect 3934 46852 3974 46892
rect 4016 46852 4056 46892
rect 6604 46852 6644 46892
rect 18124 46852 18164 46892
rect 18808 46852 18848 46892
rect 18890 46852 18930 46892
rect 18972 46852 19012 46892
rect 19054 46852 19094 46892
rect 19136 46852 19176 46892
rect 9580 46768 9620 46808
rect 18028 46684 18068 46724
rect 7084 46600 7124 46640
rect 8140 46600 8180 46640
rect 9196 46600 9236 46640
rect 5836 46516 5876 46556
rect 4684 46432 4724 46472
rect 18700 46432 18740 46472
rect 19948 46432 19988 46472
rect 4588 46348 4628 46388
rect 20716 46348 20756 46388
rect 4492 46264 4532 46304
rect 18124 46264 18164 46304
rect 21388 46264 21428 46304
rect 4928 46096 4968 46136
rect 5010 46096 5050 46136
rect 5092 46096 5132 46136
rect 5174 46096 5214 46136
rect 5256 46096 5296 46136
rect 20048 46096 20088 46136
rect 20130 46096 20170 46136
rect 20212 46096 20252 46136
rect 20294 46096 20334 46136
rect 20376 46096 20416 46136
rect 4588 45928 4628 45968
rect 5836 45844 5876 45884
rect 6604 45844 6644 45884
rect 7852 45844 7892 45884
rect 9580 45760 9620 45800
rect 4588 45676 4628 45716
rect 5932 45676 5972 45716
rect 7084 45424 7124 45464
rect 16108 45760 16148 45800
rect 17452 45676 17492 45716
rect 3688 45340 3728 45380
rect 3770 45340 3810 45380
rect 3852 45340 3892 45380
rect 3934 45340 3974 45380
rect 4016 45340 4056 45380
rect 19852 45424 19892 45464
rect 18808 45340 18848 45380
rect 18890 45340 18930 45380
rect 18972 45340 19012 45380
rect 19054 45340 19094 45380
rect 19136 45340 19176 45380
rect 13708 45256 13748 45296
rect 15052 45256 15092 45296
rect 7660 45172 7700 45212
rect 11404 45172 11444 45212
rect 19852 45172 19892 45212
rect 2764 45088 2804 45128
rect 4684 45088 4724 45128
rect 4780 45004 4820 45044
rect 7276 44920 7316 44960
rect 4492 44836 4532 44876
rect 8908 44836 8948 44876
rect 7852 44752 7892 44792
rect 8140 44752 8180 44792
rect 19276 44668 19316 44708
rect 4928 44584 4968 44624
rect 5010 44584 5050 44624
rect 5092 44584 5132 44624
rect 5174 44584 5214 44624
rect 5256 44584 5296 44624
rect 9484 44584 9524 44624
rect 20048 44584 20088 44624
rect 20130 44584 20170 44624
rect 20212 44584 20252 44624
rect 20294 44584 20334 44624
rect 20376 44584 20416 44624
rect 4588 44416 4628 44456
rect 18700 44416 18740 44456
rect 4396 44332 4436 44372
rect 5356 44248 5396 44288
rect 15052 44164 15092 44204
rect 2284 44080 2324 44120
rect 8332 44080 8372 44120
rect 3688 43828 3728 43868
rect 3770 43828 3810 43868
rect 3852 43828 3892 43868
rect 3934 43828 3974 43868
rect 4016 43828 4056 43868
rect 18808 43828 18848 43868
rect 18890 43828 18930 43868
rect 18972 43828 19012 43868
rect 19054 43828 19094 43868
rect 19136 43828 19176 43868
rect 4300 43576 4340 43616
rect 4928 43072 4968 43112
rect 5010 43072 5050 43112
rect 5092 43072 5132 43112
rect 5174 43072 5214 43112
rect 5256 43072 5296 43112
rect 20048 43072 20088 43112
rect 20130 43072 20170 43112
rect 20212 43072 20252 43112
rect 20294 43072 20334 43112
rect 20376 43072 20416 43112
rect 748 42988 788 43028
rect 10348 42820 10388 42860
rect 15724 42820 15764 42860
rect 6604 42736 6644 42776
rect 10732 42736 10772 42776
rect 12652 42736 12692 42776
rect 11980 42568 12020 42608
rect 3688 42316 3728 42356
rect 3770 42316 3810 42356
rect 3852 42316 3892 42356
rect 3934 42316 3974 42356
rect 4016 42316 4056 42356
rect 18808 42316 18848 42356
rect 18890 42316 18930 42356
rect 18972 42316 19012 42356
rect 19054 42316 19094 42356
rect 19136 42316 19176 42356
rect 11596 42232 11636 42272
rect 10732 42064 10772 42104
rect 10156 41896 10196 41936
rect 11020 41896 11060 41936
rect 3532 41560 3572 41600
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 11980 41560 12020 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 2188 41476 2228 41516
rect 13996 41476 14036 41516
rect 14860 41476 14900 41516
rect 1804 41224 1844 41264
rect 9868 41224 9908 41264
rect 14092 41224 14132 41264
rect 364 40972 404 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 14476 40720 14516 40760
rect 14764 40720 14804 40760
rect 556 40636 596 40676
rect 13804 40636 13844 40676
rect 5548 40552 5588 40592
rect 8908 40384 8948 40424
rect 14860 40384 14900 40424
rect 1804 40300 1844 40340
rect 1996 40300 2036 40340
rect 10924 40300 10964 40340
rect 13804 40300 13844 40340
rect 4684 40216 4724 40256
rect 8332 40216 8372 40256
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 1804 39796 1844 39836
rect 10540 39712 10580 39752
rect 9004 39628 9044 39668
rect 12940 39628 12980 39668
rect 16492 39628 16532 39668
rect 14092 39544 14132 39584
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 5932 39208 5972 39248
rect 844 39124 884 39164
rect 6028 39124 6068 39164
rect 4780 39040 4820 39080
rect 14956 38872 14996 38912
rect 16396 38872 16436 38912
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 10732 38368 10772 38408
rect 11980 38452 12020 38492
rect 12748 38284 12788 38324
rect 3148 38200 3188 38240
rect 10252 38200 10292 38240
rect 11116 38200 11156 38240
rect 13324 38200 13364 38240
rect 14764 38200 14804 38240
rect 10636 38116 10676 38156
rect 14092 38116 14132 38156
rect 18316 38116 18356 38156
rect 19852 38116 19892 38156
rect 4300 38032 4340 38072
rect 11980 37948 12020 37988
rect 19564 37948 19604 37988
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 12748 37780 12788 37820
rect 15820 37864 15860 37904
rect 15148 37780 15188 37820
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 12748 37612 12788 37652
rect 15148 37612 15188 37652
rect 7276 37360 7316 37400
rect 12268 37276 12308 37316
rect 1900 37192 1940 37232
rect 4108 37192 4148 37232
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 1516 36940 1556 36980
rect 5644 36940 5684 36980
rect 6604 36940 6644 36980
rect 7084 36856 7124 36896
rect 5644 36772 5684 36812
rect 1132 36688 1172 36728
rect 9772 36688 9812 36728
rect 12748 36604 12788 36644
rect 10060 36520 10100 36560
rect 10732 36520 10772 36560
rect 13228 36520 13268 36560
rect 940 36436 980 36476
rect 6220 36436 6260 36476
rect 13036 36436 13076 36476
rect 15820 36436 15860 36476
rect 10828 36352 10868 36392
rect 19660 36352 19700 36392
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 11788 36268 11828 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 19468 36268 19508 36308
rect 6604 36184 6644 36224
rect 4300 36100 4340 36140
rect 7180 36100 7220 36140
rect 9676 36100 9716 36140
rect 19852 36100 19892 36140
rect 12652 36016 12692 36056
rect 17356 36016 17396 36056
rect 9100 35848 9140 35888
rect 748 35764 788 35804
rect 9484 35764 9524 35804
rect 10828 35764 10868 35804
rect 18316 35680 18356 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 6220 35428 6260 35468
rect 7276 35344 7316 35384
rect 20716 35344 20756 35384
rect 5836 35260 5876 35300
rect 7084 35260 7124 35300
rect 16108 35260 16148 35300
rect 16684 35260 16724 35300
rect 18316 35260 18356 35300
rect 2956 35176 2996 35216
rect 3148 35092 3188 35132
rect 18028 35092 18068 35132
rect 2764 35008 2804 35048
rect 4492 35008 4532 35048
rect 5836 35008 5876 35048
rect 8236 35008 8276 35048
rect 15052 35008 15092 35048
rect 19660 35008 19700 35048
rect 19948 35008 19988 35048
rect 3532 34924 3572 34964
rect 5548 34924 5588 34964
rect 11404 34924 11444 34964
rect 15340 34840 15380 34880
rect 1708 34756 1748 34796
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 5356 34756 5396 34796
rect 10348 34756 10388 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 5548 34672 5588 34712
rect 6604 34672 6644 34712
rect 2380 34588 2420 34628
rect 11788 34588 11828 34628
rect 13132 34588 13172 34628
rect 5548 34504 5588 34544
rect 6028 34504 6068 34544
rect 17452 34504 17492 34544
rect 6220 34420 6260 34460
rect 11116 34420 11156 34460
rect 1324 34336 1364 34376
rect 10732 34336 10772 34376
rect 12844 34336 12884 34376
rect 7660 34252 7700 34292
rect 12364 34168 12404 34208
rect 19852 34168 19892 34208
rect 2860 34084 2900 34124
rect 1324 34000 1364 34040
rect 2092 34000 2132 34040
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 10348 33916 10388 33956
rect 20716 33916 20756 33956
rect 3244 33832 3284 33872
rect 19948 33832 19988 33872
rect 8140 33748 8180 33788
rect 18124 33748 18164 33788
rect 3436 33664 3476 33704
rect 10828 33664 10868 33704
rect 18700 33664 18740 33704
rect 21388 33664 21428 33704
rect 4300 33580 4340 33620
rect 16588 33580 16628 33620
rect 1228 33496 1268 33536
rect 6220 33496 6260 33536
rect 17260 33496 17300 33536
rect 5836 33412 5876 33452
rect 13324 33328 13364 33368
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 16876 33244 16916 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 21388 33160 21428 33200
rect 4684 33076 4724 33116
rect 3244 32992 3284 33032
rect 15052 32992 15092 33032
rect 16588 32992 16628 33032
rect 17452 32992 17492 33032
rect 1612 32908 1652 32948
rect 17932 32992 17972 33032
rect 2572 32824 2612 32864
rect 14092 32824 14132 32864
rect 1132 32740 1172 32780
rect 17452 32740 17492 32780
rect 3244 32656 3284 32696
rect 13420 32656 13460 32696
rect 17644 32656 17684 32696
rect 18220 32656 18260 32696
rect 2860 32572 2900 32612
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 4108 32320 4148 32360
rect 13420 32320 13460 32360
rect 20716 32320 20756 32360
rect 16972 32236 17012 32276
rect 18700 32236 18740 32276
rect 2860 32152 2900 32192
rect 18220 32152 18260 32192
rect 2956 32068 2996 32108
rect 19852 31984 19892 32024
rect 4780 31900 4820 31940
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 4684 31648 4724 31688
rect 13132 31480 13172 31520
rect 18124 31396 18164 31436
rect 5356 31312 5396 31352
rect 13996 31312 14036 31352
rect 14764 31312 14804 31352
rect 5644 31144 5684 31184
rect 2860 31060 2900 31100
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 5548 30976 5588 31016
rect 17068 30976 17108 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 13804 30892 13844 30932
rect 12268 30808 12308 30848
rect 2476 30640 2516 30680
rect 3532 30640 3572 30680
rect 5836 30640 5876 30680
rect 18028 30640 18068 30680
rect 5548 30556 5588 30596
rect 9676 30556 9716 30596
rect 12844 30556 12884 30596
rect 7276 30472 7316 30512
rect 20620 30304 20660 30344
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 11020 30220 11060 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 5452 30136 5492 30176
rect 7660 30052 7700 30092
rect 20716 30052 20756 30092
rect 5644 29884 5684 29924
rect 9676 29800 9716 29840
rect 17452 29884 17492 29924
rect 17068 29800 17108 29840
rect 13612 29716 13652 29756
rect 6028 29632 6068 29672
rect 14380 29632 14420 29672
rect 2284 29464 2324 29504
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 6220 29464 6260 29504
rect 2284 29296 2324 29336
rect 10828 29296 10868 29336
rect 17260 29716 17300 29756
rect 16972 29632 17012 29672
rect 19372 29632 19412 29672
rect 17644 29548 17684 29588
rect 18316 29548 18356 29588
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 14860 29296 14900 29336
rect 19276 29212 19316 29252
rect 19468 29212 19508 29252
rect 8236 29128 8276 29168
rect 10828 28876 10868 28916
rect 556 28792 596 28832
rect 2476 28792 2516 28832
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 19564 28624 19604 28664
rect 20620 28540 20660 28580
rect 10732 28372 10772 28412
rect 3244 28288 3284 28328
rect 4492 28288 4532 28328
rect 13996 28288 14036 28328
rect 16300 28288 16340 28328
rect 17260 28288 17300 28328
rect 19756 28204 19796 28244
rect 20716 28204 20756 28244
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 6028 27784 6068 27824
rect 15340 27784 15380 27824
rect 3532 27700 3572 27740
rect 6988 27700 7028 27740
rect 1324 27616 1364 27656
rect 6604 27616 6644 27656
rect 7084 27616 7124 27656
rect 12268 27616 12308 27656
rect 18316 27616 18356 27656
rect 4108 27532 4148 27572
rect 19468 27532 19508 27572
rect 21004 27448 21044 27488
rect 11404 27364 11444 27404
rect 1996 27280 2036 27320
rect 2476 27280 2516 27320
rect 11116 27280 11156 27320
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 16876 27196 16916 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 8236 27112 8276 27152
rect 15052 27112 15092 27152
rect 14860 27028 14900 27068
rect 17452 27028 17492 27068
rect 16972 26860 17012 26900
rect 2476 26776 2516 26816
rect 5644 26776 5684 26816
rect 2284 26440 2324 26480
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 13420 26440 13460 26480
rect 13708 26440 13748 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 9196 26356 9236 26396
rect 1420 26272 1460 26312
rect 7084 26188 7124 26228
rect 268 26104 308 26144
rect 19756 26104 19796 26144
rect 3532 26020 3572 26060
rect 16300 26020 16340 26060
rect 4588 25936 4628 25976
rect 8044 25936 8084 25976
rect 16684 25936 16724 25976
rect 17068 25936 17108 25976
rect 20524 25936 20564 25976
rect 19564 25852 19604 25892
rect 5932 25768 5972 25808
rect 7468 25768 7508 25808
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 18700 25684 18740 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 13036 25600 13076 25640
rect 16876 25600 16916 25640
rect 17452 25600 17492 25640
rect 19276 25600 19316 25640
rect 14860 25432 14900 25472
rect 5452 25180 5492 25220
rect 5356 25096 5396 25136
rect 13420 25264 13460 25304
rect 14092 25264 14132 25304
rect 18604 25180 18644 25220
rect 18796 25180 18836 25220
rect 18124 25012 18164 25052
rect 20908 25012 20948 25052
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 6988 24928 7028 24968
rect 15340 24928 15380 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 13036 24844 13076 24884
rect 19564 24760 19604 24800
rect 2476 24676 2516 24716
rect 6604 24676 6644 24716
rect 2956 24592 2996 24632
rect 5356 24592 5396 24632
rect 7372 24592 7412 24632
rect 8236 24592 8276 24632
rect 9292 24592 9332 24632
rect 10156 24592 10196 24632
rect 19276 24592 19316 24632
rect 4780 24508 4820 24548
rect 13996 24508 14036 24548
rect 20908 24508 20948 24548
rect 9964 24424 10004 24464
rect 6028 24340 6068 24380
rect 21196 24340 21236 24380
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 5836 24172 5876 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 9868 24004 9908 24044
rect 10732 24004 10772 24044
rect 9100 23920 9140 23960
rect 14092 23920 14132 23960
rect 18700 23920 18740 23960
rect 4108 23500 4148 23540
rect 7372 23836 7412 23876
rect 11020 23752 11060 23792
rect 17068 23752 17108 23792
rect 7372 23668 7412 23708
rect 12268 23668 12308 23708
rect 11308 23584 11348 23624
rect 19372 23584 19412 23624
rect 13132 23500 13172 23540
rect 172 23416 212 23456
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 7564 23332 7604 23372
rect 11308 23332 11348 23372
rect 19372 23248 19412 23288
rect 4588 23164 4628 23204
rect 7372 23164 7412 23204
rect 16492 23164 16532 23204
rect 17356 23164 17396 23204
rect 11116 23080 11156 23120
rect 17452 22996 17492 23036
rect 13036 22912 13076 22952
rect 19660 22828 19700 22868
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 14764 22660 14804 22700
rect 18604 22660 18644 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 9580 22576 9620 22616
rect 15820 22492 15860 22532
rect 7372 22324 7412 22364
rect 16396 22324 16436 22364
rect 16876 22324 16916 22364
rect 2380 22240 2420 22280
rect 2668 22240 2708 22280
rect 14092 22240 14132 22280
rect 16876 22156 16916 22196
rect 7084 22072 7124 22112
rect 7372 22072 7412 22112
rect 13132 22072 13172 22112
rect 3244 21988 3284 22028
rect 6988 21988 7028 22028
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 16972 21904 17012 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 6700 21820 6740 21860
rect 2956 21736 2996 21776
rect 9580 21652 9620 21692
rect 15340 21652 15380 21692
rect 1228 21400 1268 21440
rect 5644 21568 5684 21608
rect 7468 21568 7508 21608
rect 17644 21568 17684 21608
rect 20620 21568 20660 21608
rect 14380 21484 14420 21524
rect 21004 21484 21044 21524
rect 7564 21316 7604 21356
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 15820 21148 15860 21188
rect 18508 21148 18548 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 14188 20980 14228 21020
rect 19276 20980 19316 21020
rect 4108 20896 4148 20936
rect 9676 20728 9716 20768
rect 10732 20728 10772 20768
rect 11308 20728 11348 20768
rect 9964 20560 10004 20600
rect 2572 20476 2612 20516
rect 4108 20392 4148 20432
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 16300 20392 16340 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 17260 20308 17300 20348
rect 19564 20308 19604 20348
rect 6028 20224 6068 20264
rect 13036 20224 13076 20264
rect 17068 20224 17108 20264
rect 19276 20224 19316 20264
rect 10444 20140 10484 20180
rect 17260 20140 17300 20180
rect 2092 20056 2132 20096
rect 9676 20056 9716 20096
rect 16588 20056 16628 20096
rect 10828 19972 10868 20012
rect 11308 19972 11348 20012
rect 16396 19888 16436 19928
rect 16300 19804 16340 19844
rect 19948 19804 19988 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 10348 19636 10388 19676
rect 16588 19636 16628 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 6028 19468 6068 19508
rect 20812 19468 20852 19508
rect 11212 19384 11252 19424
rect 2572 19300 2612 19340
rect 7564 19216 7604 19256
rect 10444 19216 10484 19256
rect 5452 19132 5492 19172
rect 7468 19132 7508 19172
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 14476 18880 14516 18920
rect 15916 18880 15956 18920
rect 16300 18880 16340 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 21100 18880 21140 18920
rect 12268 18796 12308 18836
rect 1228 18712 1268 18752
rect 11116 18712 11156 18752
rect 20524 18712 20564 18752
rect 21004 18712 21044 18752
rect 14092 18628 14132 18668
rect 3724 18544 3764 18584
rect 6412 18544 6452 18584
rect 6604 18544 6644 18584
rect 8044 18544 8084 18584
rect 13708 18544 13748 18584
rect 20524 18544 20564 18584
rect 21004 18544 21044 18584
rect 7948 18460 7988 18500
rect 2572 18376 2612 18416
rect 10348 18376 10388 18416
rect 17068 18376 17108 18416
rect 14476 18292 14516 18332
rect 20524 18292 20564 18332
rect 15148 18208 15188 18248
rect 3244 18124 3284 18164
rect 1228 18040 1268 18080
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 16396 18124 16436 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 1516 18040 1556 18080
rect 13708 18040 13748 18080
rect 6412 17956 6452 17996
rect 19468 18040 19508 18080
rect 8236 17956 8276 17996
rect 17452 17956 17492 17996
rect 76 17872 116 17912
rect 15340 17872 15380 17912
rect 16492 17872 16532 17912
rect 2572 17788 2612 17828
rect 2764 17788 2804 17828
rect 9580 17788 9620 17828
rect 17260 17788 17300 17828
rect 5068 17704 5108 17744
rect 6412 17704 6452 17744
rect 7660 17620 7700 17660
rect 11788 17620 11828 17660
rect 7180 17536 7220 17576
rect 7948 17452 7988 17492
rect 10828 17452 10868 17492
rect 4204 17368 4244 17408
rect 4780 17368 4820 17408
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 8716 17368 8756 17408
rect 9580 17368 9620 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 2572 17284 2612 17324
rect 6412 17284 6452 17324
rect 7372 17284 7412 17324
rect 20620 17284 20660 17324
rect 9868 17200 9908 17240
rect 13708 17200 13748 17240
rect 2572 17116 2612 17156
rect 7564 17116 7604 17156
rect 13228 17116 13268 17156
rect 6220 17032 6260 17072
rect 7180 17032 7220 17072
rect 16684 17032 16724 17072
rect 19660 16948 19700 16988
rect 940 16696 980 16736
rect 3244 16696 3284 16736
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 15724 16780 15764 16820
rect 18508 16780 18548 16820
rect 7660 16696 7700 16736
rect 11404 16696 11444 16736
rect 13324 16696 13364 16736
rect 18700 16696 18740 16736
rect 13804 16612 13844 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 4204 16528 4244 16568
rect 16300 16528 16340 16568
rect 4876 16360 4916 16400
rect 9388 16360 9428 16400
rect 19276 16360 19316 16400
rect 21100 16276 21140 16316
rect 11020 16192 11060 16232
rect 15916 16192 15956 16232
rect 21004 16192 21044 16232
rect 4108 16024 4148 16064
rect 13036 16024 13076 16064
rect 1900 15940 1940 15980
rect 4492 15940 4532 15980
rect 18028 15940 18068 15980
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 16300 15688 16340 15728
rect 16780 15688 16820 15728
rect 1228 15604 1268 15644
rect 1900 15520 1940 15560
rect 20140 15520 20180 15560
rect 16396 15352 16436 15392
rect 18220 15352 18260 15392
rect 16492 15268 16532 15308
rect 18508 15184 18548 15224
rect 20812 15184 20852 15224
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 3244 14848 3284 14888
rect 7948 14848 7988 14888
rect 8812 14848 8852 14888
rect 5740 14764 5780 14804
rect 3244 14680 3284 14720
rect 4204 14680 4244 14720
rect 11500 14596 11540 14636
rect 12076 14596 12116 14636
rect 18508 14680 18548 14720
rect 15148 14512 15188 14552
rect 6124 14428 6164 14468
rect 19564 14428 19604 14468
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 15724 14344 15764 14384
rect 17068 14344 17108 14384
rect 19852 14344 19892 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 3532 14008 3572 14048
rect 6124 14008 6164 14048
rect 4108 13924 4148 13964
rect 11500 13840 11540 13880
rect 15724 13840 15764 13880
rect 18028 13840 18068 13880
rect 4204 13756 4244 13796
rect 19276 13756 19316 13796
rect 13996 13672 14036 13712
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 5452 13588 5492 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 8812 13504 8852 13544
rect 17260 13504 17300 13544
rect 172 13420 212 13460
rect 7756 13336 7796 13376
rect 14860 13420 14900 13460
rect 4300 13252 4340 13292
rect 19948 13252 19988 13292
rect 4396 13168 4436 13208
rect 5644 13168 5684 13208
rect 6604 13168 6644 13208
rect 14572 13084 14612 13124
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 3052 12664 3092 12704
rect 7372 12664 7412 12704
rect 3532 12580 3572 12620
rect 5452 12580 5492 12620
rect 10156 12580 10196 12620
rect 3244 12496 3284 12536
rect 3820 12496 3860 12536
rect 6220 12496 6260 12536
rect 8428 12496 8468 12536
rect 4780 12412 4820 12452
rect 16204 12328 16244 12368
rect 7276 12160 7316 12200
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 16684 12076 16724 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 1228 11992 1268 12032
rect 12172 11992 12212 12032
rect 3244 11908 3284 11948
rect 4204 11908 4244 11948
rect 21196 11824 21236 11864
rect 13228 11740 13268 11780
rect 16204 11656 16244 11696
rect 17260 11656 17300 11696
rect 6316 11404 6356 11444
rect 7948 11404 7988 11444
rect 13804 11404 13844 11444
rect 16396 11404 16436 11444
rect 16876 11404 16916 11444
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 13228 11320 13268 11360
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 9388 11236 9428 11276
rect 12844 11236 12884 11276
rect 13036 11236 13076 11276
rect 16396 11236 16436 11276
rect 13804 11152 13844 11192
rect 20140 11152 20180 11192
rect 4108 11068 4148 11108
rect 8428 11068 8468 11108
rect 12076 11068 12116 11108
rect 4684 10984 4724 11024
rect 9580 10984 9620 11024
rect 17260 10816 17300 10856
rect 268 10732 308 10772
rect 4108 10732 4148 10772
rect 11788 10732 11828 10772
rect 1516 10648 1556 10688
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18028 10480 18068 10520
rect 18508 10480 18548 10520
rect 6124 10396 6164 10436
rect 18220 10396 18260 10436
rect 17932 10312 17972 10352
rect 4108 10228 4148 10268
rect 9964 10228 10004 10268
rect 3436 10060 3476 10100
rect 4204 9976 4244 10016
rect 18700 9976 18740 10016
rect 20524 9892 20564 9932
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 8812 9808 8852 9848
rect 13996 9808 14036 9848
rect 17932 9808 17972 9848
rect 19468 9808 19508 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 20812 9808 20852 9848
rect 8524 9724 8564 9764
rect 18028 9724 18068 9764
rect 1612 9472 1652 9512
rect 4396 9472 4436 9512
rect 16204 9472 16244 9512
rect 17452 9472 17492 9512
rect 19372 9472 19407 9512
rect 19407 9472 19412 9512
rect 19564 9472 19604 9512
rect 2572 9304 2612 9344
rect 4300 9304 4340 9344
rect 6220 9304 6260 9344
rect 2860 9220 2900 9260
rect 3628 9220 3635 9260
rect 3635 9220 3668 9260
rect 4492 9220 4532 9260
rect 7372 9220 7412 9260
rect 20524 9136 20564 9176
rect 20908 9136 20948 9176
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 6604 9052 6644 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 3436 8968 3476 9008
rect 3532 8884 3572 8924
rect 3724 8800 3764 8840
rect 6316 8800 6356 8840
rect 9388 8800 9428 8840
rect 20140 8800 20180 8840
rect 5644 8716 5684 8756
rect 19468 8632 19508 8672
rect 4108 8548 4148 8588
rect 9196 8548 9236 8588
rect 4492 8464 4532 8504
rect 12844 8380 12884 8420
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4780 7960 4820 8000
rect 7564 7960 7604 8000
rect 8236 7960 8276 8000
rect 9196 7960 9236 8000
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19276 7960 19316 8000
rect 7564 7708 7604 7748
rect 19372 7708 19412 7748
rect 13420 7624 13460 7664
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 4684 7456 4724 7496
rect 5356 7456 5396 7496
rect 76 7288 116 7328
rect 2572 7288 2612 7328
rect 7468 7120 7508 7160
rect 17164 7036 17204 7076
rect 20140 7120 20180 7160
rect 19276 6952 19316 6992
rect 19564 6952 19604 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 16396 6700 16436 6740
rect 17452 6700 17492 6740
rect 16396 6532 16436 6572
rect 19852 6112 19892 6152
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 19468 5440 19508 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 12364 5020 12404 5060
rect 20716 5020 20756 5060
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 9964 3676 10004 3716
rect 6220 3424 6260 3464
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 940 2836 980 2876
rect 13804 2668 13844 2708
rect 14380 2668 14420 2708
rect 460 2332 500 2372
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 17740 2248 17780 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 1036 2164 1076 2204
rect 5740 2080 5780 2120
rect 6508 2080 6548 2120
rect 6892 2080 6932 2120
rect 7276 2080 7316 2120
rect 13900 2080 13940 2120
rect 15436 2080 15476 2120
rect 16300 2080 16340 2120
rect 17548 2080 17588 2120
rect 18124 2080 18164 2120
rect 18316 2080 18356 2120
rect 18604 2080 18644 2120
rect 19564 2080 19604 2120
rect 8140 1828 8180 1868
rect 10540 1828 10580 1868
rect 10924 1828 10964 1868
rect 11692 1828 11732 1868
rect 11980 1828 12020 1868
rect 14284 1828 14324 1868
rect 14668 1828 14708 1868
rect 15532 1828 15572 1868
rect 16012 1828 16052 1868
rect 16396 1828 16436 1868
rect 15436 1744 15476 1784
rect 16588 1828 16628 1868
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 2956 1240 2996 1280
rect 3148 1240 3188 1280
rect 6796 1240 6836 1280
rect 9772 1240 9812 1280
rect 15436 1240 15476 1280
rect 15628 1240 15668 1280
rect 17836 1240 17876 1280
rect 18412 1240 18452 1280
rect 1804 1156 1844 1196
rect 11596 1156 11636 1196
rect 13036 1156 13076 1196
rect 13420 1156 13460 1196
rect 14956 1156 14996 1196
rect 16108 1156 16148 1196
rect 3340 1072 3380 1112
rect 12748 1072 12788 1112
rect 15532 1072 15572 1112
rect 9004 988 9044 1028
rect 10636 988 10676 1028
rect 19180 904 19220 944
rect 8332 820 8372 860
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 748 568 788 608
rect 9484 568 9524 608
rect 11884 400 11924 440
rect 10060 316 10100 356
rect 5068 232 5108 272
rect 4876 148 4916 188
rect 12940 148 12980 188
rect 3340 64 3380 104
rect 13516 64 13556 104
<< metal4 >>
rect 19083 85952 19125 85961
rect 19083 85912 19084 85952
rect 19124 85912 19125 85952
rect 19083 85903 19125 85912
rect 19276 85952 19316 85961
rect 19084 85818 19124 85903
rect 19276 85793 19316 85912
rect 19275 85784 19317 85793
rect 19275 85744 19276 85784
rect 19316 85744 19317 85784
rect 19275 85735 19317 85744
rect 6508 85616 6548 85625
rect 2380 85196 2420 85205
rect 1515 83516 1557 83525
rect 1515 83476 1516 83516
rect 1556 83476 1557 83516
rect 1515 83467 1557 83476
rect 2092 83516 2132 83525
rect 1516 83382 1556 83467
rect 76 77888 116 77897
rect 76 42701 116 77848
rect 1516 77216 1556 77225
rect 651 76544 693 76553
rect 651 76504 652 76544
rect 692 76504 693 76544
rect 651 76495 693 76504
rect 652 76410 692 76495
rect 268 75872 308 75881
rect 172 72512 212 72521
rect 75 42692 117 42701
rect 75 42652 76 42692
rect 116 42652 117 42692
rect 75 42643 117 42652
rect 172 40601 212 72472
rect 268 42785 308 75832
rect 364 71168 404 71177
rect 267 42776 309 42785
rect 267 42736 268 42776
rect 308 42736 309 42776
rect 267 42727 309 42736
rect 364 41012 404 71128
rect 364 40963 404 40972
rect 556 69152 596 69161
rect 556 40676 596 69112
rect 748 68480 788 68489
rect 748 43028 788 68440
rect 1036 67136 1076 67145
rect 1036 59921 1076 67096
rect 1228 65792 1268 65801
rect 1132 61088 1172 61097
rect 1035 59912 1077 59921
rect 1035 59872 1036 59912
rect 1076 59872 1077 59912
rect 1035 59863 1077 59872
rect 748 42979 788 42988
rect 1036 54200 1076 54209
rect 556 40627 596 40636
rect 171 40592 213 40601
rect 171 40552 172 40592
rect 212 40552 213 40592
rect 171 40543 213 40552
rect 844 39164 884 39173
rect 748 35804 788 35813
rect 459 34208 501 34217
rect 459 34168 460 34208
rect 500 34168 501 34208
rect 459 34159 501 34168
rect 268 26144 308 26153
rect 172 23456 212 23465
rect 76 17912 116 17921
rect 76 7328 116 17872
rect 172 13460 212 23416
rect 172 13411 212 13420
rect 268 10772 308 26104
rect 268 10723 308 10732
rect 76 7279 116 7288
rect 460 2372 500 34159
rect 555 33704 597 33713
rect 555 33664 556 33704
rect 596 33664 597 33704
rect 555 33655 597 33664
rect 556 28832 596 33655
rect 748 29000 788 35764
rect 556 28783 596 28792
rect 652 28960 788 29000
rect 652 26480 692 28960
rect 556 26440 692 26480
rect 556 22121 596 26440
rect 844 22280 884 39124
rect 652 22240 884 22280
rect 940 36476 980 36485
rect 555 22112 597 22121
rect 555 22072 556 22112
rect 596 22072 597 22112
rect 555 22063 597 22072
rect 652 16409 692 22240
rect 747 22112 789 22121
rect 747 22072 748 22112
rect 788 22072 789 22112
rect 747 22063 789 22072
rect 651 16400 693 16409
rect 651 16360 652 16400
rect 692 16360 693 16400
rect 651 16351 693 16360
rect 460 2323 500 2332
rect 748 608 788 22063
rect 940 20180 980 36436
rect 844 20140 980 20180
rect 844 11360 884 20140
rect 939 16820 981 16829
rect 939 16780 940 16820
rect 980 16780 981 16820
rect 939 16771 981 16780
rect 940 16736 980 16771
rect 940 16685 980 16696
rect 844 11320 980 11360
rect 940 2876 980 11320
rect 940 2827 980 2836
rect 1036 2204 1076 54160
rect 1132 36728 1172 61048
rect 1132 36679 1172 36688
rect 1228 33704 1268 65752
rect 1516 36980 1556 77176
rect 1804 75200 1844 75209
rect 1516 36931 1556 36940
rect 1708 62432 1748 62441
rect 1708 34796 1748 62392
rect 1804 41264 1844 75160
rect 1804 40340 1844 41224
rect 1804 40291 1844 40300
rect 1900 71840 1940 71849
rect 1708 34747 1748 34756
rect 1804 39836 1844 39845
rect 1323 34376 1365 34385
rect 1323 34336 1324 34376
rect 1364 34336 1365 34376
rect 1323 34327 1365 34336
rect 1324 34040 1364 34327
rect 1324 33991 1364 34000
rect 1132 33664 1268 33704
rect 1132 32780 1172 33664
rect 1227 33536 1269 33545
rect 1227 33496 1228 33536
rect 1268 33496 1269 33536
rect 1227 33487 1269 33496
rect 1228 33402 1268 33487
rect 1132 32731 1172 32740
rect 1612 32948 1652 32957
rect 1324 27656 1364 27665
rect 1324 26153 1364 27616
rect 1419 26312 1461 26321
rect 1419 26272 1420 26312
rect 1460 26272 1461 26312
rect 1419 26263 1461 26272
rect 1420 26178 1460 26263
rect 1323 26144 1365 26153
rect 1323 26104 1324 26144
rect 1364 26104 1365 26144
rect 1323 26095 1365 26104
rect 1227 21440 1269 21449
rect 1227 21400 1228 21440
rect 1268 21400 1269 21440
rect 1227 21391 1269 21400
rect 1228 21306 1268 21391
rect 1227 18752 1269 18761
rect 1227 18712 1228 18752
rect 1268 18712 1269 18752
rect 1227 18703 1269 18712
rect 1228 18618 1268 18703
rect 1227 18332 1269 18341
rect 1227 18292 1228 18332
rect 1268 18292 1269 18332
rect 1227 18283 1269 18292
rect 1228 18080 1268 18283
rect 1228 18031 1268 18040
rect 1516 18080 1556 18089
rect 1228 15644 1268 15653
rect 1228 12032 1268 15604
rect 1228 11983 1268 11992
rect 1516 10688 1556 18040
rect 1516 10639 1556 10648
rect 1612 9512 1652 32908
rect 1612 9463 1652 9472
rect 1036 2155 1076 2164
rect 1804 1196 1844 39796
rect 1900 37232 1940 71800
rect 1996 54788 2036 54797
rect 1996 47648 2036 54748
rect 2092 49412 2132 83476
rect 2284 83516 2324 83525
rect 2092 49363 2132 49372
rect 2188 69824 2228 69833
rect 1996 47599 2036 47608
rect 2188 41516 2228 69784
rect 2284 52436 2324 83476
rect 2284 52387 2324 52396
rect 2380 45977 2420 85156
rect 3688 84692 4056 84701
rect 3728 84652 3770 84692
rect 3810 84652 3852 84692
rect 3892 84652 3934 84692
rect 3974 84652 4016 84692
rect 3688 84643 4056 84652
rect 5836 84440 5876 84449
rect 4928 83936 5296 83945
rect 4968 83896 5010 83936
rect 5050 83896 5092 83936
rect 5132 83896 5174 83936
rect 5214 83896 5256 83936
rect 4928 83887 5296 83896
rect 2668 83348 2708 83357
rect 2476 60920 2516 60929
rect 2476 57056 2516 60880
rect 2476 57007 2516 57016
rect 2572 58568 2612 58577
rect 2572 52856 2612 58528
rect 2668 56132 2708 83308
rect 3688 83180 4056 83189
rect 3728 83140 3770 83180
rect 3810 83140 3852 83180
rect 3892 83140 3934 83180
rect 3974 83140 4016 83180
rect 3688 83131 4056 83140
rect 2860 82844 2900 82853
rect 2764 65456 2804 65465
rect 2764 61760 2804 65416
rect 2764 61711 2804 61720
rect 2860 58316 2900 82804
rect 3244 82844 3284 82853
rect 3244 81920 3284 82804
rect 3532 82844 3572 82853
rect 3244 81880 3476 81920
rect 2956 64364 2996 64373
rect 2956 64280 2996 64324
rect 3052 64280 3092 64289
rect 2956 64240 3052 64280
rect 3052 64231 3092 64240
rect 3340 61592 3380 61601
rect 3340 60752 3380 61552
rect 3148 60080 3188 60089
rect 2860 58267 2900 58276
rect 2956 59156 2996 59165
rect 2668 56083 2708 56092
rect 2764 56384 2804 56393
rect 2572 52807 2612 52816
rect 2764 54536 2804 56344
rect 2572 48740 2612 48749
rect 2379 45968 2421 45977
rect 2379 45928 2380 45968
rect 2420 45928 2421 45968
rect 2379 45919 2421 45928
rect 2188 41467 2228 41476
rect 2284 44120 2324 44129
rect 1900 37183 1940 37192
rect 1996 40340 2036 40349
rect 1996 27320 2036 40300
rect 1996 27271 2036 27280
rect 2092 34040 2132 34049
rect 2092 20096 2132 34000
rect 2284 29504 2324 44080
rect 2284 29455 2324 29464
rect 2380 34628 2420 34637
rect 2284 29336 2324 29345
rect 2284 26480 2324 29296
rect 2284 26431 2324 26440
rect 2380 22280 2420 34588
rect 2572 32864 2612 48700
rect 2764 45128 2804 54496
rect 2859 52016 2901 52025
rect 2859 51976 2860 52016
rect 2900 51976 2901 52016
rect 2859 51967 2901 51976
rect 2860 48488 2900 51967
rect 2956 51764 2996 59116
rect 3052 55964 3092 55973
rect 3052 52100 3092 55924
rect 3052 51848 3092 52060
rect 3148 52025 3188 60040
rect 3244 59576 3284 59585
rect 3244 58484 3284 59536
rect 3244 53360 3284 58444
rect 3147 52016 3189 52025
rect 3147 51976 3148 52016
rect 3188 51976 3189 52016
rect 3147 51967 3189 51976
rect 3052 51808 3188 51848
rect 2956 51724 3092 51764
rect 2860 48236 2900 48448
rect 2860 48187 2900 48196
rect 2764 45079 2804 45088
rect 2956 35216 2996 35225
rect 2572 32815 2612 32824
rect 2764 35048 2804 35057
rect 2476 30680 2516 30689
rect 2476 28832 2516 30640
rect 2476 28783 2516 28792
rect 2476 27320 2516 27329
rect 2476 26816 2516 27280
rect 2476 24716 2516 26776
rect 2476 24667 2516 24676
rect 2380 22231 2420 22240
rect 2668 22280 2708 22289
rect 2092 20047 2132 20056
rect 2572 20516 2612 20525
rect 2572 19340 2612 20476
rect 2572 19291 2612 19300
rect 2572 18416 2612 18425
rect 2572 17828 2612 18376
rect 2572 17779 2612 17788
rect 2572 17324 2612 17333
rect 2572 17156 2612 17284
rect 2572 17107 2612 17116
rect 1900 15980 1940 15989
rect 1900 15560 1940 15940
rect 1900 15511 1940 15520
rect 2572 9344 2612 9353
rect 2572 7328 2612 9304
rect 2668 8849 2708 22240
rect 2764 17828 2804 35008
rect 2860 34124 2900 34133
rect 2860 32612 2900 34084
rect 2860 32192 2900 32572
rect 2860 32143 2900 32152
rect 2956 32108 2996 35176
rect 2956 32059 2996 32068
rect 2764 17779 2804 17788
rect 2860 31100 2900 31109
rect 2860 9260 2900 31060
rect 2956 24632 2996 24641
rect 2956 21776 2996 24592
rect 2956 21727 2996 21736
rect 2955 16400 2997 16409
rect 2955 16360 2956 16400
rect 2996 16360 2997 16400
rect 2955 16351 2997 16360
rect 2860 9211 2900 9220
rect 2667 8840 2709 8849
rect 2667 8800 2668 8840
rect 2708 8800 2709 8840
rect 2667 8791 2709 8800
rect 2572 7279 2612 7288
rect 2956 1280 2996 16351
rect 3052 12704 3092 51724
rect 3148 51260 3188 51808
rect 3148 51211 3188 51220
rect 3148 50252 3188 50261
rect 3148 50000 3188 50212
rect 3148 47648 3188 49960
rect 3148 38240 3188 47608
rect 3148 38191 3188 38200
rect 3052 12655 3092 12664
rect 3148 35132 3188 35141
rect 2956 1231 2996 1240
rect 3148 1280 3188 35092
rect 3244 33872 3284 53320
rect 3244 33823 3284 33832
rect 3244 33032 3284 33041
rect 3244 32696 3284 32992
rect 3244 32647 3284 32656
rect 3244 28328 3284 28337
rect 3244 22028 3284 28288
rect 3244 21979 3284 21988
rect 3244 18164 3284 18173
rect 3244 16736 3284 18124
rect 3244 16687 3284 16696
rect 3244 14888 3284 14897
rect 3244 14720 3284 14848
rect 3244 14671 3284 14680
rect 3244 12536 3284 12545
rect 3244 11948 3284 12496
rect 3244 11899 3284 11908
rect 3148 1231 3188 1240
rect 1804 1147 1844 1156
rect 3340 1112 3380 60712
rect 3436 57905 3476 81880
rect 3435 57896 3477 57905
rect 3435 57856 3436 57896
rect 3476 57856 3477 57896
rect 3435 57847 3477 57856
rect 3532 56897 3572 82804
rect 4928 82424 5296 82433
rect 4968 82384 5010 82424
rect 5050 82384 5092 82424
rect 5132 82384 5174 82424
rect 5214 82384 5256 82424
rect 4928 82375 5296 82384
rect 3688 81668 4056 81677
rect 3728 81628 3770 81668
rect 3810 81628 3852 81668
rect 3892 81628 3934 81668
rect 3974 81628 4016 81668
rect 3688 81619 4056 81628
rect 4928 80912 5296 80921
rect 4968 80872 5010 80912
rect 5050 80872 5092 80912
rect 5132 80872 5174 80912
rect 5214 80872 5256 80912
rect 4928 80863 5296 80872
rect 3688 80156 4056 80165
rect 3728 80116 3770 80156
rect 3810 80116 3852 80156
rect 3892 80116 3934 80156
rect 3974 80116 4016 80156
rect 3688 80107 4056 80116
rect 4928 79400 5296 79409
rect 4968 79360 5010 79400
rect 5050 79360 5092 79400
rect 5132 79360 5174 79400
rect 5214 79360 5256 79400
rect 4928 79351 5296 79360
rect 3688 78644 4056 78653
rect 3728 78604 3770 78644
rect 3810 78604 3852 78644
rect 3892 78604 3934 78644
rect 3974 78604 4016 78644
rect 3688 78595 4056 78604
rect 4928 77888 5296 77897
rect 4968 77848 5010 77888
rect 5050 77848 5092 77888
rect 5132 77848 5174 77888
rect 5214 77848 5256 77888
rect 4928 77839 5296 77848
rect 3688 77132 4056 77141
rect 3728 77092 3770 77132
rect 3810 77092 3852 77132
rect 3892 77092 3934 77132
rect 3974 77092 4016 77132
rect 3688 77083 4056 77092
rect 4928 76376 5296 76385
rect 4968 76336 5010 76376
rect 5050 76336 5092 76376
rect 5132 76336 5174 76376
rect 5214 76336 5256 76376
rect 4928 76327 5296 76336
rect 3688 75620 4056 75629
rect 3728 75580 3770 75620
rect 3810 75580 3852 75620
rect 3892 75580 3934 75620
rect 3974 75580 4016 75620
rect 3688 75571 4056 75580
rect 4928 74864 5296 74873
rect 4968 74824 5010 74864
rect 5050 74824 5092 74864
rect 5132 74824 5174 74864
rect 5214 74824 5256 74864
rect 4928 74815 5296 74824
rect 3688 74108 4056 74117
rect 3728 74068 3770 74108
rect 3810 74068 3852 74108
rect 3892 74068 3934 74108
rect 3974 74068 4016 74108
rect 3688 74059 4056 74068
rect 5356 73856 5396 73865
rect 4928 73352 5296 73361
rect 4968 73312 5010 73352
rect 5050 73312 5092 73352
rect 5132 73312 5174 73352
rect 5214 73312 5256 73352
rect 4928 73303 5296 73312
rect 3688 72596 4056 72605
rect 3728 72556 3770 72596
rect 3810 72556 3852 72596
rect 3892 72556 3934 72596
rect 3974 72556 4016 72596
rect 3688 72547 4056 72556
rect 4300 72260 4340 72269
rect 3688 71084 4056 71093
rect 3728 71044 3770 71084
rect 3810 71044 3852 71084
rect 3892 71044 3934 71084
rect 3974 71044 4016 71084
rect 3688 71035 4056 71044
rect 3688 69572 4056 69581
rect 3728 69532 3770 69572
rect 3810 69532 3852 69572
rect 3892 69532 3934 69572
rect 3974 69532 4016 69572
rect 3688 69523 4056 69532
rect 4108 69320 4148 69329
rect 4108 68396 4148 69280
rect 3688 68060 4056 68069
rect 3728 68020 3770 68060
rect 3810 68020 3852 68060
rect 3892 68020 3934 68060
rect 3974 68020 4016 68060
rect 3688 68011 4056 68020
rect 3688 66548 4056 66557
rect 3728 66508 3770 66548
rect 3810 66508 3852 66548
rect 3892 66508 3934 66548
rect 3974 66508 4016 66548
rect 3688 66499 4056 66508
rect 4108 66044 4148 68356
rect 4108 65995 4148 66004
rect 4300 65288 4340 72220
rect 4928 71840 5296 71849
rect 4968 71800 5010 71840
rect 5050 71800 5092 71840
rect 5132 71800 5174 71840
rect 5214 71800 5256 71840
rect 4928 71791 5296 71800
rect 5356 71588 5396 73816
rect 5356 71539 5396 71548
rect 5548 70664 5588 70673
rect 4492 70496 4532 70505
rect 4492 69152 4532 70456
rect 4928 70328 5296 70337
rect 4968 70288 5010 70328
rect 5050 70288 5092 70328
rect 5132 70288 5174 70328
rect 5214 70288 5256 70328
rect 4928 70279 5296 70288
rect 4492 69103 4532 69112
rect 4928 68816 5296 68825
rect 4968 68776 5010 68816
rect 5050 68776 5092 68816
rect 5132 68776 5174 68816
rect 5214 68776 5256 68816
rect 4928 68767 5296 68776
rect 5548 67556 5588 70624
rect 4928 67304 5296 67313
rect 4968 67264 5010 67304
rect 5050 67264 5092 67304
rect 5132 67264 5174 67304
rect 5214 67264 5256 67304
rect 4928 67255 5296 67264
rect 4300 65239 4340 65248
rect 4396 67052 4436 67061
rect 3688 65036 4056 65045
rect 3728 64996 3770 65036
rect 3810 64996 3852 65036
rect 3892 64996 3934 65036
rect 3974 64996 4016 65036
rect 3688 64987 4056 64996
rect 4204 63944 4244 63953
rect 3688 63524 4056 63533
rect 3728 63484 3770 63524
rect 3810 63484 3852 63524
rect 3892 63484 3934 63524
rect 3974 63484 4016 63524
rect 3688 63475 4056 63484
rect 4204 62432 4244 63904
rect 4204 62383 4244 62392
rect 3688 62012 4056 62021
rect 3728 61972 3770 62012
rect 3810 61972 3852 62012
rect 3892 61972 3934 62012
rect 3974 61972 4016 62012
rect 3688 61963 4056 61972
rect 3688 60500 4056 60509
rect 3728 60460 3770 60500
rect 3810 60460 3852 60500
rect 3892 60460 3934 60500
rect 3974 60460 4016 60500
rect 3688 60451 4056 60460
rect 4396 60248 4436 67012
rect 4928 65792 5296 65801
rect 4968 65752 5010 65792
rect 5050 65752 5092 65792
rect 5132 65752 5174 65792
rect 5214 65752 5256 65792
rect 4928 65743 5296 65752
rect 4928 64280 5296 64289
rect 4968 64240 5010 64280
rect 5050 64240 5092 64280
rect 5132 64240 5174 64280
rect 5214 64240 5256 64280
rect 4928 64231 5296 64240
rect 5548 63692 5588 67516
rect 5548 63356 5588 63652
rect 5548 63307 5588 63316
rect 5644 69152 5684 69161
rect 5548 63104 5588 63113
rect 5644 63104 5684 69112
rect 5836 64280 5876 84400
rect 6220 84440 6260 84449
rect 5588 63064 5684 63104
rect 5740 64240 5876 64280
rect 6028 73688 6068 73697
rect 4928 62768 5296 62777
rect 4968 62728 5010 62768
rect 5050 62728 5092 62768
rect 5132 62728 5174 62768
rect 5214 62728 5256 62768
rect 4928 62719 5296 62728
rect 4928 61256 5296 61265
rect 4968 61216 5010 61256
rect 5050 61216 5092 61256
rect 5132 61216 5174 61256
rect 5214 61216 5256 61256
rect 4928 61207 5296 61216
rect 4204 59240 4244 59249
rect 3688 58988 4056 58997
rect 3728 58948 3770 58988
rect 3810 58948 3852 58988
rect 3892 58948 3934 58988
rect 3974 58948 4016 58988
rect 3688 58939 4056 58948
rect 3688 57476 4056 57485
rect 3728 57436 3770 57476
rect 3810 57436 3852 57476
rect 3892 57436 3934 57476
rect 3974 57436 4016 57476
rect 3688 57427 4056 57436
rect 3531 56888 3573 56897
rect 3531 56848 3532 56888
rect 3572 56848 3573 56888
rect 3531 56839 3573 56848
rect 3532 56216 3572 56225
rect 3532 54368 3572 56176
rect 3688 55964 4056 55973
rect 3728 55924 3770 55964
rect 3810 55924 3852 55964
rect 3892 55924 3934 55964
rect 3974 55924 4016 55964
rect 3688 55915 4056 55924
rect 4108 55796 4148 55805
rect 4108 54788 4148 55756
rect 3688 54452 4056 54461
rect 3728 54412 3770 54452
rect 3810 54412 3852 54452
rect 3892 54412 3934 54452
rect 3974 54412 4016 54452
rect 3688 54403 4056 54412
rect 3436 54328 3532 54368
rect 3436 51848 3476 54328
rect 3532 54319 3572 54328
rect 3436 51799 3476 51808
rect 3532 54200 3572 54209
rect 3532 41600 3572 54160
rect 3688 52940 4056 52949
rect 3728 52900 3770 52940
rect 3810 52900 3852 52940
rect 3892 52900 3934 52940
rect 3974 52900 4016 52940
rect 3688 52891 4056 52900
rect 3688 51428 4056 51437
rect 3728 51388 3770 51428
rect 3810 51388 3852 51428
rect 3892 51388 3934 51428
rect 3974 51388 4016 51428
rect 3688 51379 4056 51388
rect 3688 49916 4056 49925
rect 3728 49876 3770 49916
rect 3810 49876 3852 49916
rect 3892 49876 3934 49916
rect 3974 49876 4016 49916
rect 3688 49867 4056 49876
rect 4108 49412 4148 54748
rect 4108 49363 4148 49372
rect 3688 48404 4056 48413
rect 3728 48364 3770 48404
rect 3810 48364 3852 48404
rect 3892 48364 3934 48404
rect 3974 48364 4016 48404
rect 3688 48355 4056 48364
rect 3688 46892 4056 46901
rect 3728 46852 3770 46892
rect 3810 46852 3852 46892
rect 3892 46852 3934 46892
rect 3974 46852 4016 46892
rect 3688 46843 4056 46852
rect 3688 45380 4056 45389
rect 3728 45340 3770 45380
rect 3810 45340 3852 45380
rect 3892 45340 3934 45380
rect 3974 45340 4016 45380
rect 3688 45331 4056 45340
rect 3688 43868 4056 43877
rect 3728 43828 3770 43868
rect 3810 43828 3852 43868
rect 3892 43828 3934 43868
rect 3974 43828 4016 43868
rect 3688 43819 4056 43828
rect 3688 42356 4056 42365
rect 3728 42316 3770 42356
rect 3810 42316 3852 42356
rect 3892 42316 3934 42356
rect 3974 42316 4016 42356
rect 3688 42307 4056 42316
rect 3532 41551 3572 41560
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 4108 37232 4148 37241
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 3532 34964 3572 34973
rect 3436 33704 3476 33713
rect 3436 12545 3476 33664
rect 3532 30680 3572 34924
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 4108 32360 4148 37192
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 3532 30631 3572 30640
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 3532 27740 3572 27749
rect 3532 26060 3572 27700
rect 4108 27572 4148 32320
rect 4108 27523 4148 27532
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 3532 26011 3572 26020
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 4108 23540 4148 23549
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 4108 20936 4148 23500
rect 4108 20432 4148 20896
rect 4108 20383 4148 20392
rect 4204 20180 4244 59200
rect 4396 56552 4436 60208
rect 4928 59744 5296 59753
rect 4968 59704 5010 59744
rect 5050 59704 5092 59744
rect 5132 59704 5174 59744
rect 5214 59704 5256 59744
rect 4928 59695 5296 59704
rect 4928 58232 5296 58241
rect 4968 58192 5010 58232
rect 5050 58192 5092 58232
rect 5132 58192 5174 58232
rect 5214 58192 5256 58232
rect 4928 58183 5296 58192
rect 5356 57812 5396 57821
rect 4299 51848 4341 51857
rect 4299 51808 4300 51848
rect 4340 51808 4341 51848
rect 4299 51799 4341 51808
rect 4300 51714 4340 51799
rect 4300 50336 4340 50345
rect 4300 43616 4340 50296
rect 4396 44372 4436 56512
rect 4492 57392 4532 57401
rect 4492 50336 4532 57352
rect 4928 56720 5296 56729
rect 4968 56680 5010 56720
rect 5050 56680 5092 56720
rect 5132 56680 5174 56720
rect 5214 56680 5256 56720
rect 4928 56671 5296 56680
rect 4928 55208 5296 55217
rect 4968 55168 5010 55208
rect 5050 55168 5092 55208
rect 5132 55168 5174 55208
rect 5214 55168 5256 55208
rect 4928 55159 5296 55168
rect 4928 53696 5296 53705
rect 4968 53656 5010 53696
rect 5050 53656 5092 53696
rect 5132 53656 5174 53696
rect 5214 53656 5256 53696
rect 4928 53647 5296 53656
rect 5356 53696 5396 57772
rect 5356 53647 5396 53656
rect 5548 52520 5588 63064
rect 4928 52184 5296 52193
rect 4968 52144 5010 52184
rect 5050 52144 5092 52184
rect 5132 52144 5174 52184
rect 5214 52144 5256 52184
rect 4928 52135 5296 52144
rect 5452 51680 5492 51689
rect 4928 50672 5296 50681
rect 4968 50632 5010 50672
rect 5050 50632 5092 50672
rect 5132 50632 5174 50672
rect 5214 50632 5256 50672
rect 4928 50623 5296 50632
rect 4492 50287 4532 50296
rect 5356 49748 5396 49757
rect 4588 49580 4628 49589
rect 4588 47312 4628 49540
rect 4588 47263 4628 47272
rect 4780 49412 4820 49421
rect 4684 46472 4724 46481
rect 4588 46388 4628 46397
rect 4492 46304 4532 46313
rect 4492 44876 4532 46264
rect 4588 45968 4628 46348
rect 4588 45919 4628 45928
rect 4587 45716 4629 45725
rect 4587 45676 4588 45716
rect 4628 45676 4629 45716
rect 4587 45667 4629 45676
rect 4588 45582 4628 45667
rect 4684 45128 4724 46432
rect 4492 44827 4532 44836
rect 4588 45088 4684 45128
rect 4588 44456 4628 45088
rect 4684 45079 4724 45088
rect 4780 45044 4820 49372
rect 4928 49160 5296 49169
rect 4968 49120 5010 49160
rect 5050 49120 5092 49160
rect 5132 49120 5174 49160
rect 5214 49120 5256 49160
rect 4928 49111 5296 49120
rect 4928 47648 5296 47657
rect 4968 47608 5010 47648
rect 5050 47608 5092 47648
rect 5132 47608 5174 47648
rect 5214 47608 5256 47648
rect 4928 47599 5296 47608
rect 4928 46136 5296 46145
rect 4968 46096 5010 46136
rect 5050 46096 5092 46136
rect 5132 46096 5174 46136
rect 5214 46096 5256 46136
rect 4928 46087 5296 46096
rect 4780 44995 4820 45004
rect 4683 44960 4725 44969
rect 4683 44920 4684 44960
rect 4724 44920 4725 44960
rect 4683 44911 4725 44920
rect 4588 44407 4628 44416
rect 4396 44323 4436 44332
rect 4300 43567 4340 43576
rect 4684 40256 4724 44911
rect 4928 44624 5296 44633
rect 4968 44584 5010 44624
rect 5050 44584 5092 44624
rect 5132 44584 5174 44624
rect 5214 44584 5256 44624
rect 4928 44575 5296 44584
rect 5356 44288 5396 49708
rect 5356 44239 5396 44248
rect 4928 43112 5296 43121
rect 4968 43072 5010 43112
rect 5050 43072 5092 43112
rect 5132 43072 5174 43112
rect 5214 43072 5256 43112
rect 4928 43063 5296 43072
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 4684 40207 4724 40216
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 4780 39080 4820 39089
rect 4300 38072 4340 38081
rect 4300 36140 4340 38032
rect 4300 36091 4340 36100
rect 4491 35048 4533 35057
rect 4491 35008 4492 35048
rect 4532 35008 4533 35048
rect 4491 34999 4533 35008
rect 4492 34914 4532 34999
rect 4300 33620 4340 33629
rect 4300 29000 4340 33580
rect 4684 33116 4724 33125
rect 4684 31688 4724 33076
rect 4780 31940 4820 39040
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 5355 35216 5397 35225
rect 5355 35176 5356 35216
rect 5396 35176 5397 35216
rect 5355 35167 5397 35176
rect 5356 34796 5396 35167
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 4780 31891 4820 31900
rect 4684 31639 4724 31648
rect 5356 31352 5396 34756
rect 5356 31303 5396 31312
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 5452 30176 5492 51640
rect 5548 51596 5588 52480
rect 5548 51547 5588 51556
rect 5644 58820 5684 58829
rect 5644 46640 5684 58780
rect 5740 54200 5780 64240
rect 5740 54151 5780 54160
rect 5836 63356 5876 63365
rect 5836 56384 5876 63316
rect 5836 50000 5876 56344
rect 5836 49748 5876 49960
rect 5836 49699 5876 49708
rect 5932 52856 5972 52865
rect 5932 49244 5972 52816
rect 5932 49195 5972 49204
rect 5932 48404 5972 48413
rect 5644 46600 5780 46640
rect 5547 40592 5589 40601
rect 5547 40552 5548 40592
rect 5588 40552 5589 40592
rect 5547 40543 5589 40552
rect 5548 40458 5588 40543
rect 5644 36980 5684 36989
rect 5644 36812 5684 36940
rect 5548 34964 5588 34973
rect 5548 34712 5588 34924
rect 5548 34663 5588 34672
rect 5548 34544 5588 34553
rect 5548 31016 5588 34504
rect 5548 30967 5588 30976
rect 5644 31184 5684 36772
rect 5452 30127 5492 30136
rect 5548 30596 5588 30605
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 4300 28960 4532 29000
rect 4108 20140 4244 20180
rect 4492 28328 4532 28960
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 3723 18584 3765 18593
rect 3723 18544 3724 18584
rect 3764 18544 3765 18584
rect 3723 18535 3765 18544
rect 3724 18450 3764 18535
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 4108 16064 4148 20140
rect 4204 17408 4244 17417
rect 4204 16568 4244 17368
rect 4204 16519 4244 16528
rect 4108 16015 4148 16024
rect 4492 15980 4532 28288
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 4588 25976 4628 25985
rect 4588 23204 4628 25936
rect 5452 25220 5492 25229
rect 5356 25136 5396 25145
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 5356 24632 5396 25096
rect 4588 23155 4628 23164
rect 4780 24548 4820 24557
rect 4780 17408 4820 24508
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 4928 20383 5296 20392
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 5067 17744 5109 17753
rect 5067 17704 5068 17744
rect 5108 17704 5109 17744
rect 5067 17695 5109 17704
rect 5068 17610 5108 17695
rect 4780 17359 4820 17368
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 4875 16400 4917 16409
rect 4875 16360 4876 16400
rect 4916 16360 4917 16400
rect 4875 16351 4917 16360
rect 4876 16266 4916 16351
rect 4492 15931 4532 15940
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 4204 14720 4244 14729
rect 3532 14048 3572 14057
rect 3532 12620 3572 14008
rect 4108 13964 4148 13973
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 3532 12571 3572 12580
rect 3435 12536 3477 12545
rect 3435 12496 3436 12536
rect 3476 12496 3477 12536
rect 3435 12487 3477 12496
rect 3819 12536 3861 12545
rect 3819 12496 3820 12536
rect 3860 12496 3861 12536
rect 3819 12487 3861 12496
rect 3820 12402 3860 12487
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 4108 11108 4148 13924
rect 4204 13796 4244 14680
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 4204 11948 4244 13756
rect 4204 11899 4244 11908
rect 4300 13292 4340 13301
rect 4108 11059 4148 11068
rect 4108 10772 4148 10781
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 4108 10268 4148 10732
rect 3436 10100 3476 10109
rect 3436 9008 3476 10060
rect 3628 9260 3668 9269
rect 3436 8959 3476 8968
rect 3532 9220 3628 9260
rect 3532 8924 3572 9220
rect 3628 9211 3668 9220
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3724 8933 3764 8935
rect 3532 8875 3572 8884
rect 3723 8924 3765 8933
rect 3723 8884 3724 8924
rect 3764 8884 3765 8924
rect 3723 8875 3765 8884
rect 3724 8840 3764 8875
rect 3724 8791 3764 8800
rect 4108 8588 4148 10228
rect 4204 10016 4244 10025
rect 4204 8933 4244 9976
rect 4300 9344 4340 13252
rect 4396 13208 4436 13217
rect 4396 9512 4436 13168
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 4780 12452 4820 12461
rect 4396 9463 4436 9472
rect 4684 11024 4724 11033
rect 4300 9295 4340 9304
rect 4492 9260 4532 9269
rect 4203 8924 4245 8933
rect 4203 8884 4204 8924
rect 4244 8884 4245 8924
rect 4203 8875 4245 8884
rect 4108 8539 4148 8548
rect 4492 8504 4532 9220
rect 4492 8455 4532 8464
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 4684 7496 4724 10984
rect 4780 8000 4820 12412
rect 4928 11360 5296 11369
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4780 7951 4820 7960
rect 4684 7447 4724 7456
rect 5356 7496 5396 24592
rect 5452 19172 5492 25180
rect 5452 19123 5492 19132
rect 5452 13628 5492 13637
rect 5452 12620 5492 13588
rect 5452 12571 5492 12580
rect 5548 10025 5588 30556
rect 5644 29924 5684 31144
rect 5644 29875 5684 29884
rect 5644 26816 5684 26825
rect 5644 21608 5684 26776
rect 5644 21559 5684 21568
rect 5740 14804 5780 46600
rect 5836 46556 5876 46565
rect 5836 45884 5876 46516
rect 5836 45835 5876 45844
rect 5932 45716 5972 48364
rect 5932 45667 5972 45676
rect 5932 39248 5972 39257
rect 5836 35300 5876 35309
rect 5836 35225 5876 35260
rect 5835 35216 5877 35225
rect 5835 35176 5836 35216
rect 5876 35176 5877 35216
rect 5835 35167 5877 35176
rect 5836 35165 5876 35167
rect 5836 35048 5876 35057
rect 5836 33452 5876 35008
rect 5836 33403 5876 33412
rect 5836 30680 5876 30689
rect 5836 24212 5876 30640
rect 5932 26321 5972 39208
rect 6028 39164 6068 73648
rect 6124 66968 6164 66977
rect 6124 65204 6164 66928
rect 6124 65155 6164 65164
rect 6028 39115 6068 39124
rect 6124 60080 6164 60089
rect 6028 34544 6068 34553
rect 6028 29672 6068 34504
rect 6028 29623 6068 29632
rect 6028 27824 6068 27833
rect 5931 26312 5973 26321
rect 5931 26272 5932 26312
rect 5972 26272 5973 26312
rect 5931 26263 5973 26272
rect 5932 25808 5972 26263
rect 5932 25759 5972 25768
rect 6028 24380 6068 27784
rect 6028 24331 6068 24340
rect 5836 24163 5876 24172
rect 6028 20264 6068 20273
rect 6028 19508 6068 20224
rect 6028 19459 6068 19468
rect 5740 14755 5780 14764
rect 6124 14468 6164 60040
rect 6220 36476 6260 84400
rect 6412 73856 6452 73865
rect 6316 67136 6356 67145
rect 6316 62768 6356 67096
rect 6316 62719 6356 62728
rect 6220 36427 6260 36436
rect 6316 58568 6356 58577
rect 6220 35468 6260 35477
rect 6220 34460 6260 35428
rect 6220 34411 6260 34420
rect 6220 33536 6260 33545
rect 6220 29504 6260 33496
rect 6220 29455 6260 29464
rect 6124 14419 6164 14428
rect 6220 17072 6260 17081
rect 6124 14048 6164 14057
rect 5644 13208 5684 13217
rect 5547 10016 5589 10025
rect 5547 9976 5548 10016
rect 5588 9976 5589 10016
rect 5547 9967 5589 9976
rect 5644 8756 5684 13168
rect 6124 10436 6164 14008
rect 6124 10387 6164 10396
rect 6220 12536 6260 17032
rect 6316 16829 6356 58528
rect 6412 18584 6452 73816
rect 6412 17996 6452 18544
rect 6412 17947 6452 17956
rect 6412 17744 6452 17753
rect 6412 17324 6452 17704
rect 6412 17275 6452 17284
rect 6315 16820 6357 16829
rect 6315 16780 6316 16820
rect 6356 16780 6357 16820
rect 6315 16771 6357 16780
rect 5644 8707 5684 8716
rect 6220 9344 6260 12496
rect 5356 7447 5396 7456
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 6220 3464 6260 9304
rect 6316 11444 6356 11453
rect 6316 8840 6356 11404
rect 6316 8791 6356 8800
rect 6220 3415 6260 3424
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 5739 2120 5781 2129
rect 5739 2080 5740 2120
rect 5780 2080 5781 2120
rect 5739 2071 5781 2080
rect 6508 2120 6548 85576
rect 16012 85616 16052 85625
rect 13900 84608 13940 84617
rect 6892 84524 6932 84533
rect 6795 84440 6837 84449
rect 6795 84400 6796 84440
rect 6836 84400 6837 84440
rect 6795 84391 6837 84400
rect 6796 84306 6836 84391
rect 6604 69992 6644 70001
rect 6604 67388 6644 69952
rect 6796 68396 6836 68405
rect 6796 68069 6836 68356
rect 6795 68060 6837 68069
rect 6795 68020 6796 68060
rect 6836 68020 6837 68060
rect 6795 68011 6837 68020
rect 6604 63104 6644 67348
rect 6604 63055 6644 63064
rect 6796 60500 6836 60509
rect 6700 60080 6740 60089
rect 6604 55124 6644 55133
rect 6604 48488 6644 55084
rect 6604 48439 6644 48448
rect 6604 46892 6644 46901
rect 6604 45884 6644 46852
rect 6604 45835 6644 45844
rect 6603 42776 6645 42785
rect 6603 42736 6604 42776
rect 6644 42736 6645 42776
rect 6603 42727 6645 42736
rect 6604 42642 6644 42727
rect 6604 36980 6644 36989
rect 6604 36224 6644 36940
rect 6604 34712 6644 36184
rect 6604 27656 6644 34672
rect 6604 27607 6644 27616
rect 6604 24716 6644 24725
rect 6604 18584 6644 24676
rect 6700 21860 6740 60040
rect 6700 21811 6740 21820
rect 6604 18535 6644 18544
rect 6604 13208 6644 13217
rect 6604 9092 6644 13168
rect 6604 9043 6644 9052
rect 6508 2071 6548 2080
rect 5740 1986 5780 2071
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 6796 1280 6836 60460
rect 6892 2120 6932 84484
rect 10636 84440 10676 84449
rect 8908 84356 8948 84365
rect 7180 83516 7220 83525
rect 6988 83180 7028 83189
rect 6988 27740 7028 83140
rect 7084 46640 7124 46649
rect 7084 45464 7124 46600
rect 7084 45415 7124 45424
rect 7084 36896 7124 36905
rect 7084 35300 7124 36856
rect 7180 36140 7220 83476
rect 7372 83516 7412 83525
rect 7275 53276 7317 53285
rect 7275 53236 7276 53276
rect 7316 53236 7317 53276
rect 7275 53227 7317 53236
rect 7276 53142 7316 53227
rect 7276 51344 7316 51353
rect 7276 44960 7316 51304
rect 7372 49832 7412 83476
rect 8140 83516 8180 83525
rect 7660 64280 7700 64289
rect 7660 62432 7700 64240
rect 7372 49783 7412 49792
rect 7564 61760 7604 61769
rect 7276 44911 7316 44920
rect 7180 36091 7220 36100
rect 7276 37400 7316 37409
rect 7276 35384 7316 37360
rect 7276 35335 7316 35344
rect 7084 35251 7124 35260
rect 7564 34217 7604 61720
rect 7660 58568 7700 62392
rect 7660 58519 7700 58528
rect 7852 58736 7892 58745
rect 7756 56300 7796 56309
rect 7660 56132 7700 56141
rect 7660 55460 7700 56092
rect 7756 55628 7796 56260
rect 7756 55579 7796 55588
rect 7852 55460 7892 58696
rect 7948 58568 7988 58577
rect 7948 57989 7988 58528
rect 7947 57980 7989 57989
rect 7947 57940 7948 57980
rect 7988 57940 7989 57980
rect 7947 57931 7989 57940
rect 7660 55411 7700 55420
rect 7756 55420 7892 55460
rect 7660 51260 7700 51269
rect 7660 49664 7700 51220
rect 7660 45212 7700 49624
rect 7660 45163 7700 45172
rect 7660 34292 7700 34301
rect 7563 34208 7605 34217
rect 7563 34168 7564 34208
rect 7604 34168 7605 34208
rect 7563 34159 7605 34168
rect 6988 27691 7028 27700
rect 7276 30512 7316 30521
rect 7084 27656 7124 27665
rect 7084 26228 7124 27616
rect 6988 24968 7028 24977
rect 6988 22028 7028 24928
rect 7084 22112 7124 26188
rect 7084 22063 7124 22072
rect 6988 21979 7028 21988
rect 7180 17576 7220 17585
rect 7180 17072 7220 17536
rect 7180 17023 7220 17032
rect 7276 12200 7316 30472
rect 7660 30092 7700 34252
rect 7660 30043 7700 30052
rect 7468 25808 7508 25817
rect 7372 24632 7412 24641
rect 7372 23876 7412 24592
rect 7372 23708 7412 23836
rect 7372 23659 7412 23668
rect 7372 23204 7412 23213
rect 7372 22364 7412 23164
rect 7372 22315 7412 22324
rect 7372 22112 7412 22121
rect 7372 17324 7412 22072
rect 7468 21608 7508 25768
rect 7468 21559 7508 21568
rect 7564 23372 7604 23381
rect 7564 21356 7604 23332
rect 7564 21307 7604 21316
rect 7564 19256 7604 19265
rect 7372 17275 7412 17284
rect 7468 19172 7508 19181
rect 7276 12151 7316 12160
rect 7372 12704 7412 12713
rect 7372 9260 7412 12664
rect 7372 9211 7412 9220
rect 7468 7160 7508 19132
rect 7564 17156 7604 19216
rect 7564 17107 7604 17116
rect 7660 17660 7700 17669
rect 7660 16736 7700 17620
rect 7660 16687 7700 16696
rect 7756 13376 7796 55420
rect 7852 51176 7892 51185
rect 7852 45884 7892 51136
rect 7852 45835 7892 45844
rect 7756 13327 7796 13336
rect 7852 44792 7892 44801
rect 7564 8000 7604 8009
rect 7564 7748 7604 7960
rect 7564 7699 7604 7708
rect 7468 7111 7508 7120
rect 6892 2071 6932 2080
rect 7275 2120 7317 2129
rect 7275 2080 7276 2120
rect 7316 2080 7317 2120
rect 7275 2071 7317 2080
rect 7276 1986 7316 2071
rect 7852 1289 7892 44752
rect 7948 18761 7988 57931
rect 8140 57308 8180 83476
rect 8140 57259 8180 57268
rect 8236 83180 8276 83189
rect 8140 57140 8180 57149
rect 8140 53108 8180 57100
rect 8140 53059 8180 53068
rect 8044 51260 8084 51269
rect 8044 50840 8084 51220
rect 8044 50791 8084 50800
rect 8236 47900 8276 83140
rect 8523 76712 8565 76721
rect 8523 76672 8524 76712
rect 8564 76672 8565 76712
rect 8523 76663 8565 76672
rect 8524 76578 8564 76663
rect 8620 74528 8660 74537
rect 8332 69992 8372 70001
rect 8332 62516 8372 69952
rect 8332 62467 8372 62476
rect 8428 66884 8468 66893
rect 8332 56720 8372 56729
rect 8332 56216 8372 56680
rect 8332 56167 8372 56176
rect 8332 51260 8372 51269
rect 8332 50756 8372 51220
rect 8332 50707 8372 50716
rect 8236 47851 8276 47860
rect 8332 49664 8372 49673
rect 8140 46640 8180 46649
rect 8140 44792 8180 46600
rect 8140 44743 8180 44752
rect 8332 44120 8372 49624
rect 8332 44071 8372 44080
rect 8332 40256 8372 40265
rect 8235 35048 8277 35057
rect 8235 35008 8236 35048
rect 8276 35008 8277 35048
rect 8235 34999 8277 35008
rect 8236 34914 8276 34999
rect 8140 33788 8180 33797
rect 8044 25976 8084 25985
rect 7947 18752 7989 18761
rect 7947 18712 7948 18752
rect 7988 18712 7989 18752
rect 7947 18703 7989 18712
rect 8044 18584 8084 25936
rect 8044 18535 8084 18544
rect 7948 18500 7988 18509
rect 7948 17492 7988 18460
rect 7948 17443 7988 17452
rect 7948 14888 7988 14897
rect 7948 11444 7988 14848
rect 7948 11395 7988 11404
rect 8140 1868 8180 33748
rect 8236 29168 8276 29177
rect 8236 27152 8276 29128
rect 8236 27103 8276 27112
rect 8236 24632 8276 24641
rect 8236 17996 8276 24592
rect 8236 8000 8276 17956
rect 8236 7951 8276 7960
rect 8140 1819 8180 1828
rect 6796 1231 6836 1240
rect 7851 1280 7893 1289
rect 7851 1240 7852 1280
rect 7892 1240 7893 1280
rect 7851 1231 7893 1240
rect 3340 1063 3380 1072
rect 8332 860 8372 40216
rect 8428 18341 8468 66844
rect 8524 65540 8564 65549
rect 8524 64028 8564 65500
rect 8524 63979 8564 63988
rect 8524 60080 8564 60089
rect 8524 53864 8564 60040
rect 8524 53815 8564 53824
rect 8524 51176 8564 51185
rect 8524 48404 8564 51136
rect 8524 48355 8564 48364
rect 8524 47900 8564 47909
rect 8524 47312 8564 47860
rect 8427 18332 8469 18341
rect 8427 18292 8428 18332
rect 8468 18292 8469 18332
rect 8427 18283 8469 18292
rect 8428 12536 8468 12545
rect 8428 11108 8468 12496
rect 8428 11059 8468 11068
rect 8524 9764 8564 47272
rect 8620 14561 8660 74488
rect 8812 74444 8852 74453
rect 8716 73688 8756 73697
rect 8716 17408 8756 73648
rect 8812 17492 8852 74404
rect 8908 44876 8948 84316
rect 10252 78140 10292 78149
rect 9003 76712 9045 76721
rect 9003 76672 9004 76712
rect 9044 76672 9045 76712
rect 9003 76663 9045 76672
rect 9004 76578 9044 76663
rect 9388 74528 9428 74537
rect 9100 73688 9140 73697
rect 9004 69320 9044 69329
rect 9004 63944 9044 69280
rect 9004 63895 9044 63904
rect 9004 63188 9044 63197
rect 9004 61676 9044 63148
rect 9004 54788 9044 61636
rect 9004 54284 9044 54748
rect 9004 54235 9044 54244
rect 9004 52352 9044 52361
rect 9004 50420 9044 52312
rect 9004 50371 9044 50380
rect 8908 44827 8948 44836
rect 8800 17452 8852 17492
rect 8908 40424 8948 40433
rect 8800 17408 8840 17452
rect 8800 17368 8852 17408
rect 8716 17359 8756 17368
rect 8812 14888 8852 17368
rect 8812 14839 8852 14848
rect 8619 14552 8661 14561
rect 8619 14512 8620 14552
rect 8660 14512 8661 14552
rect 8619 14503 8661 14512
rect 8812 13544 8852 13553
rect 8812 9848 8852 13504
rect 8812 9799 8852 9808
rect 8524 9715 8564 9724
rect 8332 811 8372 820
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 748 559 788 568
rect 8908 281 8948 40384
rect 9004 39668 9044 39677
rect 9004 17585 9044 39628
rect 9100 35888 9140 73648
rect 9292 71504 9332 71513
rect 9196 60836 9236 60845
rect 9196 53612 9236 60796
rect 9196 53563 9236 53572
rect 9196 47480 9236 47489
rect 9196 46640 9236 47440
rect 9196 46591 9236 46600
rect 9100 35839 9140 35848
rect 9196 26396 9236 26405
rect 9100 23960 9140 23969
rect 9003 17576 9045 17585
rect 9003 17536 9004 17576
rect 9044 17536 9045 17576
rect 9003 17527 9045 17536
rect 9003 13208 9045 13217
rect 9003 13168 9004 13208
rect 9044 13168 9045 13208
rect 9003 13159 9045 13168
rect 9004 1028 9044 13159
rect 9004 979 9044 988
rect 5067 272 5109 281
rect 5067 232 5068 272
rect 5108 232 5109 272
rect 5067 223 5109 232
rect 8907 272 8949 281
rect 8907 232 8908 272
rect 8948 232 8949 272
rect 8907 223 8949 232
rect 3340 113 3380 198
rect 4875 188 4917 197
rect 4875 148 4876 188
rect 4916 148 4917 188
rect 4875 139 4917 148
rect 3339 104 3381 113
rect 3339 64 3340 104
rect 3380 64 3381 104
rect 3339 55 3381 64
rect 4876 54 4916 139
rect 5068 138 5108 223
rect 9100 113 9140 23920
rect 9196 8588 9236 26356
rect 9292 24632 9332 71464
rect 9292 24583 9332 24592
rect 9291 17576 9333 17585
rect 9291 17536 9292 17576
rect 9332 17536 9333 17576
rect 9291 17527 9333 17536
rect 9292 13217 9332 17527
rect 9388 16400 9428 74488
rect 9868 70748 9908 70757
rect 9772 61760 9812 61769
rect 9484 59744 9524 59753
rect 9484 57728 9524 59704
rect 9484 57679 9524 57688
rect 9484 54284 9524 54293
rect 9484 44624 9524 54244
rect 9772 53780 9812 61720
rect 9772 53731 9812 53740
rect 9772 50840 9812 50849
rect 9580 47564 9620 47573
rect 9580 46808 9620 47524
rect 9580 45800 9620 46768
rect 9580 45751 9620 45760
rect 9484 44575 9524 44584
rect 9772 36728 9812 50800
rect 9868 41264 9908 70708
rect 10060 59240 10100 59249
rect 10060 57989 10100 59200
rect 10059 57980 10101 57989
rect 10059 57940 10060 57980
rect 10100 57940 10101 57980
rect 10059 57931 10101 57940
rect 9964 57560 10004 57569
rect 9964 55460 10004 57520
rect 10060 57140 10100 57931
rect 10060 57091 10100 57100
rect 10156 55544 10196 55553
rect 9964 55420 10100 55460
rect 10060 54704 10100 55420
rect 10060 54655 10100 54664
rect 10156 54116 10196 55504
rect 10156 54067 10196 54076
rect 10156 52940 10196 52949
rect 10156 49328 10196 52900
rect 10156 49279 10196 49288
rect 10155 41936 10197 41945
rect 10155 41896 10156 41936
rect 10196 41896 10197 41936
rect 10155 41887 10197 41896
rect 10156 41802 10196 41887
rect 9868 41215 9908 41224
rect 10252 38240 10292 78100
rect 10444 77468 10484 77477
rect 10444 76292 10484 77428
rect 10444 76243 10484 76252
rect 10348 75872 10388 75881
rect 10348 42860 10388 75832
rect 10540 65372 10580 65381
rect 10540 64868 10580 65332
rect 10348 42811 10388 42820
rect 10444 61592 10484 61601
rect 10252 38191 10292 38200
rect 9676 36140 9716 36149
rect 9388 16351 9428 16360
rect 9484 35804 9524 35813
rect 9291 13208 9333 13217
rect 9291 13168 9292 13208
rect 9332 13168 9333 13208
rect 9291 13159 9333 13168
rect 9388 11276 9428 11285
rect 9388 8840 9428 11236
rect 9388 8791 9428 8800
rect 9196 8000 9236 8548
rect 9196 7951 9236 7960
rect 9484 608 9524 35764
rect 9676 30596 9716 36100
rect 9676 29840 9716 30556
rect 9580 22616 9620 22625
rect 9580 21692 9620 22576
rect 9580 21643 9620 21652
rect 9676 20768 9716 29800
rect 9676 20719 9716 20728
rect 9676 20096 9716 20105
rect 9676 18593 9716 20056
rect 9675 18584 9717 18593
rect 9675 18544 9676 18584
rect 9716 18544 9717 18584
rect 9675 18535 9717 18544
rect 9580 17828 9620 17837
rect 9580 17408 9620 17788
rect 9580 11024 9620 17368
rect 9580 10975 9620 10984
rect 9772 1280 9812 36688
rect 10060 36560 10100 36569
rect 9964 24464 10004 24473
rect 9868 24044 9908 24053
rect 9868 17240 9908 24004
rect 9964 20600 10004 24424
rect 9964 20551 10004 20560
rect 9868 17191 9908 17200
rect 9963 10268 10005 10277
rect 9963 10228 9964 10268
rect 10004 10228 10005 10268
rect 9963 10219 10005 10228
rect 9964 3716 10004 10219
rect 9964 3667 10004 3676
rect 9772 1231 9812 1240
rect 9484 559 9524 568
rect 10060 356 10100 36520
rect 10348 34796 10388 34805
rect 10348 33956 10388 34756
rect 10348 33907 10388 33916
rect 10156 24632 10196 24641
rect 10156 12620 10196 24592
rect 10444 21449 10484 61552
rect 10540 56384 10580 64828
rect 10540 56335 10580 56344
rect 10540 53612 10580 53621
rect 10540 53276 10580 53572
rect 10540 53227 10580 53236
rect 10540 52940 10580 52949
rect 10540 52100 10580 52900
rect 10540 52051 10580 52060
rect 10636 47144 10676 84400
rect 12172 84440 12212 84449
rect 10924 83600 10964 83609
rect 10924 68732 10964 83560
rect 11116 79316 11156 79325
rect 11116 78980 11156 79276
rect 10924 68683 10964 68692
rect 11020 76544 11060 76553
rect 10924 61424 10964 61433
rect 10731 57896 10773 57905
rect 10731 57856 10732 57896
rect 10772 57856 10773 57896
rect 10731 57847 10773 57856
rect 10732 51596 10772 57847
rect 10924 56468 10964 61384
rect 10924 56419 10964 56428
rect 10732 51547 10772 51556
rect 10828 54620 10868 54629
rect 10828 47480 10868 54580
rect 10924 54200 10964 54209
rect 10924 52352 10964 54160
rect 10924 52303 10964 52312
rect 10828 47431 10868 47440
rect 10636 47095 10676 47104
rect 10732 42776 10772 42787
rect 10732 42701 10772 42736
rect 10731 42692 10773 42701
rect 10731 42652 10732 42692
rect 10772 42652 10773 42692
rect 10731 42643 10773 42652
rect 10732 42104 10772 42643
rect 10732 42055 10772 42064
rect 11020 41936 11060 76504
rect 11020 41887 11060 41896
rect 10924 40340 10964 40349
rect 10540 39752 10580 39761
rect 10443 21440 10485 21449
rect 10443 21400 10444 21440
rect 10484 21400 10485 21440
rect 10443 21391 10485 21400
rect 10444 20180 10484 20189
rect 10348 19676 10388 19685
rect 10348 18416 10388 19636
rect 10444 19256 10484 20140
rect 10444 19207 10484 19216
rect 10348 18367 10388 18376
rect 10156 12571 10196 12580
rect 10540 1868 10580 39712
rect 10732 38408 10772 38417
rect 10540 1819 10580 1828
rect 10636 38156 10676 38165
rect 10636 1028 10676 38116
rect 10732 36560 10772 38368
rect 10732 36511 10772 36520
rect 10828 36392 10868 36401
rect 10828 35804 10868 36352
rect 10732 34376 10772 34385
rect 10732 28412 10772 34336
rect 10828 33704 10868 35764
rect 10828 33655 10868 33664
rect 10828 29336 10868 29345
rect 10828 28916 10868 29296
rect 10828 28867 10868 28876
rect 10732 26312 10772 28372
rect 10732 26272 10868 26312
rect 10732 24044 10772 24053
rect 10732 20768 10772 24004
rect 10732 20719 10772 20728
rect 10828 20180 10868 26272
rect 10732 20140 10868 20180
rect 10732 11285 10772 20140
rect 10828 20012 10868 20021
rect 10828 17492 10868 19972
rect 10828 17443 10868 17452
rect 10731 11276 10773 11285
rect 10731 11236 10732 11276
rect 10772 11236 10773 11276
rect 10731 11227 10773 11236
rect 10924 1868 10964 40300
rect 11116 38240 11156 78940
rect 11980 79064 12020 79073
rect 11884 74444 11924 74453
rect 11884 73604 11924 74404
rect 11884 73555 11924 73564
rect 11596 72932 11636 72941
rect 11596 72680 11636 72892
rect 11596 72631 11636 72640
rect 11211 72260 11253 72269
rect 11211 72220 11212 72260
rect 11252 72220 11253 72260
rect 11211 72211 11253 72220
rect 11212 62096 11252 72211
rect 11884 71336 11924 71345
rect 11404 68312 11444 68321
rect 11307 68060 11349 68069
rect 11307 68020 11308 68060
rect 11348 68020 11349 68060
rect 11307 68011 11349 68020
rect 11308 63860 11348 68011
rect 11404 65456 11444 68272
rect 11404 65407 11444 65416
rect 11788 66800 11828 66809
rect 11308 63811 11348 63820
rect 11212 62047 11252 62056
rect 11692 61088 11732 61097
rect 11116 38191 11156 38200
rect 11212 60836 11252 60845
rect 11116 34460 11156 34469
rect 11020 30260 11060 30269
rect 11020 23792 11060 30220
rect 11116 27320 11156 34420
rect 11116 27271 11156 27280
rect 11020 16232 11060 23752
rect 11116 23120 11156 23129
rect 11116 18752 11156 23080
rect 11212 19424 11252 60796
rect 11308 59240 11348 59249
rect 11308 59156 11348 59200
rect 11308 59116 11444 59156
rect 11404 58568 11444 59116
rect 11404 54452 11444 58528
rect 11499 56888 11541 56897
rect 11499 56848 11500 56888
rect 11540 56848 11541 56888
rect 11499 56839 11541 56848
rect 11404 52772 11444 54412
rect 11404 52723 11444 52732
rect 11500 49412 11540 56839
rect 11500 49363 11540 49372
rect 11596 56048 11636 56057
rect 11596 51428 11636 56008
rect 11692 54620 11732 61048
rect 11692 54571 11732 54580
rect 11788 58568 11828 66760
rect 11596 49244 11636 51388
rect 11404 49204 11636 49244
rect 11692 53108 11732 53117
rect 11404 45212 11444 49204
rect 11404 44969 11444 45172
rect 11500 48908 11540 48917
rect 11403 44960 11445 44969
rect 11403 44920 11404 44960
rect 11444 44920 11445 44960
rect 11403 44911 11445 44920
rect 11404 34964 11444 34973
rect 11404 27404 11444 34924
rect 11404 27355 11444 27364
rect 11308 23624 11348 23633
rect 11308 23372 11348 23584
rect 11308 23323 11348 23332
rect 11308 20768 11348 20777
rect 11308 20012 11348 20728
rect 11308 19963 11348 19972
rect 11212 19375 11252 19384
rect 11116 18703 11156 18712
rect 11307 17744 11349 17753
rect 11500 17744 11540 48868
rect 11307 17704 11308 17744
rect 11348 17704 11540 17744
rect 11596 42272 11636 42281
rect 11307 17695 11349 17704
rect 11404 16736 11444 17704
rect 11404 16687 11444 16696
rect 11020 16183 11060 16192
rect 11500 14636 11540 14645
rect 11500 13880 11540 14596
rect 11500 13831 11540 13840
rect 10924 1819 10964 1828
rect 11596 1196 11636 42232
rect 11692 1868 11732 53068
rect 11788 52436 11828 58528
rect 11788 52387 11828 52396
rect 11788 36308 11828 36317
rect 11788 34628 11828 36268
rect 11788 34579 11828 34588
rect 11788 17660 11828 17669
rect 11788 10772 11828 17620
rect 11788 10723 11828 10732
rect 11692 1819 11732 1828
rect 11596 1147 11636 1156
rect 10636 979 10676 988
rect 11884 440 11924 71296
rect 11980 61844 12020 79024
rect 11980 61795 12020 61804
rect 12076 75704 12116 75713
rect 11980 59828 12020 59837
rect 11980 42608 12020 59788
rect 11980 41600 12020 42568
rect 11980 41551 12020 41560
rect 11980 38492 12020 38501
rect 11980 37988 12020 38452
rect 11980 1868 12020 37948
rect 12076 14636 12116 75664
rect 12172 50756 12212 84400
rect 13324 84440 13364 84449
rect 12940 76628 12980 76637
rect 12940 76292 12980 76588
rect 12940 76243 12980 76252
rect 13227 75956 13269 75965
rect 13227 75916 13228 75956
rect 13268 75916 13269 75956
rect 13227 75907 13269 75916
rect 12268 73184 12308 73193
rect 12268 73016 12308 73144
rect 12268 72967 12308 72976
rect 13228 65624 13268 75907
rect 13228 65575 13268 65584
rect 12460 61508 12500 61517
rect 12172 50707 12212 50716
rect 12268 57476 12308 57485
rect 12076 14587 12116 14596
rect 12172 50084 12212 50093
rect 12172 12032 12212 50044
rect 12268 37316 12308 57436
rect 12460 56048 12500 61468
rect 12651 59912 12693 59921
rect 12651 59872 12652 59912
rect 12692 59872 12693 59912
rect 12651 59863 12693 59872
rect 12460 55999 12500 56008
rect 12268 37267 12308 37276
rect 12556 48572 12596 48581
rect 12364 34208 12404 34217
rect 12268 30848 12308 30857
rect 12268 27656 12308 30808
rect 12268 27607 12308 27616
rect 12268 23708 12308 23717
rect 12268 18836 12308 23668
rect 12268 18787 12308 18796
rect 12172 11983 12212 11992
rect 12076 11108 12116 11117
rect 12076 10445 12116 11068
rect 12075 10436 12117 10445
rect 12075 10396 12076 10436
rect 12116 10396 12117 10436
rect 12075 10387 12117 10396
rect 12364 5060 12404 34168
rect 12556 33713 12596 48532
rect 12652 42776 12692 59863
rect 13036 58820 13076 58829
rect 12652 36056 12692 42736
rect 12748 58568 12788 58577
rect 12748 38324 12788 58528
rect 12940 54200 12980 54209
rect 12940 53528 12980 54160
rect 12940 53479 12980 53488
rect 13036 53024 13076 58780
rect 13036 52975 13076 52984
rect 13132 57308 13172 57317
rect 13132 52016 13172 57268
rect 13132 51967 13172 51976
rect 13228 53780 13268 53789
rect 12844 51764 12884 51773
rect 12844 48488 12884 51724
rect 12844 48439 12884 48448
rect 13036 51512 13076 51521
rect 12748 38275 12788 38284
rect 12940 39668 12980 39677
rect 12652 36007 12692 36016
rect 12748 37820 12788 37829
rect 12748 37652 12788 37780
rect 12748 36644 12788 37612
rect 12555 33704 12597 33713
rect 12555 33664 12556 33704
rect 12596 33664 12597 33704
rect 12555 33655 12597 33664
rect 12364 5011 12404 5020
rect 11980 1819 12020 1828
rect 12748 1112 12788 36604
rect 12844 34376 12884 34385
rect 12844 30596 12884 34336
rect 12844 30547 12884 30556
rect 12844 11276 12884 11285
rect 12844 8420 12884 11236
rect 12844 8371 12884 8380
rect 12748 1063 12788 1072
rect 11884 391 11924 400
rect 10060 307 10100 316
rect 12940 188 12980 39628
rect 13036 36476 13076 51472
rect 13228 50588 13268 53740
rect 13228 50539 13268 50548
rect 13324 38240 13364 84400
rect 13708 84440 13748 84449
rect 13612 83516 13652 83525
rect 13420 76964 13460 76973
rect 13420 75536 13460 76924
rect 13420 75487 13460 75496
rect 13516 76712 13556 76721
rect 13516 74528 13556 76672
rect 13420 70748 13460 70757
rect 13420 59660 13460 70708
rect 13420 59611 13460 59620
rect 13420 56720 13460 56729
rect 13420 55544 13460 56680
rect 13420 46976 13460 55504
rect 13420 46927 13460 46936
rect 13324 38191 13364 38200
rect 13036 36427 13076 36436
rect 13228 36560 13268 36569
rect 13132 34628 13172 34637
rect 13132 31520 13172 34588
rect 13132 31471 13172 31480
rect 13036 25640 13076 25649
rect 13036 24884 13076 25600
rect 13036 22952 13076 24844
rect 13036 22903 13076 22912
rect 13132 23540 13172 23549
rect 13132 22112 13172 23500
rect 13132 22063 13172 22072
rect 13036 20264 13076 20273
rect 13036 16064 13076 20224
rect 13228 17156 13268 36520
rect 13228 17107 13268 17116
rect 13324 33368 13364 33377
rect 13324 16736 13364 33328
rect 13420 32696 13460 32705
rect 13420 32360 13460 32656
rect 13420 32311 13460 32320
rect 13324 16687 13364 16696
rect 13420 26480 13460 26489
rect 13420 25304 13460 26440
rect 13036 16015 13076 16024
rect 13131 15728 13173 15737
rect 13131 15688 13132 15728
rect 13172 15688 13173 15728
rect 13131 15679 13173 15688
rect 13036 11276 13076 11285
rect 13036 11117 13076 11236
rect 13035 11108 13077 11117
rect 13035 11068 13036 11108
rect 13076 11068 13077 11108
rect 13035 11059 13077 11068
rect 13132 2540 13172 15679
rect 13228 11780 13268 11789
rect 13228 11360 13268 11740
rect 13228 11311 13268 11320
rect 13420 7664 13460 25264
rect 13420 7615 13460 7624
rect 13036 2500 13172 2540
rect 13036 1196 13076 2500
rect 13036 1147 13076 1156
rect 13419 1196 13461 1205
rect 13419 1156 13420 1196
rect 13460 1156 13461 1196
rect 13419 1147 13461 1156
rect 13420 1062 13460 1147
rect 12940 139 12980 148
rect 9099 104 9141 113
rect 9099 64 9100 104
rect 9140 64 9141 104
rect 9099 55 9141 64
rect 13516 104 13556 74488
rect 13612 29756 13652 83476
rect 13708 45296 13748 84400
rect 13804 64616 13844 64625
rect 13804 62852 13844 64576
rect 13804 62803 13844 62812
rect 13708 45247 13748 45256
rect 13804 61004 13844 61013
rect 13804 40676 13844 60964
rect 13804 40340 13844 40636
rect 13804 40291 13844 40300
rect 13612 29707 13652 29716
rect 13804 30932 13844 30941
rect 13708 26480 13748 26489
rect 13708 18584 13748 26440
rect 13708 18535 13748 18544
rect 13708 18080 13748 18089
rect 13708 17240 13748 18040
rect 13708 17191 13748 17200
rect 13804 16652 13844 30892
rect 13804 16603 13844 16612
rect 13804 11444 13844 11453
rect 13804 11192 13844 11404
rect 13804 11143 13844 11152
rect 13803 2708 13845 2717
rect 13803 2668 13804 2708
rect 13844 2668 13845 2708
rect 13803 2659 13845 2668
rect 13804 2574 13844 2659
rect 13900 2120 13940 84568
rect 14284 84524 14324 84533
rect 13996 84440 14036 84449
rect 13996 41516 14036 84400
rect 14092 70580 14132 70589
rect 14092 68312 14132 70540
rect 14092 62852 14132 68272
rect 14092 62803 14132 62812
rect 14092 59744 14132 59753
rect 14092 46640 14132 59704
rect 14188 57140 14228 57149
rect 14188 56300 14228 57100
rect 14188 54956 14228 56260
rect 14188 54907 14228 54916
rect 14188 53948 14228 53957
rect 14188 52604 14228 53908
rect 14188 52555 14228 52564
rect 14284 48824 14324 84484
rect 14956 84524 14996 84533
rect 14668 84440 14708 84449
rect 14572 68228 14612 68237
rect 14476 62600 14516 62609
rect 14188 48784 14324 48824
rect 14380 60752 14420 60761
rect 14188 47648 14228 48784
rect 14283 47900 14325 47909
rect 14283 47860 14284 47900
rect 14324 47860 14325 47900
rect 14283 47851 14325 47860
rect 14284 47766 14324 47851
rect 14188 47608 14324 47648
rect 14092 46600 14228 46640
rect 13996 41467 14036 41476
rect 14092 41264 14132 41273
rect 14092 39584 14132 41224
rect 14092 38156 14132 39544
rect 14092 38107 14132 38116
rect 14092 32864 14132 32873
rect 13996 31352 14036 31361
rect 13996 28328 14036 31312
rect 13996 24548 14036 28288
rect 13996 24499 14036 24508
rect 14092 25304 14132 32824
rect 14092 23960 14132 25264
rect 14092 23911 14132 23920
rect 14092 22280 14132 22289
rect 14092 18668 14132 22240
rect 14188 21020 14228 46600
rect 14188 20971 14228 20980
rect 14092 18619 14132 18628
rect 13996 13712 14036 13721
rect 13996 9848 14036 13672
rect 13996 9799 14036 9808
rect 13900 2071 13940 2080
rect 14284 1868 14324 47608
rect 14380 29672 14420 60712
rect 14476 40760 14516 62560
rect 14572 53948 14612 68188
rect 14572 53899 14612 53908
rect 14476 40711 14516 40720
rect 14572 52436 14612 52445
rect 14380 29623 14420 29632
rect 14380 21524 14420 21533
rect 14380 2708 14420 21484
rect 14476 18920 14516 18929
rect 14476 18332 14516 18880
rect 14476 18283 14516 18292
rect 14572 13124 14612 52396
rect 14572 13075 14612 13084
rect 14380 2659 14420 2668
rect 14284 1819 14324 1828
rect 14668 1868 14708 84400
rect 14956 81920 14996 84484
rect 15051 84440 15093 84449
rect 15051 84400 15052 84440
rect 15092 84400 15093 84440
rect 15051 84391 15093 84400
rect 15532 84440 15572 84449
rect 15052 84306 15092 84391
rect 15340 83516 15380 83525
rect 14956 81880 15092 81920
rect 14860 71840 14900 71849
rect 14860 71084 14900 71800
rect 14860 71035 14900 71044
rect 14860 70580 14900 70589
rect 14860 64616 14900 70540
rect 14956 69908 14996 69917
rect 14956 67388 14996 69868
rect 15052 68648 15092 81880
rect 15148 76040 15188 76049
rect 15148 74024 15188 76000
rect 15148 73975 15188 73984
rect 15052 68599 15092 68608
rect 15148 69908 15188 69917
rect 14956 67339 14996 67348
rect 15148 66800 15188 69868
rect 14860 64567 14900 64576
rect 15052 66760 15188 66800
rect 15052 63860 15092 66760
rect 15052 63811 15092 63820
rect 15244 60164 15284 60173
rect 15244 59744 15284 60124
rect 14860 55628 14900 55637
rect 14860 55460 14900 55588
rect 14860 55411 14900 55420
rect 15244 54452 15284 59704
rect 15244 54403 15284 54412
rect 14860 51764 14900 51773
rect 14860 48404 14900 51724
rect 15340 49748 15380 83476
rect 15436 71840 15476 71849
rect 15436 71504 15476 71800
rect 15436 71455 15476 71464
rect 15340 49699 15380 49708
rect 15436 68648 15476 68657
rect 14860 48355 14900 48364
rect 15052 45296 15092 45305
rect 15052 44204 15092 45256
rect 15052 44155 15092 44164
rect 14860 41516 14900 41525
rect 14764 40760 14804 40769
rect 14764 38240 14804 40720
rect 14860 40424 14900 41476
rect 14860 40375 14900 40384
rect 14764 31352 14804 38200
rect 14764 31303 14804 31312
rect 14956 38912 14996 38921
rect 14860 29336 14900 29345
rect 14860 27068 14900 29296
rect 14860 27019 14900 27028
rect 14860 25472 14900 25481
rect 14764 22700 14804 22709
rect 14764 7169 14804 22660
rect 14860 13460 14900 25432
rect 14860 13411 14900 13420
rect 14763 7160 14805 7169
rect 14763 7120 14764 7160
rect 14804 7120 14805 7160
rect 14763 7111 14805 7120
rect 14668 1819 14708 1828
rect 14956 1196 14996 38872
rect 15148 37820 15188 37829
rect 15148 37652 15188 37780
rect 15148 37603 15188 37612
rect 15052 35048 15092 35057
rect 15052 33032 15092 35008
rect 15052 32983 15092 32992
rect 15340 34880 15380 34889
rect 15340 27824 15380 34840
rect 15340 27775 15380 27784
rect 15052 27152 15092 27161
rect 15052 26480 15092 27112
rect 15052 26440 15188 26480
rect 15148 18248 15188 26440
rect 15148 18199 15188 18208
rect 15340 24968 15380 24977
rect 15340 21692 15380 24928
rect 15340 17912 15380 21652
rect 15340 17863 15380 17872
rect 15147 14552 15189 14561
rect 15147 14512 15148 14552
rect 15188 14512 15189 14552
rect 15147 14503 15189 14512
rect 15148 14418 15188 14503
rect 15436 2120 15476 68608
rect 15436 2071 15476 2080
rect 15532 1868 15572 84400
rect 15820 69824 15860 69833
rect 15628 69236 15668 69245
rect 15628 61760 15668 69196
rect 15628 61711 15668 61720
rect 15436 1784 15476 1793
rect 15436 1280 15476 1744
rect 15436 1231 15476 1240
rect 14956 1147 14996 1156
rect 15532 1112 15572 1828
rect 15628 60920 15668 60929
rect 15628 1280 15668 60880
rect 15820 55040 15860 69784
rect 15916 59660 15956 59669
rect 15916 58988 15956 59620
rect 15916 58939 15956 58948
rect 15820 54991 15860 55000
rect 15916 55208 15956 55217
rect 15916 53696 15956 55168
rect 15916 53647 15956 53656
rect 15724 50672 15764 50681
rect 15724 47396 15764 50632
rect 15724 47347 15764 47356
rect 15724 42860 15764 42869
rect 15724 17669 15764 42820
rect 15820 37904 15860 37913
rect 15820 36476 15860 37864
rect 15820 36427 15860 36436
rect 15820 22532 15860 22541
rect 15820 21188 15860 22492
rect 15820 21139 15860 21148
rect 15916 18920 15956 18929
rect 15723 17660 15765 17669
rect 15723 17620 15724 17660
rect 15764 17620 15765 17660
rect 15723 17611 15765 17620
rect 15723 16820 15765 16829
rect 15723 16780 15724 16820
rect 15764 16780 15765 16820
rect 15723 16771 15765 16780
rect 15724 16686 15764 16771
rect 15916 16232 15956 18880
rect 15916 16183 15956 16192
rect 15724 14384 15764 14393
rect 15724 13880 15764 14344
rect 15724 13831 15764 13840
rect 16012 1868 16052 85576
rect 16876 85616 16916 85625
rect 16396 84944 16436 84953
rect 16204 83516 16244 83525
rect 16108 70580 16148 70589
rect 16108 63104 16148 70540
rect 16108 63055 16148 63064
rect 16108 61928 16148 61937
rect 16108 57980 16148 61888
rect 16108 57931 16148 57940
rect 16108 52856 16148 52865
rect 16108 51680 16148 52816
rect 16108 51631 16148 51640
rect 16108 51092 16148 51101
rect 16108 45800 16148 51052
rect 16108 45751 16148 45760
rect 16012 1819 16052 1828
rect 16108 35300 16148 35309
rect 15628 1231 15668 1240
rect 16108 1196 16148 35260
rect 16204 12368 16244 83476
rect 16300 74024 16340 74033
rect 16300 71504 16340 73984
rect 16300 61508 16340 71464
rect 16300 61459 16340 61468
rect 16300 57056 16340 57065
rect 16300 53192 16340 57016
rect 16300 53143 16340 53152
rect 16300 52100 16340 52109
rect 16300 51596 16340 52060
rect 16300 51547 16340 51556
rect 16396 38912 16436 84904
rect 16780 84524 16820 84533
rect 16588 77468 16628 77477
rect 16492 72176 16532 72185
rect 16492 71252 16532 72136
rect 16492 71203 16532 71212
rect 16492 69824 16532 69833
rect 16492 48656 16532 69784
rect 16588 67892 16628 77428
rect 16588 67843 16628 67852
rect 16684 61424 16724 61433
rect 16684 58568 16724 61384
rect 16684 55796 16724 58528
rect 16684 55747 16724 55756
rect 16492 48488 16532 48616
rect 16492 48439 16532 48448
rect 16684 54620 16724 54629
rect 16396 38863 16436 38872
rect 16492 39668 16532 39677
rect 16300 28328 16340 28337
rect 16300 26060 16340 28288
rect 16300 26011 16340 26020
rect 16492 23204 16532 39628
rect 16684 35300 16724 54580
rect 16684 35251 16724 35260
rect 16492 23155 16532 23164
rect 16588 33620 16628 33629
rect 16588 33032 16628 33580
rect 16396 22364 16436 22373
rect 16300 20432 16340 20441
rect 16300 19844 16340 20392
rect 16300 18920 16340 19804
rect 16300 18871 16340 18880
rect 16396 19928 16436 22324
rect 16588 20096 16628 32992
rect 16396 18164 16436 19888
rect 16396 17660 16436 18124
rect 16492 20056 16588 20096
rect 16492 17912 16532 20056
rect 16588 20047 16628 20056
rect 16684 25976 16724 25985
rect 16492 17863 16532 17872
rect 16588 19676 16628 19685
rect 16300 17620 16436 17660
rect 16300 16568 16340 17620
rect 16300 16519 16340 16528
rect 16204 12319 16244 12328
rect 16300 15728 16340 15737
rect 16204 11696 16244 11705
rect 16204 9512 16244 11656
rect 16204 9463 16244 9472
rect 16300 2120 16340 15688
rect 16395 15560 16437 15569
rect 16395 15520 16396 15560
rect 16436 15520 16437 15560
rect 16395 15511 16437 15520
rect 16396 15392 16436 15511
rect 16396 15343 16436 15352
rect 16492 15308 16532 15317
rect 16396 11444 16436 11453
rect 16396 11276 16436 11404
rect 16396 11227 16436 11236
rect 16396 6740 16436 6749
rect 16396 6572 16436 6700
rect 16396 6523 16436 6532
rect 16492 2540 16532 15268
rect 16300 2071 16340 2080
rect 16396 2500 16532 2540
rect 16396 1868 16436 2500
rect 16396 1819 16436 1828
rect 16588 1868 16628 19636
rect 16684 17072 16724 25936
rect 16684 12116 16724 17032
rect 16780 15728 16820 84484
rect 16876 59576 16916 85576
rect 17931 85112 17973 85121
rect 17931 85072 17932 85112
rect 17972 85072 17973 85112
rect 17931 85063 17973 85072
rect 19852 85112 19892 85121
rect 17932 84978 17972 85063
rect 18808 84692 19176 84701
rect 18848 84652 18890 84692
rect 18930 84652 18972 84692
rect 19012 84652 19054 84692
rect 19094 84652 19136 84692
rect 18808 84643 19176 84652
rect 17740 84524 17780 84533
rect 17260 84440 17300 84449
rect 16972 78140 17012 78149
rect 16972 70076 17012 78100
rect 17068 77636 17108 77645
rect 17068 77216 17108 77596
rect 17068 75200 17108 77176
rect 17068 71000 17108 75160
rect 17164 72848 17204 72857
rect 17164 72008 17204 72808
rect 17164 71959 17204 71968
rect 17068 70951 17108 70960
rect 16972 70027 17012 70036
rect 16972 67388 17012 67397
rect 16972 65960 17012 67348
rect 16972 65911 17012 65920
rect 16876 59527 16916 59536
rect 17164 61844 17204 61853
rect 16876 53948 16916 53957
rect 16876 52184 16916 53908
rect 16971 53276 17013 53285
rect 16971 53236 16972 53276
rect 17012 53236 17013 53276
rect 16971 53227 17013 53236
rect 16876 52135 16916 52144
rect 16876 33284 16916 33293
rect 16876 27236 16916 33244
rect 16972 32276 17012 53227
rect 17068 50840 17108 50849
rect 17068 33545 17108 50800
rect 17067 33536 17109 33545
rect 17067 33496 17068 33536
rect 17108 33496 17109 33536
rect 17067 33487 17109 33496
rect 16972 32227 17012 32236
rect 17068 31016 17108 31025
rect 17068 29840 17108 30976
rect 17068 29791 17108 29800
rect 16876 27187 16916 27196
rect 16972 29672 17012 29681
rect 16972 26900 17012 29632
rect 17067 28496 17109 28505
rect 17067 28456 17068 28496
rect 17108 28456 17109 28496
rect 17067 28447 17109 28456
rect 16972 26851 17012 26860
rect 17068 25976 17108 28447
rect 17068 25927 17108 25936
rect 16876 25640 16916 25649
rect 16876 22364 16916 25600
rect 16876 22315 16916 22324
rect 17068 23792 17108 23801
rect 16780 15679 16820 15688
rect 16876 22196 16916 22205
rect 16684 12067 16724 12076
rect 16876 11444 16916 22156
rect 16972 21944 17012 21953
rect 16972 20096 17012 21904
rect 17068 20264 17108 23752
rect 17068 20215 17108 20224
rect 16972 20056 17108 20096
rect 17068 18416 17108 20056
rect 17068 14384 17108 18376
rect 17068 14335 17108 14344
rect 16876 11395 16916 11404
rect 17164 7076 17204 61804
rect 17260 56552 17300 84400
rect 17548 84440 17588 84449
rect 17452 69320 17492 69329
rect 17452 57140 17492 69280
rect 17452 57091 17492 57100
rect 17260 56503 17300 56512
rect 17452 56636 17492 56645
rect 17356 56300 17396 56309
rect 17260 53780 17300 53789
rect 17260 51596 17300 53740
rect 17356 53696 17396 56260
rect 17452 54116 17492 56596
rect 17452 54067 17492 54076
rect 17356 53647 17396 53656
rect 17260 51547 17300 51556
rect 17452 53276 17492 53285
rect 17452 45716 17492 53236
rect 17452 45667 17492 45676
rect 17356 36056 17396 36065
rect 17260 33536 17300 33545
rect 17260 29756 17300 33496
rect 17260 28505 17300 29716
rect 17259 28496 17301 28505
rect 17259 28456 17260 28496
rect 17300 28456 17301 28496
rect 17259 28447 17301 28456
rect 17260 28328 17300 28337
rect 17356 28328 17396 36016
rect 17452 34544 17492 34553
rect 17452 33032 17492 34504
rect 17452 32983 17492 32992
rect 17452 32780 17492 32789
rect 17452 29924 17492 32740
rect 17452 29875 17492 29884
rect 17300 28288 17396 28328
rect 17260 20348 17300 28288
rect 17452 27068 17492 27077
rect 17452 25640 17492 27028
rect 17452 25591 17492 25600
rect 17260 20299 17300 20308
rect 17356 23204 17396 23213
rect 17260 20180 17300 20189
rect 17260 17828 17300 20140
rect 17260 13544 17300 17788
rect 17260 13495 17300 13504
rect 17260 11696 17300 11705
rect 17260 10856 17300 11656
rect 17356 11360 17396 23164
rect 17452 23036 17492 23045
rect 17452 17996 17492 22996
rect 17452 17947 17492 17956
rect 17356 11320 17492 11360
rect 17260 10807 17300 10816
rect 17164 7027 17204 7036
rect 17452 9512 17492 11320
rect 17452 6740 17492 9472
rect 17452 6691 17492 6700
rect 17548 2120 17588 84400
rect 17644 70832 17684 70841
rect 17644 68984 17684 70792
rect 17644 68935 17684 68944
rect 17644 68648 17684 68657
rect 17644 68144 17684 68608
rect 17644 68095 17684 68104
rect 17644 56720 17684 56729
rect 17644 54032 17684 56680
rect 17644 53983 17684 53992
rect 17643 51848 17685 51857
rect 17643 51808 17644 51848
rect 17684 51808 17685 51848
rect 17643 51799 17685 51808
rect 17644 51714 17684 51799
rect 17644 32696 17684 32705
rect 17644 29588 17684 32656
rect 17644 29539 17684 29548
rect 17643 29420 17685 29429
rect 17643 29380 17644 29420
rect 17684 29380 17685 29420
rect 17643 29371 17685 29380
rect 17644 21608 17684 29371
rect 17644 21559 17684 21568
rect 17740 2288 17780 84484
rect 18604 84524 18644 84533
rect 17740 2239 17780 2248
rect 17836 84440 17876 84449
rect 17548 2071 17588 2080
rect 16588 1819 16628 1828
rect 17836 1280 17876 84400
rect 18412 84440 18452 84449
rect 18124 73268 18164 73277
rect 17932 73100 17972 73109
rect 17932 71168 17972 73060
rect 18124 72848 18164 73228
rect 18124 72799 18164 72808
rect 17932 69740 17972 71128
rect 17932 69691 17972 69700
rect 18028 69236 18068 69245
rect 17932 66128 17972 66137
rect 17932 65456 17972 66088
rect 18028 65960 18068 69196
rect 18028 65911 18068 65920
rect 18124 68060 18164 68069
rect 18124 67556 18164 68020
rect 17932 63776 17972 65416
rect 17932 63727 17972 63736
rect 18124 63104 18164 67516
rect 18124 63055 18164 63064
rect 18316 61592 18356 61601
rect 18028 58568 18068 58577
rect 18028 53360 18068 58528
rect 18220 58064 18260 58073
rect 18220 54788 18260 58024
rect 18220 54739 18260 54748
rect 18028 53311 18068 53320
rect 18028 53024 18068 53033
rect 17932 52184 17972 52193
rect 17932 48992 17972 52144
rect 18028 51680 18068 52984
rect 18028 51631 18068 51640
rect 17932 48943 17972 48952
rect 18316 49496 18356 61552
rect 18316 47564 18356 49456
rect 18316 47515 18356 47524
rect 18124 46892 18164 46901
rect 18028 46724 18068 46733
rect 18028 45725 18068 46684
rect 18124 46304 18164 46852
rect 18124 46255 18164 46264
rect 18027 45716 18069 45725
rect 18027 45676 18028 45716
rect 18068 45676 18069 45716
rect 18027 45667 18069 45676
rect 18316 38156 18356 38165
rect 18316 35720 18356 38116
rect 18316 35300 18356 35680
rect 18316 35251 18356 35260
rect 18028 35132 18068 35141
rect 17932 33032 17972 33041
rect 17932 29429 17972 32992
rect 18028 30680 18068 35092
rect 18124 33788 18164 33797
rect 18124 31436 18164 33748
rect 18124 31387 18164 31396
rect 18220 32696 18260 32705
rect 18220 32192 18260 32656
rect 18028 30631 18068 30640
rect 17931 29420 17973 29429
rect 17931 29380 17932 29420
rect 17972 29380 17973 29420
rect 17931 29371 17973 29380
rect 18124 25052 18164 25061
rect 18028 15980 18068 15989
rect 18028 13880 18068 15940
rect 18028 13831 18068 13840
rect 18028 10520 18068 10529
rect 17932 10352 17972 10361
rect 17932 9848 17972 10312
rect 17932 9799 17972 9808
rect 18028 9764 18068 10480
rect 18028 9715 18068 9724
rect 18124 2120 18164 25012
rect 18220 15392 18260 32152
rect 18316 29588 18356 29597
rect 18316 27656 18356 29548
rect 18316 27607 18356 27616
rect 18315 24632 18357 24641
rect 18315 24592 18316 24632
rect 18356 24592 18357 24632
rect 18315 24583 18357 24592
rect 18220 15343 18260 15352
rect 18219 10436 18261 10445
rect 18219 10396 18220 10436
rect 18260 10396 18261 10436
rect 18219 10387 18261 10396
rect 18220 10302 18260 10387
rect 18124 2071 18164 2080
rect 18316 2120 18356 24583
rect 18316 2071 18356 2080
rect 17836 1231 17876 1240
rect 18412 1280 18452 84400
rect 18508 63776 18548 63785
rect 18508 60752 18548 63736
rect 18508 21188 18548 60712
rect 18604 25220 18644 84484
rect 19660 84440 19700 84449
rect 18808 83180 19176 83189
rect 18848 83140 18890 83180
rect 18930 83140 18972 83180
rect 19012 83140 19054 83180
rect 19094 83140 19136 83180
rect 18808 83131 19176 83140
rect 19276 82760 19316 82769
rect 18808 81668 19176 81677
rect 18848 81628 18890 81668
rect 18930 81628 18972 81668
rect 19012 81628 19054 81668
rect 19094 81628 19136 81668
rect 18808 81619 19176 81628
rect 18808 80156 19176 80165
rect 18848 80116 18890 80156
rect 18930 80116 18972 80156
rect 19012 80116 19054 80156
rect 19094 80116 19136 80156
rect 18808 80107 19176 80116
rect 18808 78644 19176 78653
rect 18848 78604 18890 78644
rect 18930 78604 18972 78644
rect 19012 78604 19054 78644
rect 19094 78604 19136 78644
rect 18808 78595 19176 78604
rect 18808 77132 19176 77141
rect 18848 77092 18890 77132
rect 18930 77092 18972 77132
rect 19012 77092 19054 77132
rect 19094 77092 19136 77132
rect 18808 77083 19176 77092
rect 18891 75956 18933 75965
rect 18891 75916 18892 75956
rect 18932 75916 18933 75956
rect 18891 75907 18933 75916
rect 18892 75822 18932 75907
rect 18808 75620 19176 75629
rect 18848 75580 18890 75620
rect 18930 75580 18972 75620
rect 19012 75580 19054 75620
rect 19094 75580 19136 75620
rect 18808 75571 19176 75580
rect 18808 74108 19176 74117
rect 18848 74068 18890 74108
rect 18930 74068 18972 74108
rect 19012 74068 19054 74108
rect 19094 74068 19136 74108
rect 18808 74059 19176 74068
rect 18700 73688 18740 73697
rect 18700 72428 18740 73648
rect 18808 72596 19176 72605
rect 18848 72556 18890 72596
rect 18930 72556 18972 72596
rect 19012 72556 19054 72596
rect 19094 72556 19136 72596
rect 18808 72547 19176 72556
rect 18700 72379 18740 72388
rect 18808 71084 19176 71093
rect 18848 71044 18890 71084
rect 18930 71044 18972 71084
rect 19012 71044 19054 71084
rect 19094 71044 19136 71084
rect 18808 71035 19176 71044
rect 18808 69572 19176 69581
rect 18848 69532 18890 69572
rect 18930 69532 18972 69572
rect 19012 69532 19054 69572
rect 19094 69532 19136 69572
rect 18808 69523 19176 69532
rect 18808 68060 19176 68069
rect 18848 68020 18890 68060
rect 18930 68020 18972 68060
rect 19012 68020 19054 68060
rect 19094 68020 19136 68060
rect 18808 68011 19176 68020
rect 18808 66548 19176 66557
rect 18848 66508 18890 66548
rect 18930 66508 18972 66548
rect 19012 66508 19054 66548
rect 19094 66508 19136 66548
rect 18808 66499 19176 66508
rect 18808 65036 19176 65045
rect 18848 64996 18890 65036
rect 18930 64996 18972 65036
rect 19012 64996 19054 65036
rect 19094 64996 19136 65036
rect 18808 64987 19176 64996
rect 18808 63524 19176 63533
rect 18848 63484 18890 63524
rect 18930 63484 18972 63524
rect 19012 63484 19054 63524
rect 19094 63484 19136 63524
rect 18808 63475 19176 63484
rect 18808 62012 19176 62021
rect 18848 61972 18890 62012
rect 18930 61972 18972 62012
rect 19012 61972 19054 62012
rect 19094 61972 19136 62012
rect 18808 61963 19176 61972
rect 18808 60500 19176 60509
rect 18848 60460 18890 60500
rect 18930 60460 18972 60500
rect 19012 60460 19054 60500
rect 19094 60460 19136 60500
rect 18808 60451 19176 60460
rect 18700 59324 18740 59333
rect 18700 55460 18740 59284
rect 18808 58988 19176 58997
rect 18848 58948 18890 58988
rect 18930 58948 18972 58988
rect 19012 58948 19054 58988
rect 19094 58948 19136 58988
rect 18808 58939 19176 58948
rect 18808 57476 19176 57485
rect 18848 57436 18890 57476
rect 18930 57436 18972 57476
rect 19012 57436 19054 57476
rect 19094 57436 19136 57476
rect 18808 57427 19176 57436
rect 18808 55964 19176 55973
rect 18848 55924 18890 55964
rect 18930 55924 18972 55964
rect 19012 55924 19054 55964
rect 19094 55924 19136 55964
rect 18808 55915 19176 55924
rect 18700 55411 18740 55420
rect 18808 54452 19176 54461
rect 18848 54412 18890 54452
rect 18930 54412 18972 54452
rect 19012 54412 19054 54452
rect 19094 54412 19136 54452
rect 18808 54403 19176 54412
rect 18699 53276 18741 53285
rect 18699 53236 18700 53276
rect 18740 53236 18741 53276
rect 18699 53227 18741 53236
rect 18700 53024 18740 53227
rect 18700 52975 18740 52984
rect 18808 52940 19176 52949
rect 18848 52900 18890 52940
rect 18930 52900 18972 52940
rect 19012 52900 19054 52940
rect 19094 52900 19136 52940
rect 18808 52891 19176 52900
rect 19276 51680 19316 82720
rect 19564 78392 19604 78401
rect 19468 76544 19508 76553
rect 19468 75536 19508 76504
rect 19564 76460 19604 78352
rect 19564 76411 19604 76420
rect 19468 75487 19508 75496
rect 19660 64280 19700 84400
rect 19756 77468 19796 77477
rect 19756 75704 19796 77428
rect 19756 75655 19796 75664
rect 19852 73940 19892 85072
rect 20620 84944 20660 84953
rect 20048 83936 20416 83945
rect 20088 83896 20130 83936
rect 20170 83896 20212 83936
rect 20252 83896 20294 83936
rect 20334 83896 20376 83936
rect 20048 83887 20416 83896
rect 20048 82424 20416 82433
rect 20088 82384 20130 82424
rect 20170 82384 20212 82424
rect 20252 82384 20294 82424
rect 20334 82384 20376 82424
rect 20048 82375 20416 82384
rect 20048 80912 20416 80921
rect 20088 80872 20130 80912
rect 20170 80872 20212 80912
rect 20252 80872 20294 80912
rect 20334 80872 20376 80912
rect 20048 80863 20416 80872
rect 20048 79400 20416 79409
rect 20088 79360 20130 79400
rect 20170 79360 20212 79400
rect 20252 79360 20294 79400
rect 20334 79360 20376 79400
rect 20048 79351 20416 79360
rect 20524 78812 20564 78821
rect 20048 77888 20416 77897
rect 20088 77848 20130 77888
rect 20170 77848 20212 77888
rect 20252 77848 20294 77888
rect 20334 77848 20376 77888
rect 20048 77839 20416 77848
rect 20524 77720 20564 78772
rect 20524 77671 20564 77680
rect 20620 77552 20660 84904
rect 20524 77512 20660 77552
rect 20716 84608 20756 84617
rect 19948 76796 19988 76805
rect 19948 74024 19988 76756
rect 20048 76376 20416 76385
rect 20088 76336 20130 76376
rect 20170 76336 20212 76376
rect 20252 76336 20294 76376
rect 20334 76336 20376 76376
rect 20048 76327 20416 76336
rect 20048 74864 20416 74873
rect 20088 74824 20130 74864
rect 20170 74824 20212 74864
rect 20252 74824 20294 74864
rect 20334 74824 20376 74864
rect 20048 74815 20416 74824
rect 19948 73975 19988 73984
rect 19852 73891 19892 73900
rect 20048 73352 20416 73361
rect 20088 73312 20130 73352
rect 20170 73312 20212 73352
rect 20252 73312 20294 73352
rect 20334 73312 20376 73352
rect 20048 73303 20416 73312
rect 20140 73100 20180 73109
rect 20140 72932 20180 73060
rect 20140 72883 20180 72892
rect 19755 72260 19797 72269
rect 19755 72220 19756 72260
rect 19796 72220 19797 72260
rect 19755 72211 19797 72220
rect 19948 72260 19988 72269
rect 19756 72126 19796 72211
rect 19948 71672 19988 72220
rect 20048 71840 20416 71849
rect 20088 71800 20130 71840
rect 20170 71800 20212 71840
rect 20252 71800 20294 71840
rect 20334 71800 20376 71840
rect 20048 71791 20416 71800
rect 19948 71623 19988 71632
rect 20048 70328 20416 70337
rect 20088 70288 20130 70328
rect 20170 70288 20212 70328
rect 20252 70288 20294 70328
rect 20334 70288 20376 70328
rect 20048 70279 20416 70288
rect 20048 68816 20416 68825
rect 20088 68776 20130 68816
rect 20170 68776 20212 68816
rect 20252 68776 20294 68816
rect 20334 68776 20376 68816
rect 20048 68767 20416 68776
rect 20048 67304 20416 67313
rect 20088 67264 20130 67304
rect 20170 67264 20212 67304
rect 20252 67264 20294 67304
rect 20334 67264 20376 67304
rect 20048 67255 20416 67264
rect 20048 65792 20416 65801
rect 20088 65752 20130 65792
rect 20170 65752 20212 65792
rect 20252 65752 20294 65792
rect 20334 65752 20376 65792
rect 20048 65743 20416 65752
rect 20048 64280 20416 64289
rect 19660 64240 19796 64280
rect 19372 60668 19412 60677
rect 19372 56888 19412 60628
rect 19372 56839 19412 56848
rect 19564 56888 19604 56897
rect 19372 56552 19412 56561
rect 19372 53612 19412 56512
rect 19372 53563 19412 53572
rect 19468 55460 19508 55469
rect 19276 51631 19316 51640
rect 19372 52436 19412 52445
rect 18808 51428 19176 51437
rect 18848 51388 18890 51428
rect 18930 51388 18972 51428
rect 19012 51388 19054 51428
rect 19094 51388 19136 51428
rect 18808 51379 19176 51388
rect 19276 51008 19316 51017
rect 18808 49916 19176 49925
rect 18848 49876 18890 49916
rect 18930 49876 18972 49916
rect 19012 49876 19054 49916
rect 19094 49876 19136 49916
rect 18808 49867 19176 49876
rect 18808 48404 19176 48413
rect 18848 48364 18890 48404
rect 18930 48364 18972 48404
rect 19012 48364 19054 48404
rect 19094 48364 19136 48404
rect 18808 48355 19176 48364
rect 18808 46892 19176 46901
rect 18848 46852 18890 46892
rect 18930 46852 18972 46892
rect 19012 46852 19054 46892
rect 19094 46852 19136 46892
rect 18808 46843 19176 46852
rect 18700 46472 18740 46481
rect 18700 44456 18740 46432
rect 18808 45380 19176 45389
rect 18848 45340 18890 45380
rect 18930 45340 18972 45380
rect 19012 45340 19054 45380
rect 19094 45340 19136 45380
rect 18808 45331 19176 45340
rect 19276 44708 19316 50968
rect 19372 48908 19412 52396
rect 19372 48859 19412 48868
rect 19468 48068 19508 55420
rect 19564 49832 19604 56848
rect 19660 55124 19700 55133
rect 19660 52016 19700 55084
rect 19660 50084 19700 51976
rect 19660 50035 19700 50044
rect 19564 49783 19604 49792
rect 19468 48019 19508 48028
rect 19276 44659 19316 44668
rect 18700 44407 18740 44416
rect 18808 43868 19176 43877
rect 18848 43828 18890 43868
rect 18930 43828 18972 43868
rect 19012 43828 19054 43868
rect 19094 43828 19136 43868
rect 18808 43819 19176 43828
rect 18808 42356 19176 42365
rect 18848 42316 18890 42356
rect 18930 42316 18972 42356
rect 19012 42316 19054 42356
rect 19094 42316 19136 42356
rect 18808 42307 19176 42316
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 19564 37988 19604 37997
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 19468 36308 19508 36317
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 18700 33704 18740 33713
rect 18700 32276 18740 33664
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 18700 32227 18740 32236
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 19372 29672 19412 29681
rect 19276 29252 19316 29261
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 18604 25171 18644 25180
rect 18700 25724 18740 25733
rect 18700 25220 18740 25684
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 19276 25640 19316 29212
rect 19276 25591 19316 25600
rect 18796 25220 18836 25229
rect 18700 25180 18796 25220
rect 18700 23960 18740 25180
rect 18796 25171 18836 25180
rect 19276 24632 19316 24641
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 18700 23911 18740 23920
rect 18508 21139 18548 21148
rect 18604 22700 18644 22709
rect 18508 16820 18548 16829
rect 18508 15224 18548 16780
rect 18508 15175 18548 15184
rect 18508 14720 18548 14729
rect 18508 10520 18548 14680
rect 18508 10471 18548 10480
rect 18604 2120 18644 22660
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 19276 21020 19316 24592
rect 19372 23624 19412 29632
rect 19468 29252 19508 36268
rect 19468 29203 19508 29212
rect 19564 28664 19604 37948
rect 19660 36392 19700 36401
rect 19660 35048 19700 36352
rect 19660 34999 19700 35008
rect 19564 28615 19604 28624
rect 19756 28244 19796 64240
rect 20088 64240 20130 64280
rect 20170 64240 20212 64280
rect 20252 64240 20294 64280
rect 20334 64240 20376 64280
rect 20048 64231 20416 64240
rect 20048 62768 20416 62777
rect 20088 62728 20130 62768
rect 20170 62728 20212 62768
rect 20252 62728 20294 62768
rect 20334 62728 20376 62768
rect 20048 62719 20416 62728
rect 20048 61256 20416 61265
rect 20088 61216 20130 61256
rect 20170 61216 20212 61256
rect 20252 61216 20294 61256
rect 20334 61216 20376 61256
rect 20048 61207 20416 61216
rect 20048 59744 20416 59753
rect 20088 59704 20130 59744
rect 20170 59704 20212 59744
rect 20252 59704 20294 59744
rect 20334 59704 20376 59744
rect 20048 59695 20416 59704
rect 20048 58232 20416 58241
rect 20088 58192 20130 58232
rect 20170 58192 20212 58232
rect 20252 58192 20294 58232
rect 20334 58192 20376 58232
rect 20048 58183 20416 58192
rect 20048 56720 20416 56729
rect 20088 56680 20130 56720
rect 20170 56680 20212 56720
rect 20252 56680 20294 56720
rect 20334 56680 20376 56720
rect 20048 56671 20416 56680
rect 20048 55208 20416 55217
rect 20088 55168 20130 55208
rect 20170 55168 20212 55208
rect 20252 55168 20294 55208
rect 20334 55168 20376 55208
rect 20048 55159 20416 55168
rect 19948 54032 19988 54041
rect 19852 53612 19892 53621
rect 19852 50924 19892 53572
rect 19948 53192 19988 53992
rect 20048 53696 20416 53705
rect 20088 53656 20130 53696
rect 20170 53656 20212 53696
rect 20252 53656 20294 53696
rect 20334 53656 20376 53696
rect 20048 53647 20416 53656
rect 19948 53143 19988 53152
rect 20139 53192 20181 53201
rect 20139 53152 20140 53192
rect 20180 53152 20181 53192
rect 20139 53143 20181 53152
rect 20140 53058 20180 53143
rect 19948 52856 19988 52865
rect 19948 52184 19988 52816
rect 19948 52135 19988 52144
rect 20048 52184 20416 52193
rect 20088 52144 20130 52184
rect 20170 52144 20212 52184
rect 20252 52144 20294 52184
rect 20334 52144 20376 52184
rect 20048 52135 20416 52144
rect 19852 50875 19892 50884
rect 19948 50840 19988 50849
rect 19852 50672 19892 50681
rect 19852 45464 19892 50632
rect 19948 50420 19988 50800
rect 20048 50672 20416 50681
rect 20088 50632 20130 50672
rect 20170 50632 20212 50672
rect 20252 50632 20294 50672
rect 20334 50632 20376 50672
rect 20048 50623 20416 50632
rect 19948 50371 19988 50380
rect 19948 49328 19988 49337
rect 19948 46472 19988 49288
rect 20048 49160 20416 49169
rect 20088 49120 20130 49160
rect 20170 49120 20212 49160
rect 20252 49120 20294 49160
rect 20334 49120 20376 49160
rect 20048 49111 20416 49120
rect 20048 47648 20416 47657
rect 20088 47608 20130 47648
rect 20170 47608 20212 47648
rect 20252 47608 20294 47648
rect 20334 47608 20376 47648
rect 20048 47599 20416 47608
rect 19948 46423 19988 46432
rect 20048 46136 20416 46145
rect 20088 46096 20130 46136
rect 20170 46096 20212 46136
rect 20252 46096 20294 46136
rect 20334 46096 20376 46136
rect 20048 46087 20416 46096
rect 19852 45212 19892 45424
rect 19852 45163 19892 45172
rect 20048 44624 20416 44633
rect 20088 44584 20130 44624
rect 20170 44584 20212 44624
rect 20252 44584 20294 44624
rect 20334 44584 20376 44624
rect 20048 44575 20416 44584
rect 20048 43112 20416 43121
rect 20088 43072 20130 43112
rect 20170 43072 20212 43112
rect 20252 43072 20294 43112
rect 20334 43072 20376 43112
rect 20048 43063 20416 43072
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 19852 38156 19892 38165
rect 19852 36140 19892 38116
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 19852 36091 19892 36100
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 19948 35048 19988 35057
rect 19852 34208 19892 34217
rect 19852 32024 19892 34168
rect 19948 33872 19988 35008
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 19948 33823 19988 33832
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 19852 31975 19892 31984
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 20524 28412 20564 77512
rect 20716 76880 20756 84568
rect 21388 82088 21428 82097
rect 20812 78560 20852 78569
rect 20812 77972 20852 78520
rect 20812 77923 20852 77932
rect 20620 76840 20756 76880
rect 20620 32780 20660 76840
rect 21388 72848 21428 82048
rect 21388 72799 21428 72808
rect 20716 68732 20756 68741
rect 20716 46388 20756 68692
rect 20812 57224 20852 57233
rect 20812 52352 20852 57184
rect 21388 54200 21428 54209
rect 20812 52303 20852 52312
rect 21292 53444 21332 53453
rect 20812 50168 20852 50177
rect 20812 48908 20852 50128
rect 20812 48859 20852 48868
rect 21292 48488 21332 53404
rect 21292 48439 21332 48448
rect 20716 46339 20756 46348
rect 21388 46304 21428 54160
rect 21388 46255 21428 46264
rect 20716 35384 20756 35393
rect 20716 33956 20756 35344
rect 20716 33907 20756 33916
rect 21388 33704 21428 33713
rect 21388 33200 21428 33664
rect 21388 33151 21428 33160
rect 20620 32740 20948 32780
rect 20716 32360 20756 32369
rect 20620 30344 20660 30353
rect 20620 28580 20660 30304
rect 20716 30092 20756 32320
rect 20716 30043 20756 30052
rect 20620 28531 20660 28540
rect 20524 28372 20852 28412
rect 19756 28195 19796 28204
rect 20716 28244 20756 28253
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 19372 23575 19412 23584
rect 19468 27572 19508 27581
rect 19276 20971 19316 20980
rect 19372 23288 19412 23297
rect 19276 20264 19316 20273
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 18700 16736 18740 16745
rect 18700 10016 18740 16696
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 19276 16400 19316 20224
rect 19276 16351 19316 16360
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 19276 13796 19316 13805
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 18700 9967 18740 9976
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 19276 8000 19316 13756
rect 19372 9512 19412 23248
rect 19468 18080 19508 27532
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 19755 26144 19797 26153
rect 19755 26104 19756 26144
rect 19796 26104 19797 26144
rect 19755 26095 19797 26104
rect 19756 26010 19796 26095
rect 20524 25976 20564 25985
rect 19564 25892 19604 25901
rect 19564 24800 19604 25852
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 19564 24751 19604 24760
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 19660 22868 19700 22877
rect 19468 18031 19508 18040
rect 19564 20348 19604 20357
rect 19564 14468 19604 20308
rect 19660 16988 19700 22828
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 19660 16939 19700 16948
rect 19948 19844 19988 19853
rect 19564 14419 19604 14428
rect 19852 14384 19892 14393
rect 19372 9463 19412 9472
rect 19468 9848 19508 9857
rect 19468 8840 19508 9808
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 19276 6992 19316 7960
rect 19372 8800 19508 8840
rect 19564 9512 19604 9521
rect 19372 7748 19412 8800
rect 19372 7699 19412 7708
rect 19468 8672 19508 8681
rect 19276 6943 19316 6952
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19468 5480 19508 8632
rect 19564 6992 19604 9472
rect 19564 6943 19604 6952
rect 19852 6152 19892 14344
rect 19948 13292 19988 19804
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 20524 18752 20564 25936
rect 20524 18703 20564 18712
rect 20620 21608 20660 21617
rect 20524 18584 20564 18593
rect 20524 18332 20564 18544
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 20139 15560 20181 15569
rect 20139 15520 20140 15560
rect 20180 15520 20181 15560
rect 20139 15511 20181 15520
rect 20140 15426 20180 15511
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 19948 13243 19988 13252
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 20048 11360 20416 11369
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 20139 11192 20181 11201
rect 20139 11152 20140 11192
rect 20180 11152 20181 11192
rect 20139 11143 20181 11152
rect 20140 11058 20180 11143
rect 20524 9932 20564 18292
rect 20620 17324 20660 21568
rect 20620 17275 20660 17284
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 20524 9176 20564 9892
rect 20524 9127 20564 9136
rect 20139 8840 20181 8849
rect 20139 8800 20140 8840
rect 20180 8800 20181 8840
rect 20139 8791 20181 8800
rect 20140 8706 20180 8791
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 20139 7160 20181 7169
rect 20139 7120 20140 7160
rect 20180 7120 20181 7160
rect 20139 7111 20181 7120
rect 20140 7026 20180 7111
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 19852 6103 19892 6112
rect 19468 5431 19508 5440
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 20716 5060 20756 28204
rect 20812 19508 20852 28372
rect 20908 25052 20948 32740
rect 20908 25003 20948 25012
rect 21004 27488 21044 27497
rect 20812 19459 20852 19468
rect 20908 24548 20948 24557
rect 20811 16820 20853 16829
rect 20811 16780 20812 16820
rect 20852 16780 20853 16820
rect 20811 16771 20853 16780
rect 20812 15224 20852 16771
rect 20812 15175 20852 15184
rect 20811 10016 20853 10025
rect 20811 9976 20812 10016
rect 20852 9976 20853 10016
rect 20811 9967 20853 9976
rect 20812 9848 20852 9967
rect 20812 9799 20852 9808
rect 20908 9176 20948 24508
rect 21004 21524 21044 27448
rect 21004 18752 21044 21484
rect 21196 24380 21236 24389
rect 21004 18703 21044 18712
rect 21100 18920 21140 18929
rect 21004 18584 21044 18593
rect 21004 16232 21044 18544
rect 21100 16316 21140 18880
rect 21100 16267 21140 16276
rect 21004 16183 21044 16192
rect 21196 11864 21236 24340
rect 21196 11815 21236 11824
rect 20908 9127 20948 9136
rect 20716 5011 20756 5020
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 18604 2071 18644 2080
rect 19563 2120 19605 2129
rect 19563 2080 19564 2120
rect 19604 2080 19605 2120
rect 19563 2071 19605 2080
rect 19564 1986 19604 2071
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 18412 1231 18452 1240
rect 16108 1147 16148 1156
rect 15532 1063 15572 1072
rect 19179 944 19221 953
rect 19179 904 19180 944
rect 19220 904 19221 944
rect 19179 895 19221 904
rect 19180 810 19220 895
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 13516 55 13556 64
<< via4 >>
rect 19084 85912 19124 85952
rect 19276 85744 19316 85784
rect 1516 83476 1556 83516
rect 652 76504 692 76544
rect 76 42652 116 42692
rect 268 42736 308 42776
rect 1036 59872 1076 59912
rect 172 40552 212 40592
rect 460 34168 500 34208
rect 556 33664 596 33704
rect 556 22072 596 22112
rect 748 22072 788 22112
rect 652 16360 692 16400
rect 940 16780 980 16820
rect 1324 34336 1364 34376
rect 1228 33496 1268 33536
rect 1420 26272 1460 26312
rect 1324 26104 1364 26144
rect 1228 21400 1268 21440
rect 1228 18712 1268 18752
rect 1228 18292 1268 18332
rect 3688 84652 3728 84692
rect 3770 84652 3810 84692
rect 3852 84652 3892 84692
rect 3934 84652 3974 84692
rect 4016 84652 4056 84692
rect 4928 83896 4968 83936
rect 5010 83896 5050 83936
rect 5092 83896 5132 83936
rect 5174 83896 5214 83936
rect 5256 83896 5296 83936
rect 3688 83140 3728 83180
rect 3770 83140 3810 83180
rect 3852 83140 3892 83180
rect 3934 83140 3974 83180
rect 4016 83140 4056 83180
rect 2380 45928 2420 45968
rect 2860 51976 2900 52016
rect 3148 51976 3188 52016
rect 2956 16360 2996 16400
rect 2668 8800 2708 8840
rect 3436 57856 3476 57896
rect 4928 82384 4968 82424
rect 5010 82384 5050 82424
rect 5092 82384 5132 82424
rect 5174 82384 5214 82424
rect 5256 82384 5296 82424
rect 3688 81628 3728 81668
rect 3770 81628 3810 81668
rect 3852 81628 3892 81668
rect 3934 81628 3974 81668
rect 4016 81628 4056 81668
rect 4928 80872 4968 80912
rect 5010 80872 5050 80912
rect 5092 80872 5132 80912
rect 5174 80872 5214 80912
rect 5256 80872 5296 80912
rect 3688 80116 3728 80156
rect 3770 80116 3810 80156
rect 3852 80116 3892 80156
rect 3934 80116 3974 80156
rect 4016 80116 4056 80156
rect 4928 79360 4968 79400
rect 5010 79360 5050 79400
rect 5092 79360 5132 79400
rect 5174 79360 5214 79400
rect 5256 79360 5296 79400
rect 3688 78604 3728 78644
rect 3770 78604 3810 78644
rect 3852 78604 3892 78644
rect 3934 78604 3974 78644
rect 4016 78604 4056 78644
rect 4928 77848 4968 77888
rect 5010 77848 5050 77888
rect 5092 77848 5132 77888
rect 5174 77848 5214 77888
rect 5256 77848 5296 77888
rect 3688 77092 3728 77132
rect 3770 77092 3810 77132
rect 3852 77092 3892 77132
rect 3934 77092 3974 77132
rect 4016 77092 4056 77132
rect 4928 76336 4968 76376
rect 5010 76336 5050 76376
rect 5092 76336 5132 76376
rect 5174 76336 5214 76376
rect 5256 76336 5296 76376
rect 3688 75580 3728 75620
rect 3770 75580 3810 75620
rect 3852 75580 3892 75620
rect 3934 75580 3974 75620
rect 4016 75580 4056 75620
rect 4928 74824 4968 74864
rect 5010 74824 5050 74864
rect 5092 74824 5132 74864
rect 5174 74824 5214 74864
rect 5256 74824 5296 74864
rect 3688 74068 3728 74108
rect 3770 74068 3810 74108
rect 3852 74068 3892 74108
rect 3934 74068 3974 74108
rect 4016 74068 4056 74108
rect 4928 73312 4968 73352
rect 5010 73312 5050 73352
rect 5092 73312 5132 73352
rect 5174 73312 5214 73352
rect 5256 73312 5296 73352
rect 3688 72556 3728 72596
rect 3770 72556 3810 72596
rect 3852 72556 3892 72596
rect 3934 72556 3974 72596
rect 4016 72556 4056 72596
rect 3688 71044 3728 71084
rect 3770 71044 3810 71084
rect 3852 71044 3892 71084
rect 3934 71044 3974 71084
rect 4016 71044 4056 71084
rect 3688 69532 3728 69572
rect 3770 69532 3810 69572
rect 3852 69532 3892 69572
rect 3934 69532 3974 69572
rect 4016 69532 4056 69572
rect 3688 68020 3728 68060
rect 3770 68020 3810 68060
rect 3852 68020 3892 68060
rect 3934 68020 3974 68060
rect 4016 68020 4056 68060
rect 3688 66508 3728 66548
rect 3770 66508 3810 66548
rect 3852 66508 3892 66548
rect 3934 66508 3974 66548
rect 4016 66508 4056 66548
rect 4928 71800 4968 71840
rect 5010 71800 5050 71840
rect 5092 71800 5132 71840
rect 5174 71800 5214 71840
rect 5256 71800 5296 71840
rect 4928 70288 4968 70328
rect 5010 70288 5050 70328
rect 5092 70288 5132 70328
rect 5174 70288 5214 70328
rect 5256 70288 5296 70328
rect 4928 68776 4968 68816
rect 5010 68776 5050 68816
rect 5092 68776 5132 68816
rect 5174 68776 5214 68816
rect 5256 68776 5296 68816
rect 4928 67264 4968 67304
rect 5010 67264 5050 67304
rect 5092 67264 5132 67304
rect 5174 67264 5214 67304
rect 5256 67264 5296 67304
rect 3688 64996 3728 65036
rect 3770 64996 3810 65036
rect 3852 64996 3892 65036
rect 3934 64996 3974 65036
rect 4016 64996 4056 65036
rect 3688 63484 3728 63524
rect 3770 63484 3810 63524
rect 3852 63484 3892 63524
rect 3934 63484 3974 63524
rect 4016 63484 4056 63524
rect 3688 61972 3728 62012
rect 3770 61972 3810 62012
rect 3852 61972 3892 62012
rect 3934 61972 3974 62012
rect 4016 61972 4056 62012
rect 3688 60460 3728 60500
rect 3770 60460 3810 60500
rect 3852 60460 3892 60500
rect 3934 60460 3974 60500
rect 4016 60460 4056 60500
rect 4928 65752 4968 65792
rect 5010 65752 5050 65792
rect 5092 65752 5132 65792
rect 5174 65752 5214 65792
rect 5256 65752 5296 65792
rect 4928 64240 4968 64280
rect 5010 64240 5050 64280
rect 5092 64240 5132 64280
rect 5174 64240 5214 64280
rect 5256 64240 5296 64280
rect 4928 62728 4968 62768
rect 5010 62728 5050 62768
rect 5092 62728 5132 62768
rect 5174 62728 5214 62768
rect 5256 62728 5296 62768
rect 4928 61216 4968 61256
rect 5010 61216 5050 61256
rect 5092 61216 5132 61256
rect 5174 61216 5214 61256
rect 5256 61216 5296 61256
rect 3688 58948 3728 58988
rect 3770 58948 3810 58988
rect 3852 58948 3892 58988
rect 3934 58948 3974 58988
rect 4016 58948 4056 58988
rect 3688 57436 3728 57476
rect 3770 57436 3810 57476
rect 3852 57436 3892 57476
rect 3934 57436 3974 57476
rect 4016 57436 4056 57476
rect 3532 56848 3572 56888
rect 3688 55924 3728 55964
rect 3770 55924 3810 55964
rect 3852 55924 3892 55964
rect 3934 55924 3974 55964
rect 4016 55924 4056 55964
rect 3688 54412 3728 54452
rect 3770 54412 3810 54452
rect 3852 54412 3892 54452
rect 3934 54412 3974 54452
rect 4016 54412 4056 54452
rect 3688 52900 3728 52940
rect 3770 52900 3810 52940
rect 3852 52900 3892 52940
rect 3934 52900 3974 52940
rect 4016 52900 4056 52940
rect 3688 51388 3728 51428
rect 3770 51388 3810 51428
rect 3852 51388 3892 51428
rect 3934 51388 3974 51428
rect 4016 51388 4056 51428
rect 3688 49876 3728 49916
rect 3770 49876 3810 49916
rect 3852 49876 3892 49916
rect 3934 49876 3974 49916
rect 4016 49876 4056 49916
rect 3688 48364 3728 48404
rect 3770 48364 3810 48404
rect 3852 48364 3892 48404
rect 3934 48364 3974 48404
rect 4016 48364 4056 48404
rect 3688 46852 3728 46892
rect 3770 46852 3810 46892
rect 3852 46852 3892 46892
rect 3934 46852 3974 46892
rect 4016 46852 4056 46892
rect 3688 45340 3728 45380
rect 3770 45340 3810 45380
rect 3852 45340 3892 45380
rect 3934 45340 3974 45380
rect 4016 45340 4056 45380
rect 3688 43828 3728 43868
rect 3770 43828 3810 43868
rect 3852 43828 3892 43868
rect 3934 43828 3974 43868
rect 4016 43828 4056 43868
rect 3688 42316 3728 42356
rect 3770 42316 3810 42356
rect 3852 42316 3892 42356
rect 3934 42316 3974 42356
rect 4016 42316 4056 42356
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 4928 59704 4968 59744
rect 5010 59704 5050 59744
rect 5092 59704 5132 59744
rect 5174 59704 5214 59744
rect 5256 59704 5296 59744
rect 4928 58192 4968 58232
rect 5010 58192 5050 58232
rect 5092 58192 5132 58232
rect 5174 58192 5214 58232
rect 5256 58192 5296 58232
rect 4300 51808 4340 51848
rect 4928 56680 4968 56720
rect 5010 56680 5050 56720
rect 5092 56680 5132 56720
rect 5174 56680 5214 56720
rect 5256 56680 5296 56720
rect 4928 55168 4968 55208
rect 5010 55168 5050 55208
rect 5092 55168 5132 55208
rect 5174 55168 5214 55208
rect 5256 55168 5296 55208
rect 4928 53656 4968 53696
rect 5010 53656 5050 53696
rect 5092 53656 5132 53696
rect 5174 53656 5214 53696
rect 5256 53656 5296 53696
rect 4928 52144 4968 52184
rect 5010 52144 5050 52184
rect 5092 52144 5132 52184
rect 5174 52144 5214 52184
rect 5256 52144 5296 52184
rect 4928 50632 4968 50672
rect 5010 50632 5050 50672
rect 5092 50632 5132 50672
rect 5174 50632 5214 50672
rect 5256 50632 5296 50672
rect 4588 45676 4628 45716
rect 4928 49120 4968 49160
rect 5010 49120 5050 49160
rect 5092 49120 5132 49160
rect 5174 49120 5214 49160
rect 5256 49120 5296 49160
rect 4928 47608 4968 47648
rect 5010 47608 5050 47648
rect 5092 47608 5132 47648
rect 5174 47608 5214 47648
rect 5256 47608 5296 47648
rect 4928 46096 4968 46136
rect 5010 46096 5050 46136
rect 5092 46096 5132 46136
rect 5174 46096 5214 46136
rect 5256 46096 5296 46136
rect 4684 44920 4724 44960
rect 4928 44584 4968 44624
rect 5010 44584 5050 44624
rect 5092 44584 5132 44624
rect 5174 44584 5214 44624
rect 5256 44584 5296 44624
rect 4928 43072 4968 43112
rect 5010 43072 5050 43112
rect 5092 43072 5132 43112
rect 5174 43072 5214 43112
rect 5256 43072 5296 43112
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 4492 35008 4532 35048
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 5356 35176 5396 35216
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 5548 40552 5588 40592
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 3724 18544 3764 18584
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 5068 17704 5108 17744
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 4876 16360 4916 16400
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 3436 12496 3476 12536
rect 3820 12496 3860 12536
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3724 8884 3764 8924
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 4204 8884 4244 8924
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 5836 35176 5876 35216
rect 5932 26272 5972 26312
rect 5548 9976 5588 10016
rect 6316 16780 6356 16820
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 5740 2080 5780 2120
rect 6796 84400 6836 84440
rect 6796 68020 6836 68060
rect 6604 42736 6644 42776
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 7276 53236 7316 53276
rect 7948 57940 7988 57980
rect 7564 34168 7604 34208
rect 7276 2080 7316 2120
rect 8524 76672 8564 76712
rect 8236 35008 8276 35048
rect 7948 18712 7988 18752
rect 7852 1240 7892 1280
rect 8428 18292 8468 18332
rect 9004 76672 9044 76712
rect 8620 14512 8660 14552
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 9004 17536 9044 17576
rect 9004 13168 9044 13208
rect 5068 232 5108 272
rect 8908 232 8948 272
rect 4876 148 4916 188
rect 3340 64 3380 104
rect 9292 17536 9332 17576
rect 10060 57940 10100 57980
rect 10156 41896 10196 41936
rect 9292 13168 9332 13208
rect 9676 18544 9716 18584
rect 9964 10228 10004 10268
rect 10732 57856 10772 57896
rect 10732 42652 10772 42692
rect 10444 21400 10484 21440
rect 10732 11236 10772 11276
rect 11212 72220 11252 72260
rect 11308 68020 11348 68060
rect 11500 56848 11540 56888
rect 11404 44920 11444 44960
rect 11308 17704 11348 17744
rect 13228 75916 13268 75956
rect 12652 59872 12692 59912
rect 12076 10396 12116 10436
rect 12556 33664 12596 33704
rect 13132 15688 13172 15728
rect 13036 11068 13076 11108
rect 13420 1156 13460 1196
rect 9100 64 9140 104
rect 13804 2668 13844 2708
rect 14284 47860 14324 47900
rect 15052 84400 15092 84440
rect 14764 7120 14804 7160
rect 15148 14512 15188 14552
rect 15724 17620 15764 17660
rect 15724 16780 15764 16820
rect 16396 15520 16436 15560
rect 17932 85072 17972 85112
rect 18808 84652 18848 84692
rect 18890 84652 18930 84692
rect 18972 84652 19012 84692
rect 19054 84652 19094 84692
rect 19136 84652 19176 84692
rect 16972 53236 17012 53276
rect 17068 33496 17108 33536
rect 17068 28456 17108 28496
rect 17260 28456 17300 28496
rect 17644 51808 17684 51848
rect 17644 29380 17684 29420
rect 18028 45676 18068 45716
rect 17932 29380 17972 29420
rect 18316 24592 18356 24632
rect 18220 10396 18260 10436
rect 18808 83140 18848 83180
rect 18890 83140 18930 83180
rect 18972 83140 19012 83180
rect 19054 83140 19094 83180
rect 19136 83140 19176 83180
rect 18808 81628 18848 81668
rect 18890 81628 18930 81668
rect 18972 81628 19012 81668
rect 19054 81628 19094 81668
rect 19136 81628 19176 81668
rect 18808 80116 18848 80156
rect 18890 80116 18930 80156
rect 18972 80116 19012 80156
rect 19054 80116 19094 80156
rect 19136 80116 19176 80156
rect 18808 78604 18848 78644
rect 18890 78604 18930 78644
rect 18972 78604 19012 78644
rect 19054 78604 19094 78644
rect 19136 78604 19176 78644
rect 18808 77092 18848 77132
rect 18890 77092 18930 77132
rect 18972 77092 19012 77132
rect 19054 77092 19094 77132
rect 19136 77092 19176 77132
rect 18892 75916 18932 75956
rect 18808 75580 18848 75620
rect 18890 75580 18930 75620
rect 18972 75580 19012 75620
rect 19054 75580 19094 75620
rect 19136 75580 19176 75620
rect 18808 74068 18848 74108
rect 18890 74068 18930 74108
rect 18972 74068 19012 74108
rect 19054 74068 19094 74108
rect 19136 74068 19176 74108
rect 18808 72556 18848 72596
rect 18890 72556 18930 72596
rect 18972 72556 19012 72596
rect 19054 72556 19094 72596
rect 19136 72556 19176 72596
rect 18808 71044 18848 71084
rect 18890 71044 18930 71084
rect 18972 71044 19012 71084
rect 19054 71044 19094 71084
rect 19136 71044 19176 71084
rect 18808 69532 18848 69572
rect 18890 69532 18930 69572
rect 18972 69532 19012 69572
rect 19054 69532 19094 69572
rect 19136 69532 19176 69572
rect 18808 68020 18848 68060
rect 18890 68020 18930 68060
rect 18972 68020 19012 68060
rect 19054 68020 19094 68060
rect 19136 68020 19176 68060
rect 18808 66508 18848 66548
rect 18890 66508 18930 66548
rect 18972 66508 19012 66548
rect 19054 66508 19094 66548
rect 19136 66508 19176 66548
rect 18808 64996 18848 65036
rect 18890 64996 18930 65036
rect 18972 64996 19012 65036
rect 19054 64996 19094 65036
rect 19136 64996 19176 65036
rect 18808 63484 18848 63524
rect 18890 63484 18930 63524
rect 18972 63484 19012 63524
rect 19054 63484 19094 63524
rect 19136 63484 19176 63524
rect 18808 61972 18848 62012
rect 18890 61972 18930 62012
rect 18972 61972 19012 62012
rect 19054 61972 19094 62012
rect 19136 61972 19176 62012
rect 18808 60460 18848 60500
rect 18890 60460 18930 60500
rect 18972 60460 19012 60500
rect 19054 60460 19094 60500
rect 19136 60460 19176 60500
rect 18808 58948 18848 58988
rect 18890 58948 18930 58988
rect 18972 58948 19012 58988
rect 19054 58948 19094 58988
rect 19136 58948 19176 58988
rect 18808 57436 18848 57476
rect 18890 57436 18930 57476
rect 18972 57436 19012 57476
rect 19054 57436 19094 57476
rect 19136 57436 19176 57476
rect 18808 55924 18848 55964
rect 18890 55924 18930 55964
rect 18972 55924 19012 55964
rect 19054 55924 19094 55964
rect 19136 55924 19176 55964
rect 18808 54412 18848 54452
rect 18890 54412 18930 54452
rect 18972 54412 19012 54452
rect 19054 54412 19094 54452
rect 19136 54412 19176 54452
rect 18700 53236 18740 53276
rect 18808 52900 18848 52940
rect 18890 52900 18930 52940
rect 18972 52900 19012 52940
rect 19054 52900 19094 52940
rect 19136 52900 19176 52940
rect 20048 83896 20088 83936
rect 20130 83896 20170 83936
rect 20212 83896 20252 83936
rect 20294 83896 20334 83936
rect 20376 83896 20416 83936
rect 20048 82384 20088 82424
rect 20130 82384 20170 82424
rect 20212 82384 20252 82424
rect 20294 82384 20334 82424
rect 20376 82384 20416 82424
rect 20048 80872 20088 80912
rect 20130 80872 20170 80912
rect 20212 80872 20252 80912
rect 20294 80872 20334 80912
rect 20376 80872 20416 80912
rect 20048 79360 20088 79400
rect 20130 79360 20170 79400
rect 20212 79360 20252 79400
rect 20294 79360 20334 79400
rect 20376 79360 20416 79400
rect 20048 77848 20088 77888
rect 20130 77848 20170 77888
rect 20212 77848 20252 77888
rect 20294 77848 20334 77888
rect 20376 77848 20416 77888
rect 20048 76336 20088 76376
rect 20130 76336 20170 76376
rect 20212 76336 20252 76376
rect 20294 76336 20334 76376
rect 20376 76336 20416 76376
rect 20048 74824 20088 74864
rect 20130 74824 20170 74864
rect 20212 74824 20252 74864
rect 20294 74824 20334 74864
rect 20376 74824 20416 74864
rect 20048 73312 20088 73352
rect 20130 73312 20170 73352
rect 20212 73312 20252 73352
rect 20294 73312 20334 73352
rect 20376 73312 20416 73352
rect 19756 72220 19796 72260
rect 20048 71800 20088 71840
rect 20130 71800 20170 71840
rect 20212 71800 20252 71840
rect 20294 71800 20334 71840
rect 20376 71800 20416 71840
rect 20048 70288 20088 70328
rect 20130 70288 20170 70328
rect 20212 70288 20252 70328
rect 20294 70288 20334 70328
rect 20376 70288 20416 70328
rect 20048 68776 20088 68816
rect 20130 68776 20170 68816
rect 20212 68776 20252 68816
rect 20294 68776 20334 68816
rect 20376 68776 20416 68816
rect 20048 67264 20088 67304
rect 20130 67264 20170 67304
rect 20212 67264 20252 67304
rect 20294 67264 20334 67304
rect 20376 67264 20416 67304
rect 20048 65752 20088 65792
rect 20130 65752 20170 65792
rect 20212 65752 20252 65792
rect 20294 65752 20334 65792
rect 20376 65752 20416 65792
rect 18808 51388 18848 51428
rect 18890 51388 18930 51428
rect 18972 51388 19012 51428
rect 19054 51388 19094 51428
rect 19136 51388 19176 51428
rect 18808 49876 18848 49916
rect 18890 49876 18930 49916
rect 18972 49876 19012 49916
rect 19054 49876 19094 49916
rect 19136 49876 19176 49916
rect 18808 48364 18848 48404
rect 18890 48364 18930 48404
rect 18972 48364 19012 48404
rect 19054 48364 19094 48404
rect 19136 48364 19176 48404
rect 18808 46852 18848 46892
rect 18890 46852 18930 46892
rect 18972 46852 19012 46892
rect 19054 46852 19094 46892
rect 19136 46852 19176 46892
rect 18808 45340 18848 45380
rect 18890 45340 18930 45380
rect 18972 45340 19012 45380
rect 19054 45340 19094 45380
rect 19136 45340 19176 45380
rect 18808 43828 18848 43868
rect 18890 43828 18930 43868
rect 18972 43828 19012 43868
rect 19054 43828 19094 43868
rect 19136 43828 19176 43868
rect 18808 42316 18848 42356
rect 18890 42316 18930 42356
rect 18972 42316 19012 42356
rect 19054 42316 19094 42356
rect 19136 42316 19176 42356
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 20048 64240 20088 64280
rect 20130 64240 20170 64280
rect 20212 64240 20252 64280
rect 20294 64240 20334 64280
rect 20376 64240 20416 64280
rect 20048 62728 20088 62768
rect 20130 62728 20170 62768
rect 20212 62728 20252 62768
rect 20294 62728 20334 62768
rect 20376 62728 20416 62768
rect 20048 61216 20088 61256
rect 20130 61216 20170 61256
rect 20212 61216 20252 61256
rect 20294 61216 20334 61256
rect 20376 61216 20416 61256
rect 20048 59704 20088 59744
rect 20130 59704 20170 59744
rect 20212 59704 20252 59744
rect 20294 59704 20334 59744
rect 20376 59704 20416 59744
rect 20048 58192 20088 58232
rect 20130 58192 20170 58232
rect 20212 58192 20252 58232
rect 20294 58192 20334 58232
rect 20376 58192 20416 58232
rect 20048 56680 20088 56720
rect 20130 56680 20170 56720
rect 20212 56680 20252 56720
rect 20294 56680 20334 56720
rect 20376 56680 20416 56720
rect 20048 55168 20088 55208
rect 20130 55168 20170 55208
rect 20212 55168 20252 55208
rect 20294 55168 20334 55208
rect 20376 55168 20416 55208
rect 20048 53656 20088 53696
rect 20130 53656 20170 53696
rect 20212 53656 20252 53696
rect 20294 53656 20334 53696
rect 20376 53656 20416 53696
rect 20140 53152 20180 53192
rect 20048 52144 20088 52184
rect 20130 52144 20170 52184
rect 20212 52144 20252 52184
rect 20294 52144 20334 52184
rect 20376 52144 20416 52184
rect 20048 50632 20088 50672
rect 20130 50632 20170 50672
rect 20212 50632 20252 50672
rect 20294 50632 20334 50672
rect 20376 50632 20416 50672
rect 20048 49120 20088 49160
rect 20130 49120 20170 49160
rect 20212 49120 20252 49160
rect 20294 49120 20334 49160
rect 20376 49120 20416 49160
rect 20048 47608 20088 47648
rect 20130 47608 20170 47648
rect 20212 47608 20252 47648
rect 20294 47608 20334 47648
rect 20376 47608 20416 47648
rect 20048 46096 20088 46136
rect 20130 46096 20170 46136
rect 20212 46096 20252 46136
rect 20294 46096 20334 46136
rect 20376 46096 20416 46136
rect 20048 44584 20088 44624
rect 20130 44584 20170 44624
rect 20212 44584 20252 44624
rect 20294 44584 20334 44624
rect 20376 44584 20416 44624
rect 20048 43072 20088 43112
rect 20130 43072 20170 43112
rect 20212 43072 20252 43112
rect 20294 43072 20334 43112
rect 20376 43072 20416 43112
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 19756 26104 19796 26144
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 20140 15520 20180 15560
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 20140 11152 20180 11192
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 20140 8800 20180 8840
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 20140 7120 20180 7160
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20812 16780 20852 16820
rect 20812 9976 20852 10016
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 19564 2080 19604 2120
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 19180 904 19220 944
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal5 >>
rect 15100 85912 19084 85952
rect 19124 85912 19133 85952
rect 12122 85891 12246 85910
rect 12122 85805 12141 85891
rect 12227 85868 12246 85891
rect 15100 85868 15140 85912
rect 12227 85828 15140 85868
rect 12227 85805 12246 85828
rect 12122 85786 12246 85805
rect 17138 85807 17262 85826
rect 17138 85721 17157 85807
rect 17243 85784 17262 85807
rect 17243 85744 19276 85784
rect 19316 85744 19325 85784
rect 17243 85721 17262 85744
rect 17138 85702 17262 85721
rect 16226 85135 16350 85154
rect 16226 85049 16245 85135
rect 16331 85112 16350 85135
rect 16331 85072 17932 85112
rect 17972 85072 17981 85112
rect 16331 85049 16350 85072
rect 16226 85030 16350 85049
rect 3679 84715 4065 84734
rect 3679 84692 3745 84715
rect 3831 84692 3913 84715
rect 3999 84692 4065 84715
rect 3679 84652 3688 84692
rect 3728 84652 3745 84692
rect 3831 84652 3852 84692
rect 3892 84652 3913 84692
rect 3999 84652 4016 84692
rect 4056 84652 4065 84692
rect 3679 84629 3745 84652
rect 3831 84629 3913 84652
rect 3999 84629 4065 84652
rect 3679 84610 4065 84629
rect 18799 84715 19185 84734
rect 18799 84692 18865 84715
rect 18951 84692 19033 84715
rect 19119 84692 19185 84715
rect 18799 84652 18808 84692
rect 18848 84652 18865 84692
rect 18951 84652 18972 84692
rect 19012 84652 19033 84692
rect 19119 84652 19136 84692
rect 19176 84652 19185 84692
rect 18799 84629 18865 84652
rect 18951 84629 19033 84652
rect 19119 84629 19185 84652
rect 18799 84610 19185 84629
rect 7106 84463 7230 84482
rect 7106 84440 7125 84463
rect 6787 84400 6796 84440
rect 6836 84400 7125 84440
rect 7106 84377 7125 84400
rect 7211 84377 7230 84463
rect 7106 84358 7230 84377
rect 14858 84463 14982 84482
rect 14858 84377 14877 84463
rect 14963 84440 14982 84463
rect 14963 84400 15052 84440
rect 15092 84400 15101 84440
rect 14963 84377 14982 84400
rect 14858 84358 14982 84377
rect 4919 83959 5305 83978
rect 4919 83936 4985 83959
rect 5071 83936 5153 83959
rect 5239 83936 5305 83959
rect 4919 83896 4928 83936
rect 4968 83896 4985 83936
rect 5071 83896 5092 83936
rect 5132 83896 5153 83936
rect 5239 83896 5256 83936
rect 5296 83896 5305 83936
rect 4919 83873 4985 83896
rect 5071 83873 5153 83896
rect 5239 83873 5305 83896
rect 4919 83854 5305 83873
rect 20039 83959 20425 83978
rect 20039 83936 20105 83959
rect 20191 83936 20273 83959
rect 20359 83936 20425 83959
rect 20039 83896 20048 83936
rect 20088 83896 20105 83936
rect 20191 83896 20212 83936
rect 20252 83896 20273 83936
rect 20359 83896 20376 83936
rect 20416 83896 20425 83936
rect 20039 83873 20105 83896
rect 20191 83873 20273 83896
rect 20359 83873 20425 83896
rect 20039 83854 20425 83873
rect 2090 83539 2214 83558
rect 2090 83516 2109 83539
rect 1507 83476 1516 83516
rect 1556 83476 2109 83516
rect 2090 83453 2109 83476
rect 2195 83453 2214 83539
rect 2090 83434 2214 83453
rect 3679 83203 4065 83222
rect 3679 83180 3745 83203
rect 3831 83180 3913 83203
rect 3999 83180 4065 83203
rect 3679 83140 3688 83180
rect 3728 83140 3745 83180
rect 3831 83140 3852 83180
rect 3892 83140 3913 83180
rect 3999 83140 4016 83180
rect 4056 83140 4065 83180
rect 3679 83117 3745 83140
rect 3831 83117 3913 83140
rect 3999 83117 4065 83140
rect 3679 83098 4065 83117
rect 18799 83203 19185 83222
rect 18799 83180 18865 83203
rect 18951 83180 19033 83203
rect 19119 83180 19185 83203
rect 18799 83140 18808 83180
rect 18848 83140 18865 83180
rect 18951 83140 18972 83180
rect 19012 83140 19033 83180
rect 19119 83140 19136 83180
rect 19176 83140 19185 83180
rect 18799 83117 18865 83140
rect 18951 83117 19033 83140
rect 19119 83117 19185 83140
rect 18799 83098 19185 83117
rect 4919 82447 5305 82466
rect 4919 82424 4985 82447
rect 5071 82424 5153 82447
rect 5239 82424 5305 82447
rect 4919 82384 4928 82424
rect 4968 82384 4985 82424
rect 5071 82384 5092 82424
rect 5132 82384 5153 82424
rect 5239 82384 5256 82424
rect 5296 82384 5305 82424
rect 4919 82361 4985 82384
rect 5071 82361 5153 82384
rect 5239 82361 5305 82384
rect 4919 82342 5305 82361
rect 20039 82447 20425 82466
rect 20039 82424 20105 82447
rect 20191 82424 20273 82447
rect 20359 82424 20425 82447
rect 20039 82384 20048 82424
rect 20088 82384 20105 82424
rect 20191 82384 20212 82424
rect 20252 82384 20273 82424
rect 20359 82384 20376 82424
rect 20416 82384 20425 82424
rect 20039 82361 20105 82384
rect 20191 82361 20273 82384
rect 20359 82361 20425 82384
rect 20039 82342 20425 82361
rect 3679 81691 4065 81710
rect 3679 81668 3745 81691
rect 3831 81668 3913 81691
rect 3999 81668 4065 81691
rect 3679 81628 3688 81668
rect 3728 81628 3745 81668
rect 3831 81628 3852 81668
rect 3892 81628 3913 81668
rect 3999 81628 4016 81668
rect 4056 81628 4065 81668
rect 3679 81605 3745 81628
rect 3831 81605 3913 81628
rect 3999 81605 4065 81628
rect 3679 81586 4065 81605
rect 18799 81691 19185 81710
rect 18799 81668 18865 81691
rect 18951 81668 19033 81691
rect 19119 81668 19185 81691
rect 18799 81628 18808 81668
rect 18848 81628 18865 81668
rect 18951 81628 18972 81668
rect 19012 81628 19033 81668
rect 19119 81628 19136 81668
rect 19176 81628 19185 81668
rect 18799 81605 18865 81628
rect 18951 81605 19033 81628
rect 19119 81605 19185 81628
rect 18799 81586 19185 81605
rect 4919 80935 5305 80954
rect 4919 80912 4985 80935
rect 5071 80912 5153 80935
rect 5239 80912 5305 80935
rect 4919 80872 4928 80912
rect 4968 80872 4985 80912
rect 5071 80872 5092 80912
rect 5132 80872 5153 80912
rect 5239 80872 5256 80912
rect 5296 80872 5305 80912
rect 4919 80849 4985 80872
rect 5071 80849 5153 80872
rect 5239 80849 5305 80872
rect 4919 80830 5305 80849
rect 20039 80935 20425 80954
rect 20039 80912 20105 80935
rect 20191 80912 20273 80935
rect 20359 80912 20425 80935
rect 20039 80872 20048 80912
rect 20088 80872 20105 80912
rect 20191 80872 20212 80912
rect 20252 80872 20273 80912
rect 20359 80872 20376 80912
rect 20416 80872 20425 80912
rect 20039 80849 20105 80872
rect 20191 80849 20273 80872
rect 20359 80849 20425 80872
rect 20039 80830 20425 80849
rect 3679 80179 4065 80198
rect 3679 80156 3745 80179
rect 3831 80156 3913 80179
rect 3999 80156 4065 80179
rect 3679 80116 3688 80156
rect 3728 80116 3745 80156
rect 3831 80116 3852 80156
rect 3892 80116 3913 80156
rect 3999 80116 4016 80156
rect 4056 80116 4065 80156
rect 3679 80093 3745 80116
rect 3831 80093 3913 80116
rect 3999 80093 4065 80116
rect 3679 80074 4065 80093
rect 18799 80179 19185 80198
rect 18799 80156 18865 80179
rect 18951 80156 19033 80179
rect 19119 80156 19185 80179
rect 18799 80116 18808 80156
rect 18848 80116 18865 80156
rect 18951 80116 18972 80156
rect 19012 80116 19033 80156
rect 19119 80116 19136 80156
rect 19176 80116 19185 80156
rect 18799 80093 18865 80116
rect 18951 80093 19033 80116
rect 19119 80093 19185 80116
rect 18799 80074 19185 80093
rect 4919 79423 5305 79442
rect 4919 79400 4985 79423
rect 5071 79400 5153 79423
rect 5239 79400 5305 79423
rect 4919 79360 4928 79400
rect 4968 79360 4985 79400
rect 5071 79360 5092 79400
rect 5132 79360 5153 79400
rect 5239 79360 5256 79400
rect 5296 79360 5305 79400
rect 4919 79337 4985 79360
rect 5071 79337 5153 79360
rect 5239 79337 5305 79360
rect 4919 79318 5305 79337
rect 20039 79423 20425 79442
rect 20039 79400 20105 79423
rect 20191 79400 20273 79423
rect 20359 79400 20425 79423
rect 20039 79360 20048 79400
rect 20088 79360 20105 79400
rect 20191 79360 20212 79400
rect 20252 79360 20273 79400
rect 20359 79360 20376 79400
rect 20416 79360 20425 79400
rect 20039 79337 20105 79360
rect 20191 79337 20273 79360
rect 20359 79337 20425 79360
rect 20039 79318 20425 79337
rect 3679 78667 4065 78686
rect 3679 78644 3745 78667
rect 3831 78644 3913 78667
rect 3999 78644 4065 78667
rect 3679 78604 3688 78644
rect 3728 78604 3745 78644
rect 3831 78604 3852 78644
rect 3892 78604 3913 78644
rect 3999 78604 4016 78644
rect 4056 78604 4065 78644
rect 3679 78581 3745 78604
rect 3831 78581 3913 78604
rect 3999 78581 4065 78604
rect 3679 78562 4065 78581
rect 18799 78667 19185 78686
rect 18799 78644 18865 78667
rect 18951 78644 19033 78667
rect 19119 78644 19185 78667
rect 18799 78604 18808 78644
rect 18848 78604 18865 78644
rect 18951 78604 18972 78644
rect 19012 78604 19033 78644
rect 19119 78604 19136 78644
rect 19176 78604 19185 78644
rect 18799 78581 18865 78604
rect 18951 78581 19033 78604
rect 19119 78581 19185 78604
rect 18799 78562 19185 78581
rect 4919 77911 5305 77930
rect 4919 77888 4985 77911
rect 5071 77888 5153 77911
rect 5239 77888 5305 77911
rect 4919 77848 4928 77888
rect 4968 77848 4985 77888
rect 5071 77848 5092 77888
rect 5132 77848 5153 77888
rect 5239 77848 5256 77888
rect 5296 77848 5305 77888
rect 4919 77825 4985 77848
rect 5071 77825 5153 77848
rect 5239 77825 5305 77848
rect 4919 77806 5305 77825
rect 20039 77911 20425 77930
rect 20039 77888 20105 77911
rect 20191 77888 20273 77911
rect 20359 77888 20425 77911
rect 20039 77848 20048 77888
rect 20088 77848 20105 77888
rect 20191 77848 20212 77888
rect 20252 77848 20273 77888
rect 20359 77848 20376 77888
rect 20416 77848 20425 77888
rect 20039 77825 20105 77848
rect 20191 77825 20273 77848
rect 20359 77825 20425 77848
rect 20039 77806 20425 77825
rect 3679 77155 4065 77174
rect 3679 77132 3745 77155
rect 3831 77132 3913 77155
rect 3999 77132 4065 77155
rect 3679 77092 3688 77132
rect 3728 77092 3745 77132
rect 3831 77092 3852 77132
rect 3892 77092 3913 77132
rect 3999 77092 4016 77132
rect 4056 77092 4065 77132
rect 3679 77069 3745 77092
rect 3831 77069 3913 77092
rect 3999 77069 4065 77092
rect 3679 77050 4065 77069
rect 18799 77155 19185 77174
rect 18799 77132 18865 77155
rect 18951 77132 19033 77155
rect 19119 77132 19185 77155
rect 18799 77092 18808 77132
rect 18848 77092 18865 77132
rect 18951 77092 18972 77132
rect 19012 77092 19033 77132
rect 19119 77092 19136 77132
rect 19176 77092 19185 77132
rect 18799 77069 18865 77092
rect 18951 77069 19033 77092
rect 19119 77069 19185 77092
rect 18799 77050 19185 77069
rect 8474 76735 8598 76754
rect 8474 76649 8493 76735
rect 8579 76649 8598 76735
rect 9386 76735 9510 76754
rect 9386 76712 9405 76735
rect 8995 76672 9004 76712
rect 9044 76672 9405 76712
rect 8474 76630 8598 76649
rect 9386 76649 9405 76672
rect 9491 76649 9510 76735
rect 9386 76630 9510 76649
rect 1178 76567 1302 76586
rect 1178 76544 1197 76567
rect 643 76504 652 76544
rect 692 76504 1197 76544
rect 1178 76481 1197 76504
rect 1283 76481 1302 76567
rect 1178 76462 1302 76481
rect 4919 76399 5305 76418
rect 4919 76376 4985 76399
rect 5071 76376 5153 76399
rect 5239 76376 5305 76399
rect 4919 76336 4928 76376
rect 4968 76336 4985 76376
rect 5071 76336 5092 76376
rect 5132 76336 5153 76376
rect 5239 76336 5256 76376
rect 5296 76336 5305 76376
rect 4919 76313 4985 76336
rect 5071 76313 5153 76336
rect 5239 76313 5305 76336
rect 4919 76294 5305 76313
rect 20039 76399 20425 76418
rect 20039 76376 20105 76399
rect 20191 76376 20273 76399
rect 20359 76376 20425 76399
rect 20039 76336 20048 76376
rect 20088 76336 20105 76376
rect 20191 76336 20212 76376
rect 20252 76336 20273 76376
rect 20359 76336 20376 76376
rect 20416 76336 20425 76376
rect 20039 76313 20105 76336
rect 20191 76313 20273 76336
rect 20359 76313 20425 76336
rect 20039 76294 20425 76313
rect 13219 75916 13228 75956
rect 13268 75916 18892 75956
rect 18932 75916 18941 75956
rect 3679 75643 4065 75662
rect 3679 75620 3745 75643
rect 3831 75620 3913 75643
rect 3999 75620 4065 75643
rect 3679 75580 3688 75620
rect 3728 75580 3745 75620
rect 3831 75580 3852 75620
rect 3892 75580 3913 75620
rect 3999 75580 4016 75620
rect 4056 75580 4065 75620
rect 3679 75557 3745 75580
rect 3831 75557 3913 75580
rect 3999 75557 4065 75580
rect 3679 75538 4065 75557
rect 18799 75643 19185 75662
rect 18799 75620 18865 75643
rect 18951 75620 19033 75643
rect 19119 75620 19185 75643
rect 18799 75580 18808 75620
rect 18848 75580 18865 75620
rect 18951 75580 18972 75620
rect 19012 75580 19033 75620
rect 19119 75580 19136 75620
rect 19176 75580 19185 75620
rect 18799 75557 18865 75580
rect 18951 75557 19033 75580
rect 19119 75557 19185 75580
rect 18799 75538 19185 75557
rect 4919 74887 5305 74906
rect 4919 74864 4985 74887
rect 5071 74864 5153 74887
rect 5239 74864 5305 74887
rect 4919 74824 4928 74864
rect 4968 74824 4985 74864
rect 5071 74824 5092 74864
rect 5132 74824 5153 74864
rect 5239 74824 5256 74864
rect 5296 74824 5305 74864
rect 4919 74801 4985 74824
rect 5071 74801 5153 74824
rect 5239 74801 5305 74824
rect 4919 74782 5305 74801
rect 20039 74887 20425 74906
rect 20039 74864 20105 74887
rect 20191 74864 20273 74887
rect 20359 74864 20425 74887
rect 20039 74824 20048 74864
rect 20088 74824 20105 74864
rect 20191 74824 20212 74864
rect 20252 74824 20273 74864
rect 20359 74824 20376 74864
rect 20416 74824 20425 74864
rect 20039 74801 20105 74824
rect 20191 74801 20273 74824
rect 20359 74801 20425 74824
rect 20039 74782 20425 74801
rect 3679 74131 4065 74150
rect 3679 74108 3745 74131
rect 3831 74108 3913 74131
rect 3999 74108 4065 74131
rect 3679 74068 3688 74108
rect 3728 74068 3745 74108
rect 3831 74068 3852 74108
rect 3892 74068 3913 74108
rect 3999 74068 4016 74108
rect 4056 74068 4065 74108
rect 3679 74045 3745 74068
rect 3831 74045 3913 74068
rect 3999 74045 4065 74068
rect 3679 74026 4065 74045
rect 18799 74131 19185 74150
rect 18799 74108 18865 74131
rect 18951 74108 19033 74131
rect 19119 74108 19185 74131
rect 18799 74068 18808 74108
rect 18848 74068 18865 74108
rect 18951 74068 18972 74108
rect 19012 74068 19033 74108
rect 19119 74068 19136 74108
rect 19176 74068 19185 74108
rect 18799 74045 18865 74068
rect 18951 74045 19033 74068
rect 19119 74045 19185 74068
rect 18799 74026 19185 74045
rect 4919 73375 5305 73394
rect 4919 73352 4985 73375
rect 5071 73352 5153 73375
rect 5239 73352 5305 73375
rect 4919 73312 4928 73352
rect 4968 73312 4985 73352
rect 5071 73312 5092 73352
rect 5132 73312 5153 73352
rect 5239 73312 5256 73352
rect 5296 73312 5305 73352
rect 4919 73289 4985 73312
rect 5071 73289 5153 73312
rect 5239 73289 5305 73312
rect 4919 73270 5305 73289
rect 20039 73375 20425 73394
rect 20039 73352 20105 73375
rect 20191 73352 20273 73375
rect 20359 73352 20425 73375
rect 20039 73312 20048 73352
rect 20088 73312 20105 73352
rect 20191 73312 20212 73352
rect 20252 73312 20273 73352
rect 20359 73312 20376 73352
rect 20416 73312 20425 73352
rect 20039 73289 20105 73312
rect 20191 73289 20273 73312
rect 20359 73289 20425 73312
rect 20039 73270 20425 73289
rect 3679 72619 4065 72638
rect 3679 72596 3745 72619
rect 3831 72596 3913 72619
rect 3999 72596 4065 72619
rect 3679 72556 3688 72596
rect 3728 72556 3745 72596
rect 3831 72556 3852 72596
rect 3892 72556 3913 72596
rect 3999 72556 4016 72596
rect 4056 72556 4065 72596
rect 3679 72533 3745 72556
rect 3831 72533 3913 72556
rect 3999 72533 4065 72556
rect 3679 72514 4065 72533
rect 18799 72619 19185 72638
rect 18799 72596 18865 72619
rect 18951 72596 19033 72619
rect 19119 72596 19185 72619
rect 18799 72556 18808 72596
rect 18848 72556 18865 72596
rect 18951 72556 18972 72596
rect 19012 72556 19033 72596
rect 19119 72556 19136 72596
rect 19176 72556 19185 72596
rect 18799 72533 18865 72556
rect 18951 72533 19033 72556
rect 19119 72533 19185 72556
rect 18799 72514 19185 72533
rect 11203 72220 11212 72260
rect 11252 72220 19756 72260
rect 19796 72220 19805 72260
rect 4919 71863 5305 71882
rect 4919 71840 4985 71863
rect 5071 71840 5153 71863
rect 5239 71840 5305 71863
rect 4919 71800 4928 71840
rect 4968 71800 4985 71840
rect 5071 71800 5092 71840
rect 5132 71800 5153 71840
rect 5239 71800 5256 71840
rect 5296 71800 5305 71840
rect 4919 71777 4985 71800
rect 5071 71777 5153 71800
rect 5239 71777 5305 71800
rect 4919 71758 5305 71777
rect 20039 71863 20425 71882
rect 20039 71840 20105 71863
rect 20191 71840 20273 71863
rect 20359 71840 20425 71863
rect 20039 71800 20048 71840
rect 20088 71800 20105 71840
rect 20191 71800 20212 71840
rect 20252 71800 20273 71840
rect 20359 71800 20376 71840
rect 20416 71800 20425 71840
rect 20039 71777 20105 71800
rect 20191 71777 20273 71800
rect 20359 71777 20425 71800
rect 20039 71758 20425 71777
rect 3679 71107 4065 71126
rect 3679 71084 3745 71107
rect 3831 71084 3913 71107
rect 3999 71084 4065 71107
rect 3679 71044 3688 71084
rect 3728 71044 3745 71084
rect 3831 71044 3852 71084
rect 3892 71044 3913 71084
rect 3999 71044 4016 71084
rect 4056 71044 4065 71084
rect 3679 71021 3745 71044
rect 3831 71021 3913 71044
rect 3999 71021 4065 71044
rect 3679 71002 4065 71021
rect 18799 71107 19185 71126
rect 18799 71084 18865 71107
rect 18951 71084 19033 71107
rect 19119 71084 19185 71107
rect 18799 71044 18808 71084
rect 18848 71044 18865 71084
rect 18951 71044 18972 71084
rect 19012 71044 19033 71084
rect 19119 71044 19136 71084
rect 19176 71044 19185 71084
rect 18799 71021 18865 71044
rect 18951 71021 19033 71044
rect 19119 71021 19185 71044
rect 18799 71002 19185 71021
rect 4919 70351 5305 70370
rect 4919 70328 4985 70351
rect 5071 70328 5153 70351
rect 5239 70328 5305 70351
rect 4919 70288 4928 70328
rect 4968 70288 4985 70328
rect 5071 70288 5092 70328
rect 5132 70288 5153 70328
rect 5239 70288 5256 70328
rect 5296 70288 5305 70328
rect 4919 70265 4985 70288
rect 5071 70265 5153 70288
rect 5239 70265 5305 70288
rect 4919 70246 5305 70265
rect 20039 70351 20425 70370
rect 20039 70328 20105 70351
rect 20191 70328 20273 70351
rect 20359 70328 20425 70351
rect 20039 70288 20048 70328
rect 20088 70288 20105 70328
rect 20191 70288 20212 70328
rect 20252 70288 20273 70328
rect 20359 70288 20376 70328
rect 20416 70288 20425 70328
rect 20039 70265 20105 70288
rect 20191 70265 20273 70288
rect 20359 70265 20425 70288
rect 20039 70246 20425 70265
rect 3679 69595 4065 69614
rect 3679 69572 3745 69595
rect 3831 69572 3913 69595
rect 3999 69572 4065 69595
rect 3679 69532 3688 69572
rect 3728 69532 3745 69572
rect 3831 69532 3852 69572
rect 3892 69532 3913 69572
rect 3999 69532 4016 69572
rect 4056 69532 4065 69572
rect 3679 69509 3745 69532
rect 3831 69509 3913 69532
rect 3999 69509 4065 69532
rect 3679 69490 4065 69509
rect 18799 69595 19185 69614
rect 18799 69572 18865 69595
rect 18951 69572 19033 69595
rect 19119 69572 19185 69595
rect 18799 69532 18808 69572
rect 18848 69532 18865 69572
rect 18951 69532 18972 69572
rect 19012 69532 19033 69572
rect 19119 69532 19136 69572
rect 19176 69532 19185 69572
rect 18799 69509 18865 69532
rect 18951 69509 19033 69532
rect 19119 69509 19185 69532
rect 18799 69490 19185 69509
rect 4919 68839 5305 68858
rect 4919 68816 4985 68839
rect 5071 68816 5153 68839
rect 5239 68816 5305 68839
rect 4919 68776 4928 68816
rect 4968 68776 4985 68816
rect 5071 68776 5092 68816
rect 5132 68776 5153 68816
rect 5239 68776 5256 68816
rect 5296 68776 5305 68816
rect 4919 68753 4985 68776
rect 5071 68753 5153 68776
rect 5239 68753 5305 68776
rect 4919 68734 5305 68753
rect 20039 68839 20425 68858
rect 20039 68816 20105 68839
rect 20191 68816 20273 68839
rect 20359 68816 20425 68839
rect 20039 68776 20048 68816
rect 20088 68776 20105 68816
rect 20191 68776 20212 68816
rect 20252 68776 20273 68816
rect 20359 68776 20376 68816
rect 20416 68776 20425 68816
rect 20039 68753 20105 68776
rect 20191 68753 20273 68776
rect 20359 68753 20425 68776
rect 20039 68734 20425 68753
rect 3679 68083 4065 68102
rect 3679 68060 3745 68083
rect 3831 68060 3913 68083
rect 3999 68060 4065 68083
rect 18799 68083 19185 68102
rect 18799 68060 18865 68083
rect 18951 68060 19033 68083
rect 19119 68060 19185 68083
rect 3679 68020 3688 68060
rect 3728 68020 3745 68060
rect 3831 68020 3852 68060
rect 3892 68020 3913 68060
rect 3999 68020 4016 68060
rect 4056 68020 4065 68060
rect 6787 68020 6796 68060
rect 6836 68020 11308 68060
rect 11348 68020 11357 68060
rect 18799 68020 18808 68060
rect 18848 68020 18865 68060
rect 18951 68020 18972 68060
rect 19012 68020 19033 68060
rect 19119 68020 19136 68060
rect 19176 68020 19185 68060
rect 3679 67997 3745 68020
rect 3831 67997 3913 68020
rect 3999 67997 4065 68020
rect 3679 67978 4065 67997
rect 18799 67997 18865 68020
rect 18951 67997 19033 68020
rect 19119 67997 19185 68020
rect 18799 67978 19185 67997
rect 4919 67327 5305 67346
rect 4919 67304 4985 67327
rect 5071 67304 5153 67327
rect 5239 67304 5305 67327
rect 4919 67264 4928 67304
rect 4968 67264 4985 67304
rect 5071 67264 5092 67304
rect 5132 67264 5153 67304
rect 5239 67264 5256 67304
rect 5296 67264 5305 67304
rect 4919 67241 4985 67264
rect 5071 67241 5153 67264
rect 5239 67241 5305 67264
rect 4919 67222 5305 67241
rect 20039 67327 20425 67346
rect 20039 67304 20105 67327
rect 20191 67304 20273 67327
rect 20359 67304 20425 67327
rect 20039 67264 20048 67304
rect 20088 67264 20105 67304
rect 20191 67264 20212 67304
rect 20252 67264 20273 67304
rect 20359 67264 20376 67304
rect 20416 67264 20425 67304
rect 20039 67241 20105 67264
rect 20191 67241 20273 67264
rect 20359 67241 20425 67264
rect 20039 67222 20425 67241
rect 3679 66571 4065 66590
rect 3679 66548 3745 66571
rect 3831 66548 3913 66571
rect 3999 66548 4065 66571
rect 3679 66508 3688 66548
rect 3728 66508 3745 66548
rect 3831 66508 3852 66548
rect 3892 66508 3913 66548
rect 3999 66508 4016 66548
rect 4056 66508 4065 66548
rect 3679 66485 3745 66508
rect 3831 66485 3913 66508
rect 3999 66485 4065 66508
rect 3679 66466 4065 66485
rect 18799 66571 19185 66590
rect 18799 66548 18865 66571
rect 18951 66548 19033 66571
rect 19119 66548 19185 66571
rect 18799 66508 18808 66548
rect 18848 66508 18865 66548
rect 18951 66508 18972 66548
rect 19012 66508 19033 66548
rect 19119 66508 19136 66548
rect 19176 66508 19185 66548
rect 18799 66485 18865 66508
rect 18951 66485 19033 66508
rect 19119 66485 19185 66508
rect 18799 66466 19185 66485
rect 4919 65815 5305 65834
rect 4919 65792 4985 65815
rect 5071 65792 5153 65815
rect 5239 65792 5305 65815
rect 4919 65752 4928 65792
rect 4968 65752 4985 65792
rect 5071 65752 5092 65792
rect 5132 65752 5153 65792
rect 5239 65752 5256 65792
rect 5296 65752 5305 65792
rect 4919 65729 4985 65752
rect 5071 65729 5153 65752
rect 5239 65729 5305 65752
rect 4919 65710 5305 65729
rect 20039 65815 20425 65834
rect 20039 65792 20105 65815
rect 20191 65792 20273 65815
rect 20359 65792 20425 65815
rect 20039 65752 20048 65792
rect 20088 65752 20105 65792
rect 20191 65752 20212 65792
rect 20252 65752 20273 65792
rect 20359 65752 20376 65792
rect 20416 65752 20425 65792
rect 20039 65729 20105 65752
rect 20191 65729 20273 65752
rect 20359 65729 20425 65752
rect 20039 65710 20425 65729
rect 3679 65059 4065 65078
rect 3679 65036 3745 65059
rect 3831 65036 3913 65059
rect 3999 65036 4065 65059
rect 3679 64996 3688 65036
rect 3728 64996 3745 65036
rect 3831 64996 3852 65036
rect 3892 64996 3913 65036
rect 3999 64996 4016 65036
rect 4056 64996 4065 65036
rect 3679 64973 3745 64996
rect 3831 64973 3913 64996
rect 3999 64973 4065 64996
rect 3679 64954 4065 64973
rect 18799 65059 19185 65078
rect 18799 65036 18865 65059
rect 18951 65036 19033 65059
rect 19119 65036 19185 65059
rect 18799 64996 18808 65036
rect 18848 64996 18865 65036
rect 18951 64996 18972 65036
rect 19012 64996 19033 65036
rect 19119 64996 19136 65036
rect 19176 64996 19185 65036
rect 18799 64973 18865 64996
rect 18951 64973 19033 64996
rect 19119 64973 19185 64996
rect 18799 64954 19185 64973
rect 4919 64303 5305 64322
rect 4919 64280 4985 64303
rect 5071 64280 5153 64303
rect 5239 64280 5305 64303
rect 4919 64240 4928 64280
rect 4968 64240 4985 64280
rect 5071 64240 5092 64280
rect 5132 64240 5153 64280
rect 5239 64240 5256 64280
rect 5296 64240 5305 64280
rect 4919 64217 4985 64240
rect 5071 64217 5153 64240
rect 5239 64217 5305 64240
rect 4919 64198 5305 64217
rect 20039 64303 20425 64322
rect 20039 64280 20105 64303
rect 20191 64280 20273 64303
rect 20359 64280 20425 64303
rect 20039 64240 20048 64280
rect 20088 64240 20105 64280
rect 20191 64240 20212 64280
rect 20252 64240 20273 64280
rect 20359 64240 20376 64280
rect 20416 64240 20425 64280
rect 20039 64217 20105 64240
rect 20191 64217 20273 64240
rect 20359 64217 20425 64240
rect 20039 64198 20425 64217
rect 3679 63547 4065 63566
rect 3679 63524 3745 63547
rect 3831 63524 3913 63547
rect 3999 63524 4065 63547
rect 3679 63484 3688 63524
rect 3728 63484 3745 63524
rect 3831 63484 3852 63524
rect 3892 63484 3913 63524
rect 3999 63484 4016 63524
rect 4056 63484 4065 63524
rect 3679 63461 3745 63484
rect 3831 63461 3913 63484
rect 3999 63461 4065 63484
rect 3679 63442 4065 63461
rect 18799 63547 19185 63566
rect 18799 63524 18865 63547
rect 18951 63524 19033 63547
rect 19119 63524 19185 63547
rect 18799 63484 18808 63524
rect 18848 63484 18865 63524
rect 18951 63484 18972 63524
rect 19012 63484 19033 63524
rect 19119 63484 19136 63524
rect 19176 63484 19185 63524
rect 18799 63461 18865 63484
rect 18951 63461 19033 63484
rect 19119 63461 19185 63484
rect 18799 63442 19185 63461
rect 4919 62791 5305 62810
rect 4919 62768 4985 62791
rect 5071 62768 5153 62791
rect 5239 62768 5305 62791
rect 4919 62728 4928 62768
rect 4968 62728 4985 62768
rect 5071 62728 5092 62768
rect 5132 62728 5153 62768
rect 5239 62728 5256 62768
rect 5296 62728 5305 62768
rect 4919 62705 4985 62728
rect 5071 62705 5153 62728
rect 5239 62705 5305 62728
rect 4919 62686 5305 62705
rect 20039 62791 20425 62810
rect 20039 62768 20105 62791
rect 20191 62768 20273 62791
rect 20359 62768 20425 62791
rect 20039 62728 20048 62768
rect 20088 62728 20105 62768
rect 20191 62728 20212 62768
rect 20252 62728 20273 62768
rect 20359 62728 20376 62768
rect 20416 62728 20425 62768
rect 20039 62705 20105 62728
rect 20191 62705 20273 62728
rect 20359 62705 20425 62728
rect 20039 62686 20425 62705
rect 3679 62035 4065 62054
rect 3679 62012 3745 62035
rect 3831 62012 3913 62035
rect 3999 62012 4065 62035
rect 3679 61972 3688 62012
rect 3728 61972 3745 62012
rect 3831 61972 3852 62012
rect 3892 61972 3913 62012
rect 3999 61972 4016 62012
rect 4056 61972 4065 62012
rect 3679 61949 3745 61972
rect 3831 61949 3913 61972
rect 3999 61949 4065 61972
rect 3679 61930 4065 61949
rect 18799 62035 19185 62054
rect 18799 62012 18865 62035
rect 18951 62012 19033 62035
rect 19119 62012 19185 62035
rect 18799 61972 18808 62012
rect 18848 61972 18865 62012
rect 18951 61972 18972 62012
rect 19012 61972 19033 62012
rect 19119 61972 19136 62012
rect 19176 61972 19185 62012
rect 18799 61949 18865 61972
rect 18951 61949 19033 61972
rect 19119 61949 19185 61972
rect 18799 61930 19185 61949
rect 4919 61279 5305 61298
rect 4919 61256 4985 61279
rect 5071 61256 5153 61279
rect 5239 61256 5305 61279
rect 4919 61216 4928 61256
rect 4968 61216 4985 61256
rect 5071 61216 5092 61256
rect 5132 61216 5153 61256
rect 5239 61216 5256 61256
rect 5296 61216 5305 61256
rect 4919 61193 4985 61216
rect 5071 61193 5153 61216
rect 5239 61193 5305 61216
rect 4919 61174 5305 61193
rect 20039 61279 20425 61298
rect 20039 61256 20105 61279
rect 20191 61256 20273 61279
rect 20359 61256 20425 61279
rect 20039 61216 20048 61256
rect 20088 61216 20105 61256
rect 20191 61216 20212 61256
rect 20252 61216 20273 61256
rect 20359 61216 20376 61256
rect 20416 61216 20425 61256
rect 20039 61193 20105 61216
rect 20191 61193 20273 61216
rect 20359 61193 20425 61216
rect 20039 61174 20425 61193
rect 3679 60523 4065 60542
rect 3679 60500 3745 60523
rect 3831 60500 3913 60523
rect 3999 60500 4065 60523
rect 3679 60460 3688 60500
rect 3728 60460 3745 60500
rect 3831 60460 3852 60500
rect 3892 60460 3913 60500
rect 3999 60460 4016 60500
rect 4056 60460 4065 60500
rect 3679 60437 3745 60460
rect 3831 60437 3913 60460
rect 3999 60437 4065 60460
rect 3679 60418 4065 60437
rect 18799 60523 19185 60542
rect 18799 60500 18865 60523
rect 18951 60500 19033 60523
rect 19119 60500 19185 60523
rect 18799 60460 18808 60500
rect 18848 60460 18865 60500
rect 18951 60460 18972 60500
rect 19012 60460 19033 60500
rect 19119 60460 19136 60500
rect 19176 60460 19185 60500
rect 18799 60437 18865 60460
rect 18951 60437 19033 60460
rect 19119 60437 19185 60460
rect 18799 60418 19185 60437
rect 1027 59872 1036 59912
rect 1076 59872 12652 59912
rect 12692 59872 12701 59912
rect 4919 59767 5305 59786
rect 4919 59744 4985 59767
rect 5071 59744 5153 59767
rect 5239 59744 5305 59767
rect 4919 59704 4928 59744
rect 4968 59704 4985 59744
rect 5071 59704 5092 59744
rect 5132 59704 5153 59744
rect 5239 59704 5256 59744
rect 5296 59704 5305 59744
rect 4919 59681 4985 59704
rect 5071 59681 5153 59704
rect 5239 59681 5305 59704
rect 4919 59662 5305 59681
rect 20039 59767 20425 59786
rect 20039 59744 20105 59767
rect 20191 59744 20273 59767
rect 20359 59744 20425 59767
rect 20039 59704 20048 59744
rect 20088 59704 20105 59744
rect 20191 59704 20212 59744
rect 20252 59704 20273 59744
rect 20359 59704 20376 59744
rect 20416 59704 20425 59744
rect 20039 59681 20105 59704
rect 20191 59681 20273 59704
rect 20359 59681 20425 59704
rect 20039 59662 20425 59681
rect 3679 59011 4065 59030
rect 3679 58988 3745 59011
rect 3831 58988 3913 59011
rect 3999 58988 4065 59011
rect 3679 58948 3688 58988
rect 3728 58948 3745 58988
rect 3831 58948 3852 58988
rect 3892 58948 3913 58988
rect 3999 58948 4016 58988
rect 4056 58948 4065 58988
rect 3679 58925 3745 58948
rect 3831 58925 3913 58948
rect 3999 58925 4065 58948
rect 3679 58906 4065 58925
rect 18799 59011 19185 59030
rect 18799 58988 18865 59011
rect 18951 58988 19033 59011
rect 19119 58988 19185 59011
rect 18799 58948 18808 58988
rect 18848 58948 18865 58988
rect 18951 58948 18972 58988
rect 19012 58948 19033 58988
rect 19119 58948 19136 58988
rect 19176 58948 19185 58988
rect 18799 58925 18865 58948
rect 18951 58925 19033 58948
rect 19119 58925 19185 58948
rect 18799 58906 19185 58925
rect 4919 58255 5305 58274
rect 4919 58232 4985 58255
rect 5071 58232 5153 58255
rect 5239 58232 5305 58255
rect 4919 58192 4928 58232
rect 4968 58192 4985 58232
rect 5071 58192 5092 58232
rect 5132 58192 5153 58232
rect 5239 58192 5256 58232
rect 5296 58192 5305 58232
rect 4919 58169 4985 58192
rect 5071 58169 5153 58192
rect 5239 58169 5305 58192
rect 4919 58150 5305 58169
rect 20039 58255 20425 58274
rect 20039 58232 20105 58255
rect 20191 58232 20273 58255
rect 20359 58232 20425 58255
rect 20039 58192 20048 58232
rect 20088 58192 20105 58232
rect 20191 58192 20212 58232
rect 20252 58192 20273 58232
rect 20359 58192 20376 58232
rect 20416 58192 20425 58232
rect 20039 58169 20105 58192
rect 20191 58169 20273 58192
rect 20359 58169 20425 58192
rect 20039 58150 20425 58169
rect 7939 57940 7948 57980
rect 7988 57940 10060 57980
rect 10100 57940 10109 57980
rect 3427 57856 3436 57896
rect 3476 57856 10732 57896
rect 10772 57856 10781 57896
rect 3679 57499 4065 57518
rect 3679 57476 3745 57499
rect 3831 57476 3913 57499
rect 3999 57476 4065 57499
rect 3679 57436 3688 57476
rect 3728 57436 3745 57476
rect 3831 57436 3852 57476
rect 3892 57436 3913 57476
rect 3999 57436 4016 57476
rect 4056 57436 4065 57476
rect 3679 57413 3745 57436
rect 3831 57413 3913 57436
rect 3999 57413 4065 57436
rect 3679 57394 4065 57413
rect 18799 57499 19185 57518
rect 18799 57476 18865 57499
rect 18951 57476 19033 57499
rect 19119 57476 19185 57499
rect 18799 57436 18808 57476
rect 18848 57436 18865 57476
rect 18951 57436 18972 57476
rect 19012 57436 19033 57476
rect 19119 57436 19136 57476
rect 19176 57436 19185 57476
rect 18799 57413 18865 57436
rect 18951 57413 19033 57436
rect 19119 57413 19185 57436
rect 18799 57394 19185 57413
rect 3523 56848 3532 56888
rect 3572 56848 11500 56888
rect 11540 56848 11549 56888
rect 4919 56743 5305 56762
rect 4919 56720 4985 56743
rect 5071 56720 5153 56743
rect 5239 56720 5305 56743
rect 4919 56680 4928 56720
rect 4968 56680 4985 56720
rect 5071 56680 5092 56720
rect 5132 56680 5153 56720
rect 5239 56680 5256 56720
rect 5296 56680 5305 56720
rect 4919 56657 4985 56680
rect 5071 56657 5153 56680
rect 5239 56657 5305 56680
rect 4919 56638 5305 56657
rect 20039 56743 20425 56762
rect 20039 56720 20105 56743
rect 20191 56720 20273 56743
rect 20359 56720 20425 56743
rect 20039 56680 20048 56720
rect 20088 56680 20105 56720
rect 20191 56680 20212 56720
rect 20252 56680 20273 56720
rect 20359 56680 20376 56720
rect 20416 56680 20425 56720
rect 20039 56657 20105 56680
rect 20191 56657 20273 56680
rect 20359 56657 20425 56680
rect 20039 56638 20425 56657
rect 3679 55987 4065 56006
rect 3679 55964 3745 55987
rect 3831 55964 3913 55987
rect 3999 55964 4065 55987
rect 3679 55924 3688 55964
rect 3728 55924 3745 55964
rect 3831 55924 3852 55964
rect 3892 55924 3913 55964
rect 3999 55924 4016 55964
rect 4056 55924 4065 55964
rect 3679 55901 3745 55924
rect 3831 55901 3913 55924
rect 3999 55901 4065 55924
rect 3679 55882 4065 55901
rect 18799 55987 19185 56006
rect 18799 55964 18865 55987
rect 18951 55964 19033 55987
rect 19119 55964 19185 55987
rect 18799 55924 18808 55964
rect 18848 55924 18865 55964
rect 18951 55924 18972 55964
rect 19012 55924 19033 55964
rect 19119 55924 19136 55964
rect 19176 55924 19185 55964
rect 18799 55901 18865 55924
rect 18951 55901 19033 55924
rect 19119 55901 19185 55924
rect 18799 55882 19185 55901
rect 4919 55231 5305 55250
rect 4919 55208 4985 55231
rect 5071 55208 5153 55231
rect 5239 55208 5305 55231
rect 4919 55168 4928 55208
rect 4968 55168 4985 55208
rect 5071 55168 5092 55208
rect 5132 55168 5153 55208
rect 5239 55168 5256 55208
rect 5296 55168 5305 55208
rect 4919 55145 4985 55168
rect 5071 55145 5153 55168
rect 5239 55145 5305 55168
rect 4919 55126 5305 55145
rect 20039 55231 20425 55250
rect 20039 55208 20105 55231
rect 20191 55208 20273 55231
rect 20359 55208 20425 55231
rect 20039 55168 20048 55208
rect 20088 55168 20105 55208
rect 20191 55168 20212 55208
rect 20252 55168 20273 55208
rect 20359 55168 20376 55208
rect 20416 55168 20425 55208
rect 20039 55145 20105 55168
rect 20191 55145 20273 55168
rect 20359 55145 20425 55168
rect 20039 55126 20425 55145
rect 3679 54475 4065 54494
rect 3679 54452 3745 54475
rect 3831 54452 3913 54475
rect 3999 54452 4065 54475
rect 3679 54412 3688 54452
rect 3728 54412 3745 54452
rect 3831 54412 3852 54452
rect 3892 54412 3913 54452
rect 3999 54412 4016 54452
rect 4056 54412 4065 54452
rect 3679 54389 3745 54412
rect 3831 54389 3913 54412
rect 3999 54389 4065 54412
rect 3679 54370 4065 54389
rect 18799 54475 19185 54494
rect 18799 54452 18865 54475
rect 18951 54452 19033 54475
rect 19119 54452 19185 54475
rect 18799 54412 18808 54452
rect 18848 54412 18865 54452
rect 18951 54412 18972 54452
rect 19012 54412 19033 54452
rect 19119 54412 19136 54452
rect 19176 54412 19185 54452
rect 18799 54389 18865 54412
rect 18951 54389 19033 54412
rect 19119 54389 19185 54412
rect 18799 54370 19185 54389
rect 4919 53719 5305 53738
rect 4919 53696 4985 53719
rect 5071 53696 5153 53719
rect 5239 53696 5305 53719
rect 4919 53656 4928 53696
rect 4968 53656 4985 53696
rect 5071 53656 5092 53696
rect 5132 53656 5153 53696
rect 5239 53656 5256 53696
rect 5296 53656 5305 53696
rect 4919 53633 4985 53656
rect 5071 53633 5153 53656
rect 5239 53633 5305 53656
rect 4919 53614 5305 53633
rect 20039 53719 20425 53738
rect 20039 53696 20105 53719
rect 20191 53696 20273 53719
rect 20359 53696 20425 53719
rect 20039 53656 20048 53696
rect 20088 53656 20105 53696
rect 20191 53656 20212 53696
rect 20252 53656 20273 53696
rect 20359 53656 20376 53696
rect 20416 53656 20425 53696
rect 20039 53633 20105 53656
rect 20191 53633 20273 53656
rect 20359 53633 20425 53656
rect 20039 53614 20425 53633
rect 7267 53236 7276 53276
rect 7316 53236 11360 53276
rect 16963 53236 16972 53276
rect 17012 53236 18700 53276
rect 18740 53236 18749 53276
rect 11320 53192 11360 53236
rect 11320 53152 20140 53192
rect 20180 53152 20189 53192
rect 3679 52963 4065 52982
rect 3679 52940 3745 52963
rect 3831 52940 3913 52963
rect 3999 52940 4065 52963
rect 3679 52900 3688 52940
rect 3728 52900 3745 52940
rect 3831 52900 3852 52940
rect 3892 52900 3913 52940
rect 3999 52900 4016 52940
rect 4056 52900 4065 52940
rect 3679 52877 3745 52900
rect 3831 52877 3913 52900
rect 3999 52877 4065 52900
rect 3679 52858 4065 52877
rect 18799 52963 19185 52982
rect 18799 52940 18865 52963
rect 18951 52940 19033 52963
rect 19119 52940 19185 52963
rect 18799 52900 18808 52940
rect 18848 52900 18865 52940
rect 18951 52900 18972 52940
rect 19012 52900 19033 52940
rect 19119 52900 19136 52940
rect 19176 52900 19185 52940
rect 18799 52877 18865 52900
rect 18951 52877 19033 52900
rect 19119 52877 19185 52900
rect 18799 52858 19185 52877
rect 4919 52207 5305 52226
rect 4919 52184 4985 52207
rect 5071 52184 5153 52207
rect 5239 52184 5305 52207
rect 4919 52144 4928 52184
rect 4968 52144 4985 52184
rect 5071 52144 5092 52184
rect 5132 52144 5153 52184
rect 5239 52144 5256 52184
rect 5296 52144 5305 52184
rect 4919 52121 4985 52144
rect 5071 52121 5153 52144
rect 5239 52121 5305 52144
rect 4919 52102 5305 52121
rect 20039 52207 20425 52226
rect 20039 52184 20105 52207
rect 20191 52184 20273 52207
rect 20359 52184 20425 52207
rect 20039 52144 20048 52184
rect 20088 52144 20105 52184
rect 20191 52144 20212 52184
rect 20252 52144 20273 52184
rect 20359 52144 20376 52184
rect 20416 52144 20425 52184
rect 20039 52121 20105 52144
rect 20191 52121 20273 52144
rect 20359 52121 20425 52144
rect 20039 52102 20425 52121
rect 2851 51976 2860 52016
rect 2900 51976 3148 52016
rect 3188 51976 3197 52016
rect 4291 51808 4300 51848
rect 4340 51808 17644 51848
rect 17684 51808 17693 51848
rect 3679 51451 4065 51470
rect 3679 51428 3745 51451
rect 3831 51428 3913 51451
rect 3999 51428 4065 51451
rect 3679 51388 3688 51428
rect 3728 51388 3745 51428
rect 3831 51388 3852 51428
rect 3892 51388 3913 51428
rect 3999 51388 4016 51428
rect 4056 51388 4065 51428
rect 3679 51365 3745 51388
rect 3831 51365 3913 51388
rect 3999 51365 4065 51388
rect 3679 51346 4065 51365
rect 18799 51451 19185 51470
rect 18799 51428 18865 51451
rect 18951 51428 19033 51451
rect 19119 51428 19185 51451
rect 18799 51388 18808 51428
rect 18848 51388 18865 51428
rect 18951 51388 18972 51428
rect 19012 51388 19033 51428
rect 19119 51388 19136 51428
rect 19176 51388 19185 51428
rect 18799 51365 18865 51388
rect 18951 51365 19033 51388
rect 19119 51365 19185 51388
rect 18799 51346 19185 51365
rect 4919 50695 5305 50714
rect 4919 50672 4985 50695
rect 5071 50672 5153 50695
rect 5239 50672 5305 50695
rect 4919 50632 4928 50672
rect 4968 50632 4985 50672
rect 5071 50632 5092 50672
rect 5132 50632 5153 50672
rect 5239 50632 5256 50672
rect 5296 50632 5305 50672
rect 4919 50609 4985 50632
rect 5071 50609 5153 50632
rect 5239 50609 5305 50632
rect 4919 50590 5305 50609
rect 20039 50695 20425 50714
rect 20039 50672 20105 50695
rect 20191 50672 20273 50695
rect 20359 50672 20425 50695
rect 20039 50632 20048 50672
rect 20088 50632 20105 50672
rect 20191 50632 20212 50672
rect 20252 50632 20273 50672
rect 20359 50632 20376 50672
rect 20416 50632 20425 50672
rect 20039 50609 20105 50632
rect 20191 50609 20273 50632
rect 20359 50609 20425 50632
rect 20039 50590 20425 50609
rect 3679 49939 4065 49958
rect 3679 49916 3745 49939
rect 3831 49916 3913 49939
rect 3999 49916 4065 49939
rect 3679 49876 3688 49916
rect 3728 49876 3745 49916
rect 3831 49876 3852 49916
rect 3892 49876 3913 49916
rect 3999 49876 4016 49916
rect 4056 49876 4065 49916
rect 3679 49853 3745 49876
rect 3831 49853 3913 49876
rect 3999 49853 4065 49876
rect 3679 49834 4065 49853
rect 18799 49939 19185 49958
rect 18799 49916 18865 49939
rect 18951 49916 19033 49939
rect 19119 49916 19185 49939
rect 18799 49876 18808 49916
rect 18848 49876 18865 49916
rect 18951 49876 18972 49916
rect 19012 49876 19033 49916
rect 19119 49876 19136 49916
rect 19176 49876 19185 49916
rect 18799 49853 18865 49876
rect 18951 49853 19033 49876
rect 19119 49853 19185 49876
rect 18799 49834 19185 49853
rect 4919 49183 5305 49202
rect 4919 49160 4985 49183
rect 5071 49160 5153 49183
rect 5239 49160 5305 49183
rect 4919 49120 4928 49160
rect 4968 49120 4985 49160
rect 5071 49120 5092 49160
rect 5132 49120 5153 49160
rect 5239 49120 5256 49160
rect 5296 49120 5305 49160
rect 4919 49097 4985 49120
rect 5071 49097 5153 49120
rect 5239 49097 5305 49120
rect 4919 49078 5305 49097
rect 20039 49183 20425 49202
rect 20039 49160 20105 49183
rect 20191 49160 20273 49183
rect 20359 49160 20425 49183
rect 20039 49120 20048 49160
rect 20088 49120 20105 49160
rect 20191 49120 20212 49160
rect 20252 49120 20273 49160
rect 20359 49120 20376 49160
rect 20416 49120 20425 49160
rect 20039 49097 20105 49120
rect 20191 49097 20273 49120
rect 20359 49097 20425 49120
rect 20039 49078 20425 49097
rect 3679 48427 4065 48446
rect 3679 48404 3745 48427
rect 3831 48404 3913 48427
rect 3999 48404 4065 48427
rect 3679 48364 3688 48404
rect 3728 48364 3745 48404
rect 3831 48364 3852 48404
rect 3892 48364 3913 48404
rect 3999 48364 4016 48404
rect 4056 48364 4065 48404
rect 3679 48341 3745 48364
rect 3831 48341 3913 48364
rect 3999 48341 4065 48364
rect 3679 48322 4065 48341
rect 18799 48427 19185 48446
rect 18799 48404 18865 48427
rect 18951 48404 19033 48427
rect 19119 48404 19185 48427
rect 18799 48364 18808 48404
rect 18848 48364 18865 48404
rect 18951 48364 18972 48404
rect 19012 48364 19033 48404
rect 19119 48364 19136 48404
rect 19176 48364 19185 48404
rect 18799 48341 18865 48364
rect 18951 48341 19033 48364
rect 19119 48341 19185 48364
rect 18799 48322 19185 48341
rect 2090 47923 2214 47942
rect 2090 47837 2109 47923
rect 2195 47900 2214 47923
rect 2195 47860 14284 47900
rect 14324 47860 14333 47900
rect 2195 47837 2214 47860
rect 2090 47818 2214 47837
rect 4919 47671 5305 47690
rect 4919 47648 4985 47671
rect 5071 47648 5153 47671
rect 5239 47648 5305 47671
rect 4919 47608 4928 47648
rect 4968 47608 4985 47648
rect 5071 47608 5092 47648
rect 5132 47608 5153 47648
rect 5239 47608 5256 47648
rect 5296 47608 5305 47648
rect 4919 47585 4985 47608
rect 5071 47585 5153 47608
rect 5239 47585 5305 47608
rect 4919 47566 5305 47585
rect 20039 47671 20425 47690
rect 20039 47648 20105 47671
rect 20191 47648 20273 47671
rect 20359 47648 20425 47671
rect 20039 47608 20048 47648
rect 20088 47608 20105 47648
rect 20191 47608 20212 47648
rect 20252 47608 20273 47648
rect 20359 47608 20376 47648
rect 20416 47608 20425 47648
rect 20039 47585 20105 47608
rect 20191 47585 20273 47608
rect 20359 47585 20425 47608
rect 20039 47566 20425 47585
rect 3679 46915 4065 46934
rect 3679 46892 3745 46915
rect 3831 46892 3913 46915
rect 3999 46892 4065 46915
rect 3679 46852 3688 46892
rect 3728 46852 3745 46892
rect 3831 46852 3852 46892
rect 3892 46852 3913 46892
rect 3999 46852 4016 46892
rect 4056 46852 4065 46892
rect 3679 46829 3745 46852
rect 3831 46829 3913 46852
rect 3999 46829 4065 46852
rect 3679 46810 4065 46829
rect 18799 46915 19185 46934
rect 18799 46892 18865 46915
rect 18951 46892 19033 46915
rect 19119 46892 19185 46915
rect 18799 46852 18808 46892
rect 18848 46852 18865 46892
rect 18951 46852 18972 46892
rect 19012 46852 19033 46892
rect 19119 46852 19136 46892
rect 19176 46852 19185 46892
rect 18799 46829 18865 46852
rect 18951 46829 19033 46852
rect 19119 46829 19185 46852
rect 18799 46810 19185 46829
rect 4919 46159 5305 46178
rect 4919 46136 4985 46159
rect 5071 46136 5153 46159
rect 5239 46136 5305 46159
rect 4919 46096 4928 46136
rect 4968 46096 4985 46136
rect 5071 46096 5092 46136
rect 5132 46096 5153 46136
rect 5239 46096 5256 46136
rect 5296 46096 5305 46136
rect 4919 46073 4985 46096
rect 5071 46073 5153 46096
rect 5239 46073 5305 46096
rect 4919 46054 5305 46073
rect 20039 46159 20425 46178
rect 20039 46136 20105 46159
rect 20191 46136 20273 46159
rect 20359 46136 20425 46159
rect 20039 46096 20048 46136
rect 20088 46096 20105 46136
rect 20191 46096 20212 46136
rect 20252 46096 20273 46136
rect 20359 46096 20376 46136
rect 20416 46096 20425 46136
rect 20039 46073 20105 46096
rect 20191 46073 20273 46096
rect 20359 46073 20425 46096
rect 20039 46054 20425 46073
rect 2090 45991 2214 46010
rect 2090 45905 2109 45991
rect 2195 45968 2214 45991
rect 2195 45928 2380 45968
rect 2420 45928 2429 45968
rect 2195 45905 2214 45928
rect 2090 45886 2214 45905
rect 4579 45676 4588 45716
rect 4628 45676 18028 45716
rect 18068 45676 18077 45716
rect 3679 45403 4065 45422
rect 3679 45380 3745 45403
rect 3831 45380 3913 45403
rect 3999 45380 4065 45403
rect 3679 45340 3688 45380
rect 3728 45340 3745 45380
rect 3831 45340 3852 45380
rect 3892 45340 3913 45380
rect 3999 45340 4016 45380
rect 4056 45340 4065 45380
rect 3679 45317 3745 45340
rect 3831 45317 3913 45340
rect 3999 45317 4065 45340
rect 3679 45298 4065 45317
rect 18799 45403 19185 45422
rect 18799 45380 18865 45403
rect 18951 45380 19033 45403
rect 19119 45380 19185 45403
rect 18799 45340 18808 45380
rect 18848 45340 18865 45380
rect 18951 45340 18972 45380
rect 19012 45340 19033 45380
rect 19119 45340 19136 45380
rect 19176 45340 19185 45380
rect 18799 45317 18865 45340
rect 18951 45317 19033 45340
rect 19119 45317 19185 45340
rect 18799 45298 19185 45317
rect 4675 44920 4684 44960
rect 4724 44920 11404 44960
rect 11444 44920 11453 44960
rect 4919 44647 5305 44666
rect 4919 44624 4985 44647
rect 5071 44624 5153 44647
rect 5239 44624 5305 44647
rect 4919 44584 4928 44624
rect 4968 44584 4985 44624
rect 5071 44584 5092 44624
rect 5132 44584 5153 44624
rect 5239 44584 5256 44624
rect 5296 44584 5305 44624
rect 4919 44561 4985 44584
rect 5071 44561 5153 44584
rect 5239 44561 5305 44584
rect 4919 44542 5305 44561
rect 20039 44647 20425 44666
rect 20039 44624 20105 44647
rect 20191 44624 20273 44647
rect 20359 44624 20425 44647
rect 20039 44584 20048 44624
rect 20088 44584 20105 44624
rect 20191 44584 20212 44624
rect 20252 44584 20273 44624
rect 20359 44584 20376 44624
rect 20416 44584 20425 44624
rect 20039 44561 20105 44584
rect 20191 44561 20273 44584
rect 20359 44561 20425 44584
rect 20039 44542 20425 44561
rect 3679 43891 4065 43910
rect 3679 43868 3745 43891
rect 3831 43868 3913 43891
rect 3999 43868 4065 43891
rect 3679 43828 3688 43868
rect 3728 43828 3745 43868
rect 3831 43828 3852 43868
rect 3892 43828 3913 43868
rect 3999 43828 4016 43868
rect 4056 43828 4065 43868
rect 3679 43805 3745 43828
rect 3831 43805 3913 43828
rect 3999 43805 4065 43828
rect 3679 43786 4065 43805
rect 18799 43891 19185 43910
rect 18799 43868 18865 43891
rect 18951 43868 19033 43891
rect 19119 43868 19185 43891
rect 18799 43828 18808 43868
rect 18848 43828 18865 43868
rect 18951 43828 18972 43868
rect 19012 43828 19033 43868
rect 19119 43828 19136 43868
rect 19176 43828 19185 43868
rect 18799 43805 18865 43828
rect 18951 43805 19033 43828
rect 19119 43805 19185 43828
rect 18799 43786 19185 43805
rect 4919 43135 5305 43154
rect 4919 43112 4985 43135
rect 5071 43112 5153 43135
rect 5239 43112 5305 43135
rect 4919 43072 4928 43112
rect 4968 43072 4985 43112
rect 5071 43072 5092 43112
rect 5132 43072 5153 43112
rect 5239 43072 5256 43112
rect 5296 43072 5305 43112
rect 4919 43049 4985 43072
rect 5071 43049 5153 43072
rect 5239 43049 5305 43072
rect 4919 43030 5305 43049
rect 20039 43135 20425 43154
rect 20039 43112 20105 43135
rect 20191 43112 20273 43135
rect 20359 43112 20425 43135
rect 20039 43072 20048 43112
rect 20088 43072 20105 43112
rect 20191 43072 20212 43112
rect 20252 43072 20273 43112
rect 20359 43072 20376 43112
rect 20416 43072 20425 43112
rect 20039 43049 20105 43072
rect 20191 43049 20273 43072
rect 20359 43049 20425 43072
rect 20039 43030 20425 43049
rect 259 42736 268 42776
rect 308 42736 6604 42776
rect 6644 42736 6653 42776
rect 67 42652 76 42692
rect 116 42652 10732 42692
rect 10772 42652 10781 42692
rect 3679 42379 4065 42398
rect 3679 42356 3745 42379
rect 3831 42356 3913 42379
rect 3999 42356 4065 42379
rect 3679 42316 3688 42356
rect 3728 42316 3745 42356
rect 3831 42316 3852 42356
rect 3892 42316 3913 42356
rect 3999 42316 4016 42356
rect 4056 42316 4065 42356
rect 3679 42293 3745 42316
rect 3831 42293 3913 42316
rect 3999 42293 4065 42316
rect 3679 42274 4065 42293
rect 18799 42379 19185 42398
rect 18799 42356 18865 42379
rect 18951 42356 19033 42379
rect 19119 42356 19185 42379
rect 18799 42316 18808 42356
rect 18848 42316 18865 42356
rect 18951 42316 18972 42356
rect 19012 42316 19033 42356
rect 19119 42316 19136 42356
rect 19176 42316 19185 42356
rect 18799 42293 18865 42316
rect 18951 42293 19033 42316
rect 19119 42293 19185 42316
rect 18799 42274 19185 42293
rect 10298 41959 10422 41978
rect 10298 41936 10317 41959
rect 10147 41896 10156 41936
rect 10196 41896 10317 41936
rect 10298 41873 10317 41896
rect 10403 41873 10422 41959
rect 10298 41854 10422 41873
rect 4919 41623 5305 41642
rect 4919 41600 4985 41623
rect 5071 41600 5153 41623
rect 5239 41600 5305 41623
rect 4919 41560 4928 41600
rect 4968 41560 4985 41600
rect 5071 41560 5092 41600
rect 5132 41560 5153 41600
rect 5239 41560 5256 41600
rect 5296 41560 5305 41600
rect 4919 41537 4985 41560
rect 5071 41537 5153 41560
rect 5239 41537 5305 41560
rect 4919 41518 5305 41537
rect 20039 41623 20425 41642
rect 20039 41600 20105 41623
rect 20191 41600 20273 41623
rect 20359 41600 20425 41623
rect 20039 41560 20048 41600
rect 20088 41560 20105 41600
rect 20191 41560 20212 41600
rect 20252 41560 20273 41600
rect 20359 41560 20376 41600
rect 20416 41560 20425 41600
rect 20039 41537 20105 41560
rect 20191 41537 20273 41560
rect 20359 41537 20425 41560
rect 20039 41518 20425 41537
rect 3679 40867 4065 40886
rect 3679 40844 3745 40867
rect 3831 40844 3913 40867
rect 3999 40844 4065 40867
rect 3679 40804 3688 40844
rect 3728 40804 3745 40844
rect 3831 40804 3852 40844
rect 3892 40804 3913 40844
rect 3999 40804 4016 40844
rect 4056 40804 4065 40844
rect 3679 40781 3745 40804
rect 3831 40781 3913 40804
rect 3999 40781 4065 40804
rect 3679 40762 4065 40781
rect 18799 40867 19185 40886
rect 18799 40844 18865 40867
rect 18951 40844 19033 40867
rect 19119 40844 19185 40867
rect 18799 40804 18808 40844
rect 18848 40804 18865 40844
rect 18951 40804 18972 40844
rect 19012 40804 19033 40844
rect 19119 40804 19136 40844
rect 19176 40804 19185 40844
rect 18799 40781 18865 40804
rect 18951 40781 19033 40804
rect 19119 40781 19185 40804
rect 18799 40762 19185 40781
rect 163 40552 172 40592
rect 212 40552 5548 40592
rect 5588 40552 5597 40592
rect 4919 40111 5305 40130
rect 4919 40088 4985 40111
rect 5071 40088 5153 40111
rect 5239 40088 5305 40111
rect 4919 40048 4928 40088
rect 4968 40048 4985 40088
rect 5071 40048 5092 40088
rect 5132 40048 5153 40088
rect 5239 40048 5256 40088
rect 5296 40048 5305 40088
rect 4919 40025 4985 40048
rect 5071 40025 5153 40048
rect 5239 40025 5305 40048
rect 4919 40006 5305 40025
rect 20039 40111 20425 40130
rect 20039 40088 20105 40111
rect 20191 40088 20273 40111
rect 20359 40088 20425 40111
rect 20039 40048 20048 40088
rect 20088 40048 20105 40088
rect 20191 40048 20212 40088
rect 20252 40048 20273 40088
rect 20359 40048 20376 40088
rect 20416 40048 20425 40088
rect 20039 40025 20105 40048
rect 20191 40025 20273 40048
rect 20359 40025 20425 40048
rect 20039 40006 20425 40025
rect 3679 39355 4065 39374
rect 3679 39332 3745 39355
rect 3831 39332 3913 39355
rect 3999 39332 4065 39355
rect 3679 39292 3688 39332
rect 3728 39292 3745 39332
rect 3831 39292 3852 39332
rect 3892 39292 3913 39332
rect 3999 39292 4016 39332
rect 4056 39292 4065 39332
rect 3679 39269 3745 39292
rect 3831 39269 3913 39292
rect 3999 39269 4065 39292
rect 3679 39250 4065 39269
rect 18799 39355 19185 39374
rect 18799 39332 18865 39355
rect 18951 39332 19033 39355
rect 19119 39332 19185 39355
rect 18799 39292 18808 39332
rect 18848 39292 18865 39332
rect 18951 39292 18972 39332
rect 19012 39292 19033 39332
rect 19119 39292 19136 39332
rect 19176 39292 19185 39332
rect 18799 39269 18865 39292
rect 18951 39269 19033 39292
rect 19119 39269 19185 39292
rect 18799 39250 19185 39269
rect 4919 38599 5305 38618
rect 4919 38576 4985 38599
rect 5071 38576 5153 38599
rect 5239 38576 5305 38599
rect 4919 38536 4928 38576
rect 4968 38536 4985 38576
rect 5071 38536 5092 38576
rect 5132 38536 5153 38576
rect 5239 38536 5256 38576
rect 5296 38536 5305 38576
rect 4919 38513 4985 38536
rect 5071 38513 5153 38536
rect 5239 38513 5305 38536
rect 4919 38494 5305 38513
rect 20039 38599 20425 38618
rect 20039 38576 20105 38599
rect 20191 38576 20273 38599
rect 20359 38576 20425 38599
rect 20039 38536 20048 38576
rect 20088 38536 20105 38576
rect 20191 38536 20212 38576
rect 20252 38536 20273 38576
rect 20359 38536 20376 38576
rect 20416 38536 20425 38576
rect 20039 38513 20105 38536
rect 20191 38513 20273 38536
rect 20359 38513 20425 38536
rect 20039 38494 20425 38513
rect 3679 37843 4065 37862
rect 3679 37820 3745 37843
rect 3831 37820 3913 37843
rect 3999 37820 4065 37843
rect 3679 37780 3688 37820
rect 3728 37780 3745 37820
rect 3831 37780 3852 37820
rect 3892 37780 3913 37820
rect 3999 37780 4016 37820
rect 4056 37780 4065 37820
rect 3679 37757 3745 37780
rect 3831 37757 3913 37780
rect 3999 37757 4065 37780
rect 3679 37738 4065 37757
rect 18799 37843 19185 37862
rect 18799 37820 18865 37843
rect 18951 37820 19033 37843
rect 19119 37820 19185 37843
rect 18799 37780 18808 37820
rect 18848 37780 18865 37820
rect 18951 37780 18972 37820
rect 19012 37780 19033 37820
rect 19119 37780 19136 37820
rect 19176 37780 19185 37820
rect 18799 37757 18865 37780
rect 18951 37757 19033 37780
rect 19119 37757 19185 37780
rect 18799 37738 19185 37757
rect 4919 37087 5305 37106
rect 4919 37064 4985 37087
rect 5071 37064 5153 37087
rect 5239 37064 5305 37087
rect 4919 37024 4928 37064
rect 4968 37024 4985 37064
rect 5071 37024 5092 37064
rect 5132 37024 5153 37064
rect 5239 37024 5256 37064
rect 5296 37024 5305 37064
rect 4919 37001 4985 37024
rect 5071 37001 5153 37024
rect 5239 37001 5305 37024
rect 4919 36982 5305 37001
rect 20039 37087 20425 37106
rect 20039 37064 20105 37087
rect 20191 37064 20273 37087
rect 20359 37064 20425 37087
rect 20039 37024 20048 37064
rect 20088 37024 20105 37064
rect 20191 37024 20212 37064
rect 20252 37024 20273 37064
rect 20359 37024 20376 37064
rect 20416 37024 20425 37064
rect 20039 37001 20105 37024
rect 20191 37001 20273 37024
rect 20359 37001 20425 37024
rect 20039 36982 20425 37001
rect 3679 36331 4065 36350
rect 3679 36308 3745 36331
rect 3831 36308 3913 36331
rect 3999 36308 4065 36331
rect 3679 36268 3688 36308
rect 3728 36268 3745 36308
rect 3831 36268 3852 36308
rect 3892 36268 3913 36308
rect 3999 36268 4016 36308
rect 4056 36268 4065 36308
rect 3679 36245 3745 36268
rect 3831 36245 3913 36268
rect 3999 36245 4065 36268
rect 3679 36226 4065 36245
rect 18799 36331 19185 36350
rect 18799 36308 18865 36331
rect 18951 36308 19033 36331
rect 19119 36308 19185 36331
rect 18799 36268 18808 36308
rect 18848 36268 18865 36308
rect 18951 36268 18972 36308
rect 19012 36268 19033 36308
rect 19119 36268 19136 36308
rect 19176 36268 19185 36308
rect 18799 36245 18865 36268
rect 18951 36245 19033 36268
rect 19119 36245 19185 36268
rect 18799 36226 19185 36245
rect 4919 35575 5305 35594
rect 4919 35552 4985 35575
rect 5071 35552 5153 35575
rect 5239 35552 5305 35575
rect 4919 35512 4928 35552
rect 4968 35512 4985 35552
rect 5071 35512 5092 35552
rect 5132 35512 5153 35552
rect 5239 35512 5256 35552
rect 5296 35512 5305 35552
rect 4919 35489 4985 35512
rect 5071 35489 5153 35512
rect 5239 35489 5305 35512
rect 4919 35470 5305 35489
rect 20039 35575 20425 35594
rect 20039 35552 20105 35575
rect 20191 35552 20273 35575
rect 20359 35552 20425 35575
rect 20039 35512 20048 35552
rect 20088 35512 20105 35552
rect 20191 35512 20212 35552
rect 20252 35512 20273 35552
rect 20359 35512 20376 35552
rect 20416 35512 20425 35552
rect 20039 35489 20105 35512
rect 20191 35489 20273 35512
rect 20359 35489 20425 35512
rect 20039 35470 20425 35489
rect 5347 35176 5356 35216
rect 5396 35176 5836 35216
rect 5876 35176 5885 35216
rect 4483 35008 4492 35048
rect 4532 35008 8236 35048
rect 8276 35008 8285 35048
rect 3679 34819 4065 34838
rect 3679 34796 3745 34819
rect 3831 34796 3913 34819
rect 3999 34796 4065 34819
rect 3679 34756 3688 34796
rect 3728 34756 3745 34796
rect 3831 34756 3852 34796
rect 3892 34756 3913 34796
rect 3999 34756 4016 34796
rect 4056 34756 4065 34796
rect 3679 34733 3745 34756
rect 3831 34733 3913 34756
rect 3999 34733 4065 34756
rect 3679 34714 4065 34733
rect 18799 34819 19185 34838
rect 18799 34796 18865 34819
rect 18951 34796 19033 34819
rect 19119 34796 19185 34819
rect 18799 34756 18808 34796
rect 18848 34756 18865 34796
rect 18951 34756 18972 34796
rect 19012 34756 19033 34796
rect 19119 34756 19136 34796
rect 19176 34756 19185 34796
rect 18799 34733 18865 34756
rect 18951 34733 19033 34756
rect 19119 34733 19185 34756
rect 18799 34714 19185 34733
rect 1178 34399 1302 34418
rect 1178 34313 1197 34399
rect 1283 34376 1302 34399
rect 1283 34336 1324 34376
rect 1364 34336 1373 34376
rect 1283 34313 1302 34336
rect 1178 34294 1302 34313
rect 451 34168 460 34208
rect 500 34168 7564 34208
rect 7604 34168 7613 34208
rect 4919 34063 5305 34082
rect 4919 34040 4985 34063
rect 5071 34040 5153 34063
rect 5239 34040 5305 34063
rect 4919 34000 4928 34040
rect 4968 34000 4985 34040
rect 5071 34000 5092 34040
rect 5132 34000 5153 34040
rect 5239 34000 5256 34040
rect 5296 34000 5305 34040
rect 4919 33977 4985 34000
rect 5071 33977 5153 34000
rect 5239 33977 5305 34000
rect 4919 33958 5305 33977
rect 20039 34063 20425 34082
rect 20039 34040 20105 34063
rect 20191 34040 20273 34063
rect 20359 34040 20425 34063
rect 20039 34000 20048 34040
rect 20088 34000 20105 34040
rect 20191 34000 20212 34040
rect 20252 34000 20273 34040
rect 20359 34000 20376 34040
rect 20416 34000 20425 34040
rect 20039 33977 20105 34000
rect 20191 33977 20273 34000
rect 20359 33977 20425 34000
rect 20039 33958 20425 33977
rect 547 33664 556 33704
rect 596 33664 12556 33704
rect 12596 33664 12605 33704
rect 1219 33496 1228 33536
rect 1268 33496 17068 33536
rect 17108 33496 17117 33536
rect 3679 33307 4065 33326
rect 3679 33284 3745 33307
rect 3831 33284 3913 33307
rect 3999 33284 4065 33307
rect 3679 33244 3688 33284
rect 3728 33244 3745 33284
rect 3831 33244 3852 33284
rect 3892 33244 3913 33284
rect 3999 33244 4016 33284
rect 4056 33244 4065 33284
rect 3679 33221 3745 33244
rect 3831 33221 3913 33244
rect 3999 33221 4065 33244
rect 3679 33202 4065 33221
rect 18799 33307 19185 33326
rect 18799 33284 18865 33307
rect 18951 33284 19033 33307
rect 19119 33284 19185 33307
rect 18799 33244 18808 33284
rect 18848 33244 18865 33284
rect 18951 33244 18972 33284
rect 19012 33244 19033 33284
rect 19119 33244 19136 33284
rect 19176 33244 19185 33284
rect 18799 33221 18865 33244
rect 18951 33221 19033 33244
rect 19119 33221 19185 33244
rect 18799 33202 19185 33221
rect 4919 32551 5305 32570
rect 4919 32528 4985 32551
rect 5071 32528 5153 32551
rect 5239 32528 5305 32551
rect 4919 32488 4928 32528
rect 4968 32488 4985 32528
rect 5071 32488 5092 32528
rect 5132 32488 5153 32528
rect 5239 32488 5256 32528
rect 5296 32488 5305 32528
rect 4919 32465 4985 32488
rect 5071 32465 5153 32488
rect 5239 32465 5305 32488
rect 4919 32446 5305 32465
rect 20039 32551 20425 32570
rect 20039 32528 20105 32551
rect 20191 32528 20273 32551
rect 20359 32528 20425 32551
rect 20039 32488 20048 32528
rect 20088 32488 20105 32528
rect 20191 32488 20212 32528
rect 20252 32488 20273 32528
rect 20359 32488 20376 32528
rect 20416 32488 20425 32528
rect 20039 32465 20105 32488
rect 20191 32465 20273 32488
rect 20359 32465 20425 32488
rect 20039 32446 20425 32465
rect 3679 31795 4065 31814
rect 3679 31772 3745 31795
rect 3831 31772 3913 31795
rect 3999 31772 4065 31795
rect 3679 31732 3688 31772
rect 3728 31732 3745 31772
rect 3831 31732 3852 31772
rect 3892 31732 3913 31772
rect 3999 31732 4016 31772
rect 4056 31732 4065 31772
rect 3679 31709 3745 31732
rect 3831 31709 3913 31732
rect 3999 31709 4065 31732
rect 3679 31690 4065 31709
rect 18799 31795 19185 31814
rect 18799 31772 18865 31795
rect 18951 31772 19033 31795
rect 19119 31772 19185 31795
rect 18799 31732 18808 31772
rect 18848 31732 18865 31772
rect 18951 31732 18972 31772
rect 19012 31732 19033 31772
rect 19119 31732 19136 31772
rect 19176 31732 19185 31772
rect 18799 31709 18865 31732
rect 18951 31709 19033 31732
rect 19119 31709 19185 31732
rect 18799 31690 19185 31709
rect 4919 31039 5305 31058
rect 4919 31016 4985 31039
rect 5071 31016 5153 31039
rect 5239 31016 5305 31039
rect 4919 30976 4928 31016
rect 4968 30976 4985 31016
rect 5071 30976 5092 31016
rect 5132 30976 5153 31016
rect 5239 30976 5256 31016
rect 5296 30976 5305 31016
rect 4919 30953 4985 30976
rect 5071 30953 5153 30976
rect 5239 30953 5305 30976
rect 4919 30934 5305 30953
rect 20039 31039 20425 31058
rect 20039 31016 20105 31039
rect 20191 31016 20273 31039
rect 20359 31016 20425 31039
rect 20039 30976 20048 31016
rect 20088 30976 20105 31016
rect 20191 30976 20212 31016
rect 20252 30976 20273 31016
rect 20359 30976 20376 31016
rect 20416 30976 20425 31016
rect 20039 30953 20105 30976
rect 20191 30953 20273 30976
rect 20359 30953 20425 30976
rect 20039 30934 20425 30953
rect 3679 30283 4065 30302
rect 3679 30260 3745 30283
rect 3831 30260 3913 30283
rect 3999 30260 4065 30283
rect 3679 30220 3688 30260
rect 3728 30220 3745 30260
rect 3831 30220 3852 30260
rect 3892 30220 3913 30260
rect 3999 30220 4016 30260
rect 4056 30220 4065 30260
rect 3679 30197 3745 30220
rect 3831 30197 3913 30220
rect 3999 30197 4065 30220
rect 3679 30178 4065 30197
rect 18799 30283 19185 30302
rect 18799 30260 18865 30283
rect 18951 30260 19033 30283
rect 19119 30260 19185 30283
rect 18799 30220 18808 30260
rect 18848 30220 18865 30260
rect 18951 30220 18972 30260
rect 19012 30220 19033 30260
rect 19119 30220 19136 30260
rect 19176 30220 19185 30260
rect 18799 30197 18865 30220
rect 18951 30197 19033 30220
rect 19119 30197 19185 30220
rect 18799 30178 19185 30197
rect 4919 29527 5305 29546
rect 4919 29504 4985 29527
rect 5071 29504 5153 29527
rect 5239 29504 5305 29527
rect 4919 29464 4928 29504
rect 4968 29464 4985 29504
rect 5071 29464 5092 29504
rect 5132 29464 5153 29504
rect 5239 29464 5256 29504
rect 5296 29464 5305 29504
rect 4919 29441 4985 29464
rect 5071 29441 5153 29464
rect 5239 29441 5305 29464
rect 4919 29422 5305 29441
rect 20039 29527 20425 29546
rect 20039 29504 20105 29527
rect 20191 29504 20273 29527
rect 20359 29504 20425 29527
rect 20039 29464 20048 29504
rect 20088 29464 20105 29504
rect 20191 29464 20212 29504
rect 20252 29464 20273 29504
rect 20359 29464 20376 29504
rect 20416 29464 20425 29504
rect 20039 29441 20105 29464
rect 20191 29441 20273 29464
rect 20359 29441 20425 29464
rect 20039 29422 20425 29441
rect 17635 29380 17644 29420
rect 17684 29380 17932 29420
rect 17972 29380 17981 29420
rect 3679 28771 4065 28790
rect 3679 28748 3745 28771
rect 3831 28748 3913 28771
rect 3999 28748 4065 28771
rect 3679 28708 3688 28748
rect 3728 28708 3745 28748
rect 3831 28708 3852 28748
rect 3892 28708 3913 28748
rect 3999 28708 4016 28748
rect 4056 28708 4065 28748
rect 3679 28685 3745 28708
rect 3831 28685 3913 28708
rect 3999 28685 4065 28708
rect 3679 28666 4065 28685
rect 18799 28771 19185 28790
rect 18799 28748 18865 28771
rect 18951 28748 19033 28771
rect 19119 28748 19185 28771
rect 18799 28708 18808 28748
rect 18848 28708 18865 28748
rect 18951 28708 18972 28748
rect 19012 28708 19033 28748
rect 19119 28708 19136 28748
rect 19176 28708 19185 28748
rect 18799 28685 18865 28708
rect 18951 28685 19033 28708
rect 19119 28685 19185 28708
rect 18799 28666 19185 28685
rect 17059 28456 17068 28496
rect 17108 28456 17260 28496
rect 17300 28456 17309 28496
rect 4919 28015 5305 28034
rect 4919 27992 4985 28015
rect 5071 27992 5153 28015
rect 5239 27992 5305 28015
rect 4919 27952 4928 27992
rect 4968 27952 4985 27992
rect 5071 27952 5092 27992
rect 5132 27952 5153 27992
rect 5239 27952 5256 27992
rect 5296 27952 5305 27992
rect 4919 27929 4985 27952
rect 5071 27929 5153 27952
rect 5239 27929 5305 27952
rect 4919 27910 5305 27929
rect 20039 28015 20425 28034
rect 20039 27992 20105 28015
rect 20191 27992 20273 28015
rect 20359 27992 20425 28015
rect 20039 27952 20048 27992
rect 20088 27952 20105 27992
rect 20191 27952 20212 27992
rect 20252 27952 20273 27992
rect 20359 27952 20376 27992
rect 20416 27952 20425 27992
rect 20039 27929 20105 27952
rect 20191 27929 20273 27952
rect 20359 27929 20425 27952
rect 20039 27910 20425 27929
rect 3679 27259 4065 27278
rect 3679 27236 3745 27259
rect 3831 27236 3913 27259
rect 3999 27236 4065 27259
rect 3679 27196 3688 27236
rect 3728 27196 3745 27236
rect 3831 27196 3852 27236
rect 3892 27196 3913 27236
rect 3999 27196 4016 27236
rect 4056 27196 4065 27236
rect 3679 27173 3745 27196
rect 3831 27173 3913 27196
rect 3999 27173 4065 27196
rect 3679 27154 4065 27173
rect 18799 27259 19185 27278
rect 18799 27236 18865 27259
rect 18951 27236 19033 27259
rect 19119 27236 19185 27259
rect 18799 27196 18808 27236
rect 18848 27196 18865 27236
rect 18951 27196 18972 27236
rect 19012 27196 19033 27236
rect 19119 27196 19136 27236
rect 19176 27196 19185 27236
rect 18799 27173 18865 27196
rect 18951 27173 19033 27196
rect 19119 27173 19185 27196
rect 18799 27154 19185 27173
rect 4919 26503 5305 26522
rect 4919 26480 4985 26503
rect 5071 26480 5153 26503
rect 5239 26480 5305 26503
rect 4919 26440 4928 26480
rect 4968 26440 4985 26480
rect 5071 26440 5092 26480
rect 5132 26440 5153 26480
rect 5239 26440 5256 26480
rect 5296 26440 5305 26480
rect 4919 26417 4985 26440
rect 5071 26417 5153 26440
rect 5239 26417 5305 26440
rect 4919 26398 5305 26417
rect 20039 26503 20425 26522
rect 20039 26480 20105 26503
rect 20191 26480 20273 26503
rect 20359 26480 20425 26503
rect 20039 26440 20048 26480
rect 20088 26440 20105 26480
rect 20191 26440 20212 26480
rect 20252 26440 20273 26480
rect 20359 26440 20376 26480
rect 20416 26440 20425 26480
rect 20039 26417 20105 26440
rect 20191 26417 20273 26440
rect 20359 26417 20425 26440
rect 20039 26398 20425 26417
rect 1411 26272 1420 26312
rect 1460 26272 5932 26312
rect 5972 26272 5981 26312
rect 1315 26104 1324 26144
rect 1364 26104 19756 26144
rect 19796 26104 19805 26144
rect 3679 25747 4065 25766
rect 3679 25724 3745 25747
rect 3831 25724 3913 25747
rect 3999 25724 4065 25747
rect 3679 25684 3688 25724
rect 3728 25684 3745 25724
rect 3831 25684 3852 25724
rect 3892 25684 3913 25724
rect 3999 25684 4016 25724
rect 4056 25684 4065 25724
rect 3679 25661 3745 25684
rect 3831 25661 3913 25684
rect 3999 25661 4065 25684
rect 3679 25642 4065 25661
rect 18799 25747 19185 25766
rect 18799 25724 18865 25747
rect 18951 25724 19033 25747
rect 19119 25724 19185 25747
rect 18799 25684 18808 25724
rect 18848 25684 18865 25724
rect 18951 25684 18972 25724
rect 19012 25684 19033 25724
rect 19119 25684 19136 25724
rect 19176 25684 19185 25724
rect 18799 25661 18865 25684
rect 18951 25661 19033 25684
rect 19119 25661 19185 25684
rect 18799 25642 19185 25661
rect 4919 24991 5305 25010
rect 4919 24968 4985 24991
rect 5071 24968 5153 24991
rect 5239 24968 5305 24991
rect 4919 24928 4928 24968
rect 4968 24928 4985 24968
rect 5071 24928 5092 24968
rect 5132 24928 5153 24968
rect 5239 24928 5256 24968
rect 5296 24928 5305 24968
rect 4919 24905 4985 24928
rect 5071 24905 5153 24928
rect 5239 24905 5305 24928
rect 4919 24886 5305 24905
rect 20039 24991 20425 25010
rect 20039 24968 20105 24991
rect 20191 24968 20273 24991
rect 20359 24968 20425 24991
rect 20039 24928 20048 24968
rect 20088 24928 20105 24968
rect 20191 24928 20212 24968
rect 20252 24928 20273 24968
rect 20359 24928 20376 24968
rect 20416 24928 20425 24968
rect 20039 24905 20105 24928
rect 20191 24905 20273 24928
rect 20359 24905 20425 24928
rect 20039 24886 20425 24905
rect 16226 24655 16350 24674
rect 16226 24569 16245 24655
rect 16331 24632 16350 24655
rect 16331 24592 18316 24632
rect 18356 24592 18365 24632
rect 16331 24569 16350 24592
rect 16226 24550 16350 24569
rect 3679 24235 4065 24254
rect 3679 24212 3745 24235
rect 3831 24212 3913 24235
rect 3999 24212 4065 24235
rect 3679 24172 3688 24212
rect 3728 24172 3745 24212
rect 3831 24172 3852 24212
rect 3892 24172 3913 24212
rect 3999 24172 4016 24212
rect 4056 24172 4065 24212
rect 3679 24149 3745 24172
rect 3831 24149 3913 24172
rect 3999 24149 4065 24172
rect 3679 24130 4065 24149
rect 18799 24235 19185 24254
rect 18799 24212 18865 24235
rect 18951 24212 19033 24235
rect 19119 24212 19185 24235
rect 18799 24172 18808 24212
rect 18848 24172 18865 24212
rect 18951 24172 18972 24212
rect 19012 24172 19033 24212
rect 19119 24172 19136 24212
rect 19176 24172 19185 24212
rect 18799 24149 18865 24172
rect 18951 24149 19033 24172
rect 19119 24149 19185 24172
rect 18799 24130 19185 24149
rect 4919 23479 5305 23498
rect 4919 23456 4985 23479
rect 5071 23456 5153 23479
rect 5239 23456 5305 23479
rect 4919 23416 4928 23456
rect 4968 23416 4985 23456
rect 5071 23416 5092 23456
rect 5132 23416 5153 23456
rect 5239 23416 5256 23456
rect 5296 23416 5305 23456
rect 4919 23393 4985 23416
rect 5071 23393 5153 23416
rect 5239 23393 5305 23416
rect 4919 23374 5305 23393
rect 20039 23479 20425 23498
rect 20039 23456 20105 23479
rect 20191 23456 20273 23479
rect 20359 23456 20425 23479
rect 20039 23416 20048 23456
rect 20088 23416 20105 23456
rect 20191 23416 20212 23456
rect 20252 23416 20273 23456
rect 20359 23416 20376 23456
rect 20416 23416 20425 23456
rect 20039 23393 20105 23416
rect 20191 23393 20273 23416
rect 20359 23393 20425 23416
rect 20039 23374 20425 23393
rect 3679 22723 4065 22742
rect 3679 22700 3745 22723
rect 3831 22700 3913 22723
rect 3999 22700 4065 22723
rect 3679 22660 3688 22700
rect 3728 22660 3745 22700
rect 3831 22660 3852 22700
rect 3892 22660 3913 22700
rect 3999 22660 4016 22700
rect 4056 22660 4065 22700
rect 3679 22637 3745 22660
rect 3831 22637 3913 22660
rect 3999 22637 4065 22660
rect 3679 22618 4065 22637
rect 18799 22723 19185 22742
rect 18799 22700 18865 22723
rect 18951 22700 19033 22723
rect 19119 22700 19185 22723
rect 18799 22660 18808 22700
rect 18848 22660 18865 22700
rect 18951 22660 18972 22700
rect 19012 22660 19033 22700
rect 19119 22660 19136 22700
rect 19176 22660 19185 22700
rect 18799 22637 18865 22660
rect 18951 22637 19033 22660
rect 19119 22637 19185 22660
rect 18799 22618 19185 22637
rect 547 22072 556 22112
rect 596 22072 748 22112
rect 788 22072 797 22112
rect 4919 21967 5305 21986
rect 4919 21944 4985 21967
rect 5071 21944 5153 21967
rect 5239 21944 5305 21967
rect 4919 21904 4928 21944
rect 4968 21904 4985 21944
rect 5071 21904 5092 21944
rect 5132 21904 5153 21944
rect 5239 21904 5256 21944
rect 5296 21904 5305 21944
rect 4919 21881 4985 21904
rect 5071 21881 5153 21904
rect 5239 21881 5305 21904
rect 4919 21862 5305 21881
rect 20039 21967 20425 21986
rect 20039 21944 20105 21967
rect 20191 21944 20273 21967
rect 20359 21944 20425 21967
rect 20039 21904 20048 21944
rect 20088 21904 20105 21944
rect 20191 21904 20212 21944
rect 20252 21904 20273 21944
rect 20359 21904 20376 21944
rect 20416 21904 20425 21944
rect 20039 21881 20105 21904
rect 20191 21881 20273 21904
rect 20359 21881 20425 21904
rect 20039 21862 20425 21881
rect 1219 21400 1228 21440
rect 1268 21400 10444 21440
rect 10484 21400 10493 21440
rect 3679 21211 4065 21230
rect 3679 21188 3745 21211
rect 3831 21188 3913 21211
rect 3999 21188 4065 21211
rect 3679 21148 3688 21188
rect 3728 21148 3745 21188
rect 3831 21148 3852 21188
rect 3892 21148 3913 21188
rect 3999 21148 4016 21188
rect 4056 21148 4065 21188
rect 3679 21125 3745 21148
rect 3831 21125 3913 21148
rect 3999 21125 4065 21148
rect 3679 21106 4065 21125
rect 18799 21211 19185 21230
rect 18799 21188 18865 21211
rect 18951 21188 19033 21211
rect 19119 21188 19185 21211
rect 18799 21148 18808 21188
rect 18848 21148 18865 21188
rect 18951 21148 18972 21188
rect 19012 21148 19033 21188
rect 19119 21148 19136 21188
rect 19176 21148 19185 21188
rect 18799 21125 18865 21148
rect 18951 21125 19033 21148
rect 19119 21125 19185 21148
rect 18799 21106 19185 21125
rect 4919 20455 5305 20474
rect 4919 20432 4985 20455
rect 5071 20432 5153 20455
rect 5239 20432 5305 20455
rect 4919 20392 4928 20432
rect 4968 20392 4985 20432
rect 5071 20392 5092 20432
rect 5132 20392 5153 20432
rect 5239 20392 5256 20432
rect 5296 20392 5305 20432
rect 4919 20369 4985 20392
rect 5071 20369 5153 20392
rect 5239 20369 5305 20392
rect 4919 20350 5305 20369
rect 20039 20455 20425 20474
rect 20039 20432 20105 20455
rect 20191 20432 20273 20455
rect 20359 20432 20425 20455
rect 20039 20392 20048 20432
rect 20088 20392 20105 20432
rect 20191 20392 20212 20432
rect 20252 20392 20273 20432
rect 20359 20392 20376 20432
rect 20416 20392 20425 20432
rect 20039 20369 20105 20392
rect 20191 20369 20273 20392
rect 20359 20369 20425 20392
rect 20039 20350 20425 20369
rect 3679 19699 4065 19718
rect 3679 19676 3745 19699
rect 3831 19676 3913 19699
rect 3999 19676 4065 19699
rect 3679 19636 3688 19676
rect 3728 19636 3745 19676
rect 3831 19636 3852 19676
rect 3892 19636 3913 19676
rect 3999 19636 4016 19676
rect 4056 19636 4065 19676
rect 3679 19613 3745 19636
rect 3831 19613 3913 19636
rect 3999 19613 4065 19636
rect 3679 19594 4065 19613
rect 18799 19699 19185 19718
rect 18799 19676 18865 19699
rect 18951 19676 19033 19699
rect 19119 19676 19185 19699
rect 18799 19636 18808 19676
rect 18848 19636 18865 19676
rect 18951 19636 18972 19676
rect 19012 19636 19033 19676
rect 19119 19636 19136 19676
rect 19176 19636 19185 19676
rect 18799 19613 18865 19636
rect 18951 19613 19033 19636
rect 19119 19613 19185 19636
rect 18799 19594 19185 19613
rect 4919 18943 5305 18962
rect 4919 18920 4985 18943
rect 5071 18920 5153 18943
rect 5239 18920 5305 18943
rect 4919 18880 4928 18920
rect 4968 18880 4985 18920
rect 5071 18880 5092 18920
rect 5132 18880 5153 18920
rect 5239 18880 5256 18920
rect 5296 18880 5305 18920
rect 4919 18857 4985 18880
rect 5071 18857 5153 18880
rect 5239 18857 5305 18880
rect 4919 18838 5305 18857
rect 20039 18943 20425 18962
rect 20039 18920 20105 18943
rect 20191 18920 20273 18943
rect 20359 18920 20425 18943
rect 20039 18880 20048 18920
rect 20088 18880 20105 18920
rect 20191 18880 20212 18920
rect 20252 18880 20273 18920
rect 20359 18880 20376 18920
rect 20416 18880 20425 18920
rect 20039 18857 20105 18880
rect 20191 18857 20273 18880
rect 20359 18857 20425 18880
rect 20039 18838 20425 18857
rect 1219 18712 1228 18752
rect 1268 18712 7948 18752
rect 7988 18712 7997 18752
rect 3715 18544 3724 18584
rect 3764 18544 9676 18584
rect 9716 18544 9725 18584
rect 1219 18292 1228 18332
rect 1268 18292 8428 18332
rect 8468 18292 8477 18332
rect 3679 18187 4065 18206
rect 3679 18164 3745 18187
rect 3831 18164 3913 18187
rect 3999 18164 4065 18187
rect 3679 18124 3688 18164
rect 3728 18124 3745 18164
rect 3831 18124 3852 18164
rect 3892 18124 3913 18164
rect 3999 18124 4016 18164
rect 4056 18124 4065 18164
rect 3679 18101 3745 18124
rect 3831 18101 3913 18124
rect 3999 18101 4065 18124
rect 3679 18082 4065 18101
rect 18799 18187 19185 18206
rect 18799 18164 18865 18187
rect 18951 18164 19033 18187
rect 19119 18164 19185 18187
rect 18799 18124 18808 18164
rect 18848 18124 18865 18164
rect 18951 18124 18972 18164
rect 19012 18124 19033 18164
rect 19119 18124 19136 18164
rect 19176 18124 19185 18164
rect 18799 18101 18865 18124
rect 18951 18101 19033 18124
rect 19119 18101 19185 18124
rect 18799 18082 19185 18101
rect 5059 17704 5068 17744
rect 5108 17704 11308 17744
rect 11348 17704 11357 17744
rect 13490 17683 13614 17702
rect 13490 17597 13509 17683
rect 13595 17660 13614 17683
rect 13595 17620 15724 17660
rect 15764 17620 15773 17660
rect 13595 17597 13614 17620
rect 13490 17578 13614 17597
rect 8995 17536 9004 17576
rect 9044 17536 9292 17576
rect 9332 17536 9341 17576
rect 4919 17431 5305 17450
rect 4919 17408 4985 17431
rect 5071 17408 5153 17431
rect 5239 17408 5305 17431
rect 4919 17368 4928 17408
rect 4968 17368 4985 17408
rect 5071 17368 5092 17408
rect 5132 17368 5153 17408
rect 5239 17368 5256 17408
rect 5296 17368 5305 17408
rect 4919 17345 4985 17368
rect 5071 17345 5153 17368
rect 5239 17345 5305 17368
rect 4919 17326 5305 17345
rect 20039 17431 20425 17450
rect 20039 17408 20105 17431
rect 20191 17408 20273 17431
rect 20359 17408 20425 17431
rect 20039 17368 20048 17408
rect 20088 17368 20105 17408
rect 20191 17368 20212 17408
rect 20252 17368 20273 17408
rect 20359 17368 20376 17408
rect 20416 17368 20425 17408
rect 20039 17345 20105 17368
rect 20191 17345 20273 17368
rect 20359 17345 20425 17368
rect 20039 17326 20425 17345
rect 931 16780 940 16820
rect 980 16780 6316 16820
rect 6356 16780 6365 16820
rect 15715 16780 15724 16820
rect 15764 16780 20812 16820
rect 20852 16780 20861 16820
rect 3679 16675 4065 16694
rect 3679 16652 3745 16675
rect 3831 16652 3913 16675
rect 3999 16652 4065 16675
rect 3679 16612 3688 16652
rect 3728 16612 3745 16652
rect 3831 16612 3852 16652
rect 3892 16612 3913 16652
rect 3999 16612 4016 16652
rect 4056 16612 4065 16652
rect 3679 16589 3745 16612
rect 3831 16589 3913 16612
rect 3999 16589 4065 16612
rect 3679 16570 4065 16589
rect 18799 16675 19185 16694
rect 18799 16652 18865 16675
rect 18951 16652 19033 16675
rect 19119 16652 19185 16675
rect 18799 16612 18808 16652
rect 18848 16612 18865 16652
rect 18951 16612 18972 16652
rect 19012 16612 19033 16652
rect 19119 16612 19136 16652
rect 19176 16612 19185 16652
rect 18799 16589 18865 16612
rect 18951 16589 19033 16612
rect 19119 16589 19185 16612
rect 18799 16570 19185 16589
rect 643 16360 652 16400
rect 692 16360 2956 16400
rect 2996 16360 4876 16400
rect 4916 16360 4925 16400
rect 4919 15919 5305 15938
rect 4919 15896 4985 15919
rect 5071 15896 5153 15919
rect 5239 15896 5305 15919
rect 4919 15856 4928 15896
rect 4968 15856 4985 15896
rect 5071 15856 5092 15896
rect 5132 15856 5153 15896
rect 5239 15856 5256 15896
rect 5296 15856 5305 15896
rect 4919 15833 4985 15856
rect 5071 15833 5153 15856
rect 5239 15833 5305 15856
rect 4919 15814 5305 15833
rect 20039 15919 20425 15938
rect 20039 15896 20105 15919
rect 20191 15896 20273 15919
rect 20359 15896 20425 15919
rect 20039 15856 20048 15896
rect 20088 15856 20105 15896
rect 20191 15856 20212 15896
rect 20252 15856 20273 15896
rect 20359 15856 20376 15896
rect 20416 15856 20425 15896
rect 20039 15833 20105 15856
rect 20191 15833 20273 15856
rect 20359 15833 20425 15856
rect 20039 15814 20425 15833
rect 14858 15751 14982 15770
rect 14858 15728 14877 15751
rect 13123 15688 13132 15728
rect 13172 15688 14877 15728
rect 14858 15665 14877 15688
rect 14963 15665 14982 15751
rect 14858 15646 14982 15665
rect 16387 15520 16396 15560
rect 16436 15520 20140 15560
rect 20180 15520 20189 15560
rect 3679 15163 4065 15182
rect 3679 15140 3745 15163
rect 3831 15140 3913 15163
rect 3999 15140 4065 15163
rect 3679 15100 3688 15140
rect 3728 15100 3745 15140
rect 3831 15100 3852 15140
rect 3892 15100 3913 15140
rect 3999 15100 4016 15140
rect 4056 15100 4065 15140
rect 3679 15077 3745 15100
rect 3831 15077 3913 15100
rect 3999 15077 4065 15100
rect 3679 15058 4065 15077
rect 18799 15163 19185 15182
rect 18799 15140 18865 15163
rect 18951 15140 19033 15163
rect 19119 15140 19185 15163
rect 18799 15100 18808 15140
rect 18848 15100 18865 15140
rect 18951 15100 18972 15140
rect 19012 15100 19033 15140
rect 19119 15100 19136 15140
rect 19176 15100 19185 15140
rect 18799 15077 18865 15100
rect 18951 15077 19033 15100
rect 19119 15077 19185 15100
rect 18799 15058 19185 15077
rect 8611 14512 8620 14552
rect 8660 14512 15148 14552
rect 15188 14512 15197 14552
rect 4919 14407 5305 14426
rect 4919 14384 4985 14407
rect 5071 14384 5153 14407
rect 5239 14384 5305 14407
rect 4919 14344 4928 14384
rect 4968 14344 4985 14384
rect 5071 14344 5092 14384
rect 5132 14344 5153 14384
rect 5239 14344 5256 14384
rect 5296 14344 5305 14384
rect 4919 14321 4985 14344
rect 5071 14321 5153 14344
rect 5239 14321 5305 14344
rect 4919 14302 5305 14321
rect 20039 14407 20425 14426
rect 20039 14384 20105 14407
rect 20191 14384 20273 14407
rect 20359 14384 20425 14407
rect 20039 14344 20048 14384
rect 20088 14344 20105 14384
rect 20191 14344 20212 14384
rect 20252 14344 20273 14384
rect 20359 14344 20376 14384
rect 20416 14344 20425 14384
rect 20039 14321 20105 14344
rect 20191 14321 20273 14344
rect 20359 14321 20425 14344
rect 20039 14302 20425 14321
rect 3679 13651 4065 13670
rect 3679 13628 3745 13651
rect 3831 13628 3913 13651
rect 3999 13628 4065 13651
rect 3679 13588 3688 13628
rect 3728 13588 3745 13628
rect 3831 13588 3852 13628
rect 3892 13588 3913 13628
rect 3999 13588 4016 13628
rect 4056 13588 4065 13628
rect 3679 13565 3745 13588
rect 3831 13565 3913 13588
rect 3999 13565 4065 13588
rect 3679 13546 4065 13565
rect 18799 13651 19185 13670
rect 18799 13628 18865 13651
rect 18951 13628 19033 13651
rect 19119 13628 19185 13651
rect 18799 13588 18808 13628
rect 18848 13588 18865 13628
rect 18951 13588 18972 13628
rect 19012 13588 19033 13628
rect 19119 13588 19136 13628
rect 19176 13588 19185 13628
rect 18799 13565 18865 13588
rect 18951 13565 19033 13588
rect 19119 13565 19185 13588
rect 18799 13546 19185 13565
rect 8995 13168 9004 13208
rect 9044 13168 9292 13208
rect 9332 13168 9341 13208
rect 4919 12895 5305 12914
rect 4919 12872 4985 12895
rect 5071 12872 5153 12895
rect 5239 12872 5305 12895
rect 4919 12832 4928 12872
rect 4968 12832 4985 12872
rect 5071 12832 5092 12872
rect 5132 12832 5153 12872
rect 5239 12832 5256 12872
rect 5296 12832 5305 12872
rect 4919 12809 4985 12832
rect 5071 12809 5153 12832
rect 5239 12809 5305 12832
rect 4919 12790 5305 12809
rect 20039 12895 20425 12914
rect 20039 12872 20105 12895
rect 20191 12872 20273 12895
rect 20359 12872 20425 12895
rect 20039 12832 20048 12872
rect 20088 12832 20105 12872
rect 20191 12832 20212 12872
rect 20252 12832 20273 12872
rect 20359 12832 20376 12872
rect 20416 12832 20425 12872
rect 20039 12809 20105 12832
rect 20191 12809 20273 12832
rect 20359 12809 20425 12832
rect 20039 12790 20425 12809
rect 3427 12496 3436 12536
rect 3476 12496 3820 12536
rect 3860 12496 3869 12536
rect 3679 12139 4065 12158
rect 3679 12116 3745 12139
rect 3831 12116 3913 12139
rect 3999 12116 4065 12139
rect 3679 12076 3688 12116
rect 3728 12076 3745 12116
rect 3831 12076 3852 12116
rect 3892 12076 3913 12116
rect 3999 12076 4016 12116
rect 4056 12076 4065 12116
rect 3679 12053 3745 12076
rect 3831 12053 3913 12076
rect 3999 12053 4065 12076
rect 3679 12034 4065 12053
rect 18799 12139 19185 12158
rect 18799 12116 18865 12139
rect 18951 12116 19033 12139
rect 19119 12116 19185 12139
rect 18799 12076 18808 12116
rect 18848 12076 18865 12116
rect 18951 12076 18972 12116
rect 19012 12076 19033 12116
rect 19119 12076 19136 12116
rect 19176 12076 19185 12116
rect 18799 12053 18865 12076
rect 18951 12053 19033 12076
rect 19119 12053 19185 12076
rect 18799 12034 19185 12053
rect 4919 11383 5305 11402
rect 4919 11360 4985 11383
rect 5071 11360 5153 11383
rect 5239 11360 5305 11383
rect 4919 11320 4928 11360
rect 4968 11320 4985 11360
rect 5071 11320 5092 11360
rect 5132 11320 5153 11360
rect 5239 11320 5256 11360
rect 5296 11320 5305 11360
rect 4919 11297 4985 11320
rect 5071 11297 5153 11320
rect 5239 11297 5305 11320
rect 4919 11278 5305 11297
rect 20039 11383 20425 11402
rect 20039 11360 20105 11383
rect 20191 11360 20273 11383
rect 20359 11360 20425 11383
rect 20039 11320 20048 11360
rect 20088 11320 20105 11360
rect 20191 11320 20212 11360
rect 20252 11320 20273 11360
rect 20359 11320 20376 11360
rect 20416 11320 20425 11360
rect 20039 11297 20105 11320
rect 20191 11297 20273 11320
rect 20359 11297 20425 11320
rect 20039 11278 20425 11297
rect 10723 11236 10732 11276
rect 10772 11236 15852 11276
rect 15812 11192 15852 11236
rect 15812 11152 20140 11192
rect 20180 11152 20189 11192
rect 8474 11131 8598 11150
rect 8474 11045 8493 11131
rect 8579 11108 8598 11131
rect 8579 11068 13036 11108
rect 13076 11068 13085 11108
rect 8579 11045 8598 11068
rect 8474 11026 8598 11045
rect 3679 10627 4065 10646
rect 3679 10604 3745 10627
rect 3831 10604 3913 10627
rect 3999 10604 4065 10627
rect 3679 10564 3688 10604
rect 3728 10564 3745 10604
rect 3831 10564 3852 10604
rect 3892 10564 3913 10604
rect 3999 10564 4016 10604
rect 4056 10564 4065 10604
rect 3679 10541 3745 10564
rect 3831 10541 3913 10564
rect 3999 10541 4065 10564
rect 3679 10522 4065 10541
rect 18799 10627 19185 10646
rect 18799 10604 18865 10627
rect 18951 10604 19033 10627
rect 19119 10604 19185 10627
rect 18799 10564 18808 10604
rect 18848 10564 18865 10604
rect 18951 10564 18972 10604
rect 19012 10564 19033 10604
rect 19119 10564 19136 10604
rect 19176 10564 19185 10604
rect 18799 10541 18865 10564
rect 18951 10541 19033 10564
rect 19119 10541 19185 10564
rect 18799 10522 19185 10541
rect 12067 10396 12076 10436
rect 12116 10396 18220 10436
rect 18260 10396 18269 10436
rect 9386 10291 9510 10310
rect 9386 10205 9405 10291
rect 9491 10268 9510 10291
rect 9491 10228 9964 10268
rect 10004 10228 10013 10268
rect 9491 10205 9510 10228
rect 9386 10186 9510 10205
rect 5539 9976 5548 10016
rect 5588 9976 20812 10016
rect 20852 9976 20861 10016
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 3715 8884 3724 8924
rect 3764 8884 4204 8924
rect 4244 8884 4253 8924
rect 2659 8800 2668 8840
rect 2708 8800 20140 8840
rect 20180 8800 20189 8840
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 14755 7120 14764 7160
rect 14804 7120 20140 7160
rect 20180 7120 20189 7160
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 4919 5230 5305 5249
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 13490 2731 13614 2750
rect 13490 2645 13509 2731
rect 13595 2708 13614 2731
rect 13595 2668 13804 2708
rect 13844 2668 13853 2708
rect 13595 2645 13614 2668
rect 13490 2626 13614 2645
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 2090 2143 2214 2162
rect 2090 2057 2109 2143
rect 2195 2120 2214 2143
rect 7106 2143 7230 2162
rect 2195 2080 5740 2120
rect 5780 2080 5789 2120
rect 2195 2057 2214 2080
rect 2090 2038 2214 2057
rect 7106 2057 7125 2143
rect 7211 2120 7230 2143
rect 12122 2143 12246 2162
rect 7211 2080 7276 2120
rect 7316 2080 7325 2120
rect 7211 2057 7230 2080
rect 7106 2038 7230 2057
rect 12122 2057 12141 2143
rect 12227 2120 12246 2143
rect 12227 2080 19564 2120
rect 19604 2080 19613 2120
rect 12227 2057 12246 2080
rect 12122 2038 12246 2057
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 3679 1450 4065 1469
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 7843 1240 7852 1280
rect 7892 1240 11360 1280
rect 11320 1196 11360 1240
rect 11320 1156 13420 1196
rect 13460 1156 13469 1196
rect 17138 967 17262 986
rect 17138 881 17157 967
rect 17243 944 17262 967
rect 17243 904 19180 944
rect 19220 904 19229 944
rect 17243 881 17262 904
rect 17138 862 17262 881
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 4919 694 5305 713
rect 20039 799 20425 818
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
rect 5059 232 5068 272
rect 5108 232 8908 272
rect 8948 232 8957 272
rect 10298 211 10422 230
rect 10298 188 10317 211
rect 4867 148 4876 188
rect 4916 148 10317 188
rect 10298 125 10317 148
rect 10403 125 10422 211
rect 10298 106 10422 125
rect 3331 64 3340 104
rect 3380 64 9100 104
rect 9140 64 9149 104
<< via5 >>
rect 12141 85805 12227 85891
rect 17157 85721 17243 85807
rect 16245 85049 16331 85135
rect 3745 84692 3831 84715
rect 3913 84692 3999 84715
rect 3745 84652 3770 84692
rect 3770 84652 3810 84692
rect 3810 84652 3831 84692
rect 3913 84652 3934 84692
rect 3934 84652 3974 84692
rect 3974 84652 3999 84692
rect 3745 84629 3831 84652
rect 3913 84629 3999 84652
rect 18865 84692 18951 84715
rect 19033 84692 19119 84715
rect 18865 84652 18890 84692
rect 18890 84652 18930 84692
rect 18930 84652 18951 84692
rect 19033 84652 19054 84692
rect 19054 84652 19094 84692
rect 19094 84652 19119 84692
rect 18865 84629 18951 84652
rect 19033 84629 19119 84652
rect 7125 84377 7211 84463
rect 14877 84377 14963 84463
rect 4985 83936 5071 83959
rect 5153 83936 5239 83959
rect 4985 83896 5010 83936
rect 5010 83896 5050 83936
rect 5050 83896 5071 83936
rect 5153 83896 5174 83936
rect 5174 83896 5214 83936
rect 5214 83896 5239 83936
rect 4985 83873 5071 83896
rect 5153 83873 5239 83896
rect 20105 83936 20191 83959
rect 20273 83936 20359 83959
rect 20105 83896 20130 83936
rect 20130 83896 20170 83936
rect 20170 83896 20191 83936
rect 20273 83896 20294 83936
rect 20294 83896 20334 83936
rect 20334 83896 20359 83936
rect 20105 83873 20191 83896
rect 20273 83873 20359 83896
rect 2109 83453 2195 83539
rect 3745 83180 3831 83203
rect 3913 83180 3999 83203
rect 3745 83140 3770 83180
rect 3770 83140 3810 83180
rect 3810 83140 3831 83180
rect 3913 83140 3934 83180
rect 3934 83140 3974 83180
rect 3974 83140 3999 83180
rect 3745 83117 3831 83140
rect 3913 83117 3999 83140
rect 18865 83180 18951 83203
rect 19033 83180 19119 83203
rect 18865 83140 18890 83180
rect 18890 83140 18930 83180
rect 18930 83140 18951 83180
rect 19033 83140 19054 83180
rect 19054 83140 19094 83180
rect 19094 83140 19119 83180
rect 18865 83117 18951 83140
rect 19033 83117 19119 83140
rect 4985 82424 5071 82447
rect 5153 82424 5239 82447
rect 4985 82384 5010 82424
rect 5010 82384 5050 82424
rect 5050 82384 5071 82424
rect 5153 82384 5174 82424
rect 5174 82384 5214 82424
rect 5214 82384 5239 82424
rect 4985 82361 5071 82384
rect 5153 82361 5239 82384
rect 20105 82424 20191 82447
rect 20273 82424 20359 82447
rect 20105 82384 20130 82424
rect 20130 82384 20170 82424
rect 20170 82384 20191 82424
rect 20273 82384 20294 82424
rect 20294 82384 20334 82424
rect 20334 82384 20359 82424
rect 20105 82361 20191 82384
rect 20273 82361 20359 82384
rect 3745 81668 3831 81691
rect 3913 81668 3999 81691
rect 3745 81628 3770 81668
rect 3770 81628 3810 81668
rect 3810 81628 3831 81668
rect 3913 81628 3934 81668
rect 3934 81628 3974 81668
rect 3974 81628 3999 81668
rect 3745 81605 3831 81628
rect 3913 81605 3999 81628
rect 18865 81668 18951 81691
rect 19033 81668 19119 81691
rect 18865 81628 18890 81668
rect 18890 81628 18930 81668
rect 18930 81628 18951 81668
rect 19033 81628 19054 81668
rect 19054 81628 19094 81668
rect 19094 81628 19119 81668
rect 18865 81605 18951 81628
rect 19033 81605 19119 81628
rect 4985 80912 5071 80935
rect 5153 80912 5239 80935
rect 4985 80872 5010 80912
rect 5010 80872 5050 80912
rect 5050 80872 5071 80912
rect 5153 80872 5174 80912
rect 5174 80872 5214 80912
rect 5214 80872 5239 80912
rect 4985 80849 5071 80872
rect 5153 80849 5239 80872
rect 20105 80912 20191 80935
rect 20273 80912 20359 80935
rect 20105 80872 20130 80912
rect 20130 80872 20170 80912
rect 20170 80872 20191 80912
rect 20273 80872 20294 80912
rect 20294 80872 20334 80912
rect 20334 80872 20359 80912
rect 20105 80849 20191 80872
rect 20273 80849 20359 80872
rect 3745 80156 3831 80179
rect 3913 80156 3999 80179
rect 3745 80116 3770 80156
rect 3770 80116 3810 80156
rect 3810 80116 3831 80156
rect 3913 80116 3934 80156
rect 3934 80116 3974 80156
rect 3974 80116 3999 80156
rect 3745 80093 3831 80116
rect 3913 80093 3999 80116
rect 18865 80156 18951 80179
rect 19033 80156 19119 80179
rect 18865 80116 18890 80156
rect 18890 80116 18930 80156
rect 18930 80116 18951 80156
rect 19033 80116 19054 80156
rect 19054 80116 19094 80156
rect 19094 80116 19119 80156
rect 18865 80093 18951 80116
rect 19033 80093 19119 80116
rect 4985 79400 5071 79423
rect 5153 79400 5239 79423
rect 4985 79360 5010 79400
rect 5010 79360 5050 79400
rect 5050 79360 5071 79400
rect 5153 79360 5174 79400
rect 5174 79360 5214 79400
rect 5214 79360 5239 79400
rect 4985 79337 5071 79360
rect 5153 79337 5239 79360
rect 20105 79400 20191 79423
rect 20273 79400 20359 79423
rect 20105 79360 20130 79400
rect 20130 79360 20170 79400
rect 20170 79360 20191 79400
rect 20273 79360 20294 79400
rect 20294 79360 20334 79400
rect 20334 79360 20359 79400
rect 20105 79337 20191 79360
rect 20273 79337 20359 79360
rect 3745 78644 3831 78667
rect 3913 78644 3999 78667
rect 3745 78604 3770 78644
rect 3770 78604 3810 78644
rect 3810 78604 3831 78644
rect 3913 78604 3934 78644
rect 3934 78604 3974 78644
rect 3974 78604 3999 78644
rect 3745 78581 3831 78604
rect 3913 78581 3999 78604
rect 18865 78644 18951 78667
rect 19033 78644 19119 78667
rect 18865 78604 18890 78644
rect 18890 78604 18930 78644
rect 18930 78604 18951 78644
rect 19033 78604 19054 78644
rect 19054 78604 19094 78644
rect 19094 78604 19119 78644
rect 18865 78581 18951 78604
rect 19033 78581 19119 78604
rect 4985 77888 5071 77911
rect 5153 77888 5239 77911
rect 4985 77848 5010 77888
rect 5010 77848 5050 77888
rect 5050 77848 5071 77888
rect 5153 77848 5174 77888
rect 5174 77848 5214 77888
rect 5214 77848 5239 77888
rect 4985 77825 5071 77848
rect 5153 77825 5239 77848
rect 20105 77888 20191 77911
rect 20273 77888 20359 77911
rect 20105 77848 20130 77888
rect 20130 77848 20170 77888
rect 20170 77848 20191 77888
rect 20273 77848 20294 77888
rect 20294 77848 20334 77888
rect 20334 77848 20359 77888
rect 20105 77825 20191 77848
rect 20273 77825 20359 77848
rect 3745 77132 3831 77155
rect 3913 77132 3999 77155
rect 3745 77092 3770 77132
rect 3770 77092 3810 77132
rect 3810 77092 3831 77132
rect 3913 77092 3934 77132
rect 3934 77092 3974 77132
rect 3974 77092 3999 77132
rect 3745 77069 3831 77092
rect 3913 77069 3999 77092
rect 18865 77132 18951 77155
rect 19033 77132 19119 77155
rect 18865 77092 18890 77132
rect 18890 77092 18930 77132
rect 18930 77092 18951 77132
rect 19033 77092 19054 77132
rect 19054 77092 19094 77132
rect 19094 77092 19119 77132
rect 18865 77069 18951 77092
rect 19033 77069 19119 77092
rect 8493 76712 8579 76735
rect 8493 76672 8524 76712
rect 8524 76672 8564 76712
rect 8564 76672 8579 76712
rect 8493 76649 8579 76672
rect 9405 76649 9491 76735
rect 1197 76481 1283 76567
rect 4985 76376 5071 76399
rect 5153 76376 5239 76399
rect 4985 76336 5010 76376
rect 5010 76336 5050 76376
rect 5050 76336 5071 76376
rect 5153 76336 5174 76376
rect 5174 76336 5214 76376
rect 5214 76336 5239 76376
rect 4985 76313 5071 76336
rect 5153 76313 5239 76336
rect 20105 76376 20191 76399
rect 20273 76376 20359 76399
rect 20105 76336 20130 76376
rect 20130 76336 20170 76376
rect 20170 76336 20191 76376
rect 20273 76336 20294 76376
rect 20294 76336 20334 76376
rect 20334 76336 20359 76376
rect 20105 76313 20191 76336
rect 20273 76313 20359 76336
rect 3745 75620 3831 75643
rect 3913 75620 3999 75643
rect 3745 75580 3770 75620
rect 3770 75580 3810 75620
rect 3810 75580 3831 75620
rect 3913 75580 3934 75620
rect 3934 75580 3974 75620
rect 3974 75580 3999 75620
rect 3745 75557 3831 75580
rect 3913 75557 3999 75580
rect 18865 75620 18951 75643
rect 19033 75620 19119 75643
rect 18865 75580 18890 75620
rect 18890 75580 18930 75620
rect 18930 75580 18951 75620
rect 19033 75580 19054 75620
rect 19054 75580 19094 75620
rect 19094 75580 19119 75620
rect 18865 75557 18951 75580
rect 19033 75557 19119 75580
rect 4985 74864 5071 74887
rect 5153 74864 5239 74887
rect 4985 74824 5010 74864
rect 5010 74824 5050 74864
rect 5050 74824 5071 74864
rect 5153 74824 5174 74864
rect 5174 74824 5214 74864
rect 5214 74824 5239 74864
rect 4985 74801 5071 74824
rect 5153 74801 5239 74824
rect 20105 74864 20191 74887
rect 20273 74864 20359 74887
rect 20105 74824 20130 74864
rect 20130 74824 20170 74864
rect 20170 74824 20191 74864
rect 20273 74824 20294 74864
rect 20294 74824 20334 74864
rect 20334 74824 20359 74864
rect 20105 74801 20191 74824
rect 20273 74801 20359 74824
rect 3745 74108 3831 74131
rect 3913 74108 3999 74131
rect 3745 74068 3770 74108
rect 3770 74068 3810 74108
rect 3810 74068 3831 74108
rect 3913 74068 3934 74108
rect 3934 74068 3974 74108
rect 3974 74068 3999 74108
rect 3745 74045 3831 74068
rect 3913 74045 3999 74068
rect 18865 74108 18951 74131
rect 19033 74108 19119 74131
rect 18865 74068 18890 74108
rect 18890 74068 18930 74108
rect 18930 74068 18951 74108
rect 19033 74068 19054 74108
rect 19054 74068 19094 74108
rect 19094 74068 19119 74108
rect 18865 74045 18951 74068
rect 19033 74045 19119 74068
rect 4985 73352 5071 73375
rect 5153 73352 5239 73375
rect 4985 73312 5010 73352
rect 5010 73312 5050 73352
rect 5050 73312 5071 73352
rect 5153 73312 5174 73352
rect 5174 73312 5214 73352
rect 5214 73312 5239 73352
rect 4985 73289 5071 73312
rect 5153 73289 5239 73312
rect 20105 73352 20191 73375
rect 20273 73352 20359 73375
rect 20105 73312 20130 73352
rect 20130 73312 20170 73352
rect 20170 73312 20191 73352
rect 20273 73312 20294 73352
rect 20294 73312 20334 73352
rect 20334 73312 20359 73352
rect 20105 73289 20191 73312
rect 20273 73289 20359 73312
rect 3745 72596 3831 72619
rect 3913 72596 3999 72619
rect 3745 72556 3770 72596
rect 3770 72556 3810 72596
rect 3810 72556 3831 72596
rect 3913 72556 3934 72596
rect 3934 72556 3974 72596
rect 3974 72556 3999 72596
rect 3745 72533 3831 72556
rect 3913 72533 3999 72556
rect 18865 72596 18951 72619
rect 19033 72596 19119 72619
rect 18865 72556 18890 72596
rect 18890 72556 18930 72596
rect 18930 72556 18951 72596
rect 19033 72556 19054 72596
rect 19054 72556 19094 72596
rect 19094 72556 19119 72596
rect 18865 72533 18951 72556
rect 19033 72533 19119 72556
rect 4985 71840 5071 71863
rect 5153 71840 5239 71863
rect 4985 71800 5010 71840
rect 5010 71800 5050 71840
rect 5050 71800 5071 71840
rect 5153 71800 5174 71840
rect 5174 71800 5214 71840
rect 5214 71800 5239 71840
rect 4985 71777 5071 71800
rect 5153 71777 5239 71800
rect 20105 71840 20191 71863
rect 20273 71840 20359 71863
rect 20105 71800 20130 71840
rect 20130 71800 20170 71840
rect 20170 71800 20191 71840
rect 20273 71800 20294 71840
rect 20294 71800 20334 71840
rect 20334 71800 20359 71840
rect 20105 71777 20191 71800
rect 20273 71777 20359 71800
rect 3745 71084 3831 71107
rect 3913 71084 3999 71107
rect 3745 71044 3770 71084
rect 3770 71044 3810 71084
rect 3810 71044 3831 71084
rect 3913 71044 3934 71084
rect 3934 71044 3974 71084
rect 3974 71044 3999 71084
rect 3745 71021 3831 71044
rect 3913 71021 3999 71044
rect 18865 71084 18951 71107
rect 19033 71084 19119 71107
rect 18865 71044 18890 71084
rect 18890 71044 18930 71084
rect 18930 71044 18951 71084
rect 19033 71044 19054 71084
rect 19054 71044 19094 71084
rect 19094 71044 19119 71084
rect 18865 71021 18951 71044
rect 19033 71021 19119 71044
rect 4985 70328 5071 70351
rect 5153 70328 5239 70351
rect 4985 70288 5010 70328
rect 5010 70288 5050 70328
rect 5050 70288 5071 70328
rect 5153 70288 5174 70328
rect 5174 70288 5214 70328
rect 5214 70288 5239 70328
rect 4985 70265 5071 70288
rect 5153 70265 5239 70288
rect 20105 70328 20191 70351
rect 20273 70328 20359 70351
rect 20105 70288 20130 70328
rect 20130 70288 20170 70328
rect 20170 70288 20191 70328
rect 20273 70288 20294 70328
rect 20294 70288 20334 70328
rect 20334 70288 20359 70328
rect 20105 70265 20191 70288
rect 20273 70265 20359 70288
rect 3745 69572 3831 69595
rect 3913 69572 3999 69595
rect 3745 69532 3770 69572
rect 3770 69532 3810 69572
rect 3810 69532 3831 69572
rect 3913 69532 3934 69572
rect 3934 69532 3974 69572
rect 3974 69532 3999 69572
rect 3745 69509 3831 69532
rect 3913 69509 3999 69532
rect 18865 69572 18951 69595
rect 19033 69572 19119 69595
rect 18865 69532 18890 69572
rect 18890 69532 18930 69572
rect 18930 69532 18951 69572
rect 19033 69532 19054 69572
rect 19054 69532 19094 69572
rect 19094 69532 19119 69572
rect 18865 69509 18951 69532
rect 19033 69509 19119 69532
rect 4985 68816 5071 68839
rect 5153 68816 5239 68839
rect 4985 68776 5010 68816
rect 5010 68776 5050 68816
rect 5050 68776 5071 68816
rect 5153 68776 5174 68816
rect 5174 68776 5214 68816
rect 5214 68776 5239 68816
rect 4985 68753 5071 68776
rect 5153 68753 5239 68776
rect 20105 68816 20191 68839
rect 20273 68816 20359 68839
rect 20105 68776 20130 68816
rect 20130 68776 20170 68816
rect 20170 68776 20191 68816
rect 20273 68776 20294 68816
rect 20294 68776 20334 68816
rect 20334 68776 20359 68816
rect 20105 68753 20191 68776
rect 20273 68753 20359 68776
rect 3745 68060 3831 68083
rect 3913 68060 3999 68083
rect 18865 68060 18951 68083
rect 19033 68060 19119 68083
rect 3745 68020 3770 68060
rect 3770 68020 3810 68060
rect 3810 68020 3831 68060
rect 3913 68020 3934 68060
rect 3934 68020 3974 68060
rect 3974 68020 3999 68060
rect 18865 68020 18890 68060
rect 18890 68020 18930 68060
rect 18930 68020 18951 68060
rect 19033 68020 19054 68060
rect 19054 68020 19094 68060
rect 19094 68020 19119 68060
rect 3745 67997 3831 68020
rect 3913 67997 3999 68020
rect 18865 67997 18951 68020
rect 19033 67997 19119 68020
rect 4985 67304 5071 67327
rect 5153 67304 5239 67327
rect 4985 67264 5010 67304
rect 5010 67264 5050 67304
rect 5050 67264 5071 67304
rect 5153 67264 5174 67304
rect 5174 67264 5214 67304
rect 5214 67264 5239 67304
rect 4985 67241 5071 67264
rect 5153 67241 5239 67264
rect 20105 67304 20191 67327
rect 20273 67304 20359 67327
rect 20105 67264 20130 67304
rect 20130 67264 20170 67304
rect 20170 67264 20191 67304
rect 20273 67264 20294 67304
rect 20294 67264 20334 67304
rect 20334 67264 20359 67304
rect 20105 67241 20191 67264
rect 20273 67241 20359 67264
rect 3745 66548 3831 66571
rect 3913 66548 3999 66571
rect 3745 66508 3770 66548
rect 3770 66508 3810 66548
rect 3810 66508 3831 66548
rect 3913 66508 3934 66548
rect 3934 66508 3974 66548
rect 3974 66508 3999 66548
rect 3745 66485 3831 66508
rect 3913 66485 3999 66508
rect 18865 66548 18951 66571
rect 19033 66548 19119 66571
rect 18865 66508 18890 66548
rect 18890 66508 18930 66548
rect 18930 66508 18951 66548
rect 19033 66508 19054 66548
rect 19054 66508 19094 66548
rect 19094 66508 19119 66548
rect 18865 66485 18951 66508
rect 19033 66485 19119 66508
rect 4985 65792 5071 65815
rect 5153 65792 5239 65815
rect 4985 65752 5010 65792
rect 5010 65752 5050 65792
rect 5050 65752 5071 65792
rect 5153 65752 5174 65792
rect 5174 65752 5214 65792
rect 5214 65752 5239 65792
rect 4985 65729 5071 65752
rect 5153 65729 5239 65752
rect 20105 65792 20191 65815
rect 20273 65792 20359 65815
rect 20105 65752 20130 65792
rect 20130 65752 20170 65792
rect 20170 65752 20191 65792
rect 20273 65752 20294 65792
rect 20294 65752 20334 65792
rect 20334 65752 20359 65792
rect 20105 65729 20191 65752
rect 20273 65729 20359 65752
rect 3745 65036 3831 65059
rect 3913 65036 3999 65059
rect 3745 64996 3770 65036
rect 3770 64996 3810 65036
rect 3810 64996 3831 65036
rect 3913 64996 3934 65036
rect 3934 64996 3974 65036
rect 3974 64996 3999 65036
rect 3745 64973 3831 64996
rect 3913 64973 3999 64996
rect 18865 65036 18951 65059
rect 19033 65036 19119 65059
rect 18865 64996 18890 65036
rect 18890 64996 18930 65036
rect 18930 64996 18951 65036
rect 19033 64996 19054 65036
rect 19054 64996 19094 65036
rect 19094 64996 19119 65036
rect 18865 64973 18951 64996
rect 19033 64973 19119 64996
rect 4985 64280 5071 64303
rect 5153 64280 5239 64303
rect 4985 64240 5010 64280
rect 5010 64240 5050 64280
rect 5050 64240 5071 64280
rect 5153 64240 5174 64280
rect 5174 64240 5214 64280
rect 5214 64240 5239 64280
rect 4985 64217 5071 64240
rect 5153 64217 5239 64240
rect 20105 64280 20191 64303
rect 20273 64280 20359 64303
rect 20105 64240 20130 64280
rect 20130 64240 20170 64280
rect 20170 64240 20191 64280
rect 20273 64240 20294 64280
rect 20294 64240 20334 64280
rect 20334 64240 20359 64280
rect 20105 64217 20191 64240
rect 20273 64217 20359 64240
rect 3745 63524 3831 63547
rect 3913 63524 3999 63547
rect 3745 63484 3770 63524
rect 3770 63484 3810 63524
rect 3810 63484 3831 63524
rect 3913 63484 3934 63524
rect 3934 63484 3974 63524
rect 3974 63484 3999 63524
rect 3745 63461 3831 63484
rect 3913 63461 3999 63484
rect 18865 63524 18951 63547
rect 19033 63524 19119 63547
rect 18865 63484 18890 63524
rect 18890 63484 18930 63524
rect 18930 63484 18951 63524
rect 19033 63484 19054 63524
rect 19054 63484 19094 63524
rect 19094 63484 19119 63524
rect 18865 63461 18951 63484
rect 19033 63461 19119 63484
rect 4985 62768 5071 62791
rect 5153 62768 5239 62791
rect 4985 62728 5010 62768
rect 5010 62728 5050 62768
rect 5050 62728 5071 62768
rect 5153 62728 5174 62768
rect 5174 62728 5214 62768
rect 5214 62728 5239 62768
rect 4985 62705 5071 62728
rect 5153 62705 5239 62728
rect 20105 62768 20191 62791
rect 20273 62768 20359 62791
rect 20105 62728 20130 62768
rect 20130 62728 20170 62768
rect 20170 62728 20191 62768
rect 20273 62728 20294 62768
rect 20294 62728 20334 62768
rect 20334 62728 20359 62768
rect 20105 62705 20191 62728
rect 20273 62705 20359 62728
rect 3745 62012 3831 62035
rect 3913 62012 3999 62035
rect 3745 61972 3770 62012
rect 3770 61972 3810 62012
rect 3810 61972 3831 62012
rect 3913 61972 3934 62012
rect 3934 61972 3974 62012
rect 3974 61972 3999 62012
rect 3745 61949 3831 61972
rect 3913 61949 3999 61972
rect 18865 62012 18951 62035
rect 19033 62012 19119 62035
rect 18865 61972 18890 62012
rect 18890 61972 18930 62012
rect 18930 61972 18951 62012
rect 19033 61972 19054 62012
rect 19054 61972 19094 62012
rect 19094 61972 19119 62012
rect 18865 61949 18951 61972
rect 19033 61949 19119 61972
rect 4985 61256 5071 61279
rect 5153 61256 5239 61279
rect 4985 61216 5010 61256
rect 5010 61216 5050 61256
rect 5050 61216 5071 61256
rect 5153 61216 5174 61256
rect 5174 61216 5214 61256
rect 5214 61216 5239 61256
rect 4985 61193 5071 61216
rect 5153 61193 5239 61216
rect 20105 61256 20191 61279
rect 20273 61256 20359 61279
rect 20105 61216 20130 61256
rect 20130 61216 20170 61256
rect 20170 61216 20191 61256
rect 20273 61216 20294 61256
rect 20294 61216 20334 61256
rect 20334 61216 20359 61256
rect 20105 61193 20191 61216
rect 20273 61193 20359 61216
rect 3745 60500 3831 60523
rect 3913 60500 3999 60523
rect 3745 60460 3770 60500
rect 3770 60460 3810 60500
rect 3810 60460 3831 60500
rect 3913 60460 3934 60500
rect 3934 60460 3974 60500
rect 3974 60460 3999 60500
rect 3745 60437 3831 60460
rect 3913 60437 3999 60460
rect 18865 60500 18951 60523
rect 19033 60500 19119 60523
rect 18865 60460 18890 60500
rect 18890 60460 18930 60500
rect 18930 60460 18951 60500
rect 19033 60460 19054 60500
rect 19054 60460 19094 60500
rect 19094 60460 19119 60500
rect 18865 60437 18951 60460
rect 19033 60437 19119 60460
rect 4985 59744 5071 59767
rect 5153 59744 5239 59767
rect 4985 59704 5010 59744
rect 5010 59704 5050 59744
rect 5050 59704 5071 59744
rect 5153 59704 5174 59744
rect 5174 59704 5214 59744
rect 5214 59704 5239 59744
rect 4985 59681 5071 59704
rect 5153 59681 5239 59704
rect 20105 59744 20191 59767
rect 20273 59744 20359 59767
rect 20105 59704 20130 59744
rect 20130 59704 20170 59744
rect 20170 59704 20191 59744
rect 20273 59704 20294 59744
rect 20294 59704 20334 59744
rect 20334 59704 20359 59744
rect 20105 59681 20191 59704
rect 20273 59681 20359 59704
rect 3745 58988 3831 59011
rect 3913 58988 3999 59011
rect 3745 58948 3770 58988
rect 3770 58948 3810 58988
rect 3810 58948 3831 58988
rect 3913 58948 3934 58988
rect 3934 58948 3974 58988
rect 3974 58948 3999 58988
rect 3745 58925 3831 58948
rect 3913 58925 3999 58948
rect 18865 58988 18951 59011
rect 19033 58988 19119 59011
rect 18865 58948 18890 58988
rect 18890 58948 18930 58988
rect 18930 58948 18951 58988
rect 19033 58948 19054 58988
rect 19054 58948 19094 58988
rect 19094 58948 19119 58988
rect 18865 58925 18951 58948
rect 19033 58925 19119 58948
rect 4985 58232 5071 58255
rect 5153 58232 5239 58255
rect 4985 58192 5010 58232
rect 5010 58192 5050 58232
rect 5050 58192 5071 58232
rect 5153 58192 5174 58232
rect 5174 58192 5214 58232
rect 5214 58192 5239 58232
rect 4985 58169 5071 58192
rect 5153 58169 5239 58192
rect 20105 58232 20191 58255
rect 20273 58232 20359 58255
rect 20105 58192 20130 58232
rect 20130 58192 20170 58232
rect 20170 58192 20191 58232
rect 20273 58192 20294 58232
rect 20294 58192 20334 58232
rect 20334 58192 20359 58232
rect 20105 58169 20191 58192
rect 20273 58169 20359 58192
rect 3745 57476 3831 57499
rect 3913 57476 3999 57499
rect 3745 57436 3770 57476
rect 3770 57436 3810 57476
rect 3810 57436 3831 57476
rect 3913 57436 3934 57476
rect 3934 57436 3974 57476
rect 3974 57436 3999 57476
rect 3745 57413 3831 57436
rect 3913 57413 3999 57436
rect 18865 57476 18951 57499
rect 19033 57476 19119 57499
rect 18865 57436 18890 57476
rect 18890 57436 18930 57476
rect 18930 57436 18951 57476
rect 19033 57436 19054 57476
rect 19054 57436 19094 57476
rect 19094 57436 19119 57476
rect 18865 57413 18951 57436
rect 19033 57413 19119 57436
rect 4985 56720 5071 56743
rect 5153 56720 5239 56743
rect 4985 56680 5010 56720
rect 5010 56680 5050 56720
rect 5050 56680 5071 56720
rect 5153 56680 5174 56720
rect 5174 56680 5214 56720
rect 5214 56680 5239 56720
rect 4985 56657 5071 56680
rect 5153 56657 5239 56680
rect 20105 56720 20191 56743
rect 20273 56720 20359 56743
rect 20105 56680 20130 56720
rect 20130 56680 20170 56720
rect 20170 56680 20191 56720
rect 20273 56680 20294 56720
rect 20294 56680 20334 56720
rect 20334 56680 20359 56720
rect 20105 56657 20191 56680
rect 20273 56657 20359 56680
rect 3745 55964 3831 55987
rect 3913 55964 3999 55987
rect 3745 55924 3770 55964
rect 3770 55924 3810 55964
rect 3810 55924 3831 55964
rect 3913 55924 3934 55964
rect 3934 55924 3974 55964
rect 3974 55924 3999 55964
rect 3745 55901 3831 55924
rect 3913 55901 3999 55924
rect 18865 55964 18951 55987
rect 19033 55964 19119 55987
rect 18865 55924 18890 55964
rect 18890 55924 18930 55964
rect 18930 55924 18951 55964
rect 19033 55924 19054 55964
rect 19054 55924 19094 55964
rect 19094 55924 19119 55964
rect 18865 55901 18951 55924
rect 19033 55901 19119 55924
rect 4985 55208 5071 55231
rect 5153 55208 5239 55231
rect 4985 55168 5010 55208
rect 5010 55168 5050 55208
rect 5050 55168 5071 55208
rect 5153 55168 5174 55208
rect 5174 55168 5214 55208
rect 5214 55168 5239 55208
rect 4985 55145 5071 55168
rect 5153 55145 5239 55168
rect 20105 55208 20191 55231
rect 20273 55208 20359 55231
rect 20105 55168 20130 55208
rect 20130 55168 20170 55208
rect 20170 55168 20191 55208
rect 20273 55168 20294 55208
rect 20294 55168 20334 55208
rect 20334 55168 20359 55208
rect 20105 55145 20191 55168
rect 20273 55145 20359 55168
rect 3745 54452 3831 54475
rect 3913 54452 3999 54475
rect 3745 54412 3770 54452
rect 3770 54412 3810 54452
rect 3810 54412 3831 54452
rect 3913 54412 3934 54452
rect 3934 54412 3974 54452
rect 3974 54412 3999 54452
rect 3745 54389 3831 54412
rect 3913 54389 3999 54412
rect 18865 54452 18951 54475
rect 19033 54452 19119 54475
rect 18865 54412 18890 54452
rect 18890 54412 18930 54452
rect 18930 54412 18951 54452
rect 19033 54412 19054 54452
rect 19054 54412 19094 54452
rect 19094 54412 19119 54452
rect 18865 54389 18951 54412
rect 19033 54389 19119 54412
rect 4985 53696 5071 53719
rect 5153 53696 5239 53719
rect 4985 53656 5010 53696
rect 5010 53656 5050 53696
rect 5050 53656 5071 53696
rect 5153 53656 5174 53696
rect 5174 53656 5214 53696
rect 5214 53656 5239 53696
rect 4985 53633 5071 53656
rect 5153 53633 5239 53656
rect 20105 53696 20191 53719
rect 20273 53696 20359 53719
rect 20105 53656 20130 53696
rect 20130 53656 20170 53696
rect 20170 53656 20191 53696
rect 20273 53656 20294 53696
rect 20294 53656 20334 53696
rect 20334 53656 20359 53696
rect 20105 53633 20191 53656
rect 20273 53633 20359 53656
rect 3745 52940 3831 52963
rect 3913 52940 3999 52963
rect 3745 52900 3770 52940
rect 3770 52900 3810 52940
rect 3810 52900 3831 52940
rect 3913 52900 3934 52940
rect 3934 52900 3974 52940
rect 3974 52900 3999 52940
rect 3745 52877 3831 52900
rect 3913 52877 3999 52900
rect 18865 52940 18951 52963
rect 19033 52940 19119 52963
rect 18865 52900 18890 52940
rect 18890 52900 18930 52940
rect 18930 52900 18951 52940
rect 19033 52900 19054 52940
rect 19054 52900 19094 52940
rect 19094 52900 19119 52940
rect 18865 52877 18951 52900
rect 19033 52877 19119 52900
rect 4985 52184 5071 52207
rect 5153 52184 5239 52207
rect 4985 52144 5010 52184
rect 5010 52144 5050 52184
rect 5050 52144 5071 52184
rect 5153 52144 5174 52184
rect 5174 52144 5214 52184
rect 5214 52144 5239 52184
rect 4985 52121 5071 52144
rect 5153 52121 5239 52144
rect 20105 52184 20191 52207
rect 20273 52184 20359 52207
rect 20105 52144 20130 52184
rect 20130 52144 20170 52184
rect 20170 52144 20191 52184
rect 20273 52144 20294 52184
rect 20294 52144 20334 52184
rect 20334 52144 20359 52184
rect 20105 52121 20191 52144
rect 20273 52121 20359 52144
rect 3745 51428 3831 51451
rect 3913 51428 3999 51451
rect 3745 51388 3770 51428
rect 3770 51388 3810 51428
rect 3810 51388 3831 51428
rect 3913 51388 3934 51428
rect 3934 51388 3974 51428
rect 3974 51388 3999 51428
rect 3745 51365 3831 51388
rect 3913 51365 3999 51388
rect 18865 51428 18951 51451
rect 19033 51428 19119 51451
rect 18865 51388 18890 51428
rect 18890 51388 18930 51428
rect 18930 51388 18951 51428
rect 19033 51388 19054 51428
rect 19054 51388 19094 51428
rect 19094 51388 19119 51428
rect 18865 51365 18951 51388
rect 19033 51365 19119 51388
rect 4985 50672 5071 50695
rect 5153 50672 5239 50695
rect 4985 50632 5010 50672
rect 5010 50632 5050 50672
rect 5050 50632 5071 50672
rect 5153 50632 5174 50672
rect 5174 50632 5214 50672
rect 5214 50632 5239 50672
rect 4985 50609 5071 50632
rect 5153 50609 5239 50632
rect 20105 50672 20191 50695
rect 20273 50672 20359 50695
rect 20105 50632 20130 50672
rect 20130 50632 20170 50672
rect 20170 50632 20191 50672
rect 20273 50632 20294 50672
rect 20294 50632 20334 50672
rect 20334 50632 20359 50672
rect 20105 50609 20191 50632
rect 20273 50609 20359 50632
rect 3745 49916 3831 49939
rect 3913 49916 3999 49939
rect 3745 49876 3770 49916
rect 3770 49876 3810 49916
rect 3810 49876 3831 49916
rect 3913 49876 3934 49916
rect 3934 49876 3974 49916
rect 3974 49876 3999 49916
rect 3745 49853 3831 49876
rect 3913 49853 3999 49876
rect 18865 49916 18951 49939
rect 19033 49916 19119 49939
rect 18865 49876 18890 49916
rect 18890 49876 18930 49916
rect 18930 49876 18951 49916
rect 19033 49876 19054 49916
rect 19054 49876 19094 49916
rect 19094 49876 19119 49916
rect 18865 49853 18951 49876
rect 19033 49853 19119 49876
rect 4985 49160 5071 49183
rect 5153 49160 5239 49183
rect 4985 49120 5010 49160
rect 5010 49120 5050 49160
rect 5050 49120 5071 49160
rect 5153 49120 5174 49160
rect 5174 49120 5214 49160
rect 5214 49120 5239 49160
rect 4985 49097 5071 49120
rect 5153 49097 5239 49120
rect 20105 49160 20191 49183
rect 20273 49160 20359 49183
rect 20105 49120 20130 49160
rect 20130 49120 20170 49160
rect 20170 49120 20191 49160
rect 20273 49120 20294 49160
rect 20294 49120 20334 49160
rect 20334 49120 20359 49160
rect 20105 49097 20191 49120
rect 20273 49097 20359 49120
rect 3745 48404 3831 48427
rect 3913 48404 3999 48427
rect 3745 48364 3770 48404
rect 3770 48364 3810 48404
rect 3810 48364 3831 48404
rect 3913 48364 3934 48404
rect 3934 48364 3974 48404
rect 3974 48364 3999 48404
rect 3745 48341 3831 48364
rect 3913 48341 3999 48364
rect 18865 48404 18951 48427
rect 19033 48404 19119 48427
rect 18865 48364 18890 48404
rect 18890 48364 18930 48404
rect 18930 48364 18951 48404
rect 19033 48364 19054 48404
rect 19054 48364 19094 48404
rect 19094 48364 19119 48404
rect 18865 48341 18951 48364
rect 19033 48341 19119 48364
rect 2109 47837 2195 47923
rect 4985 47648 5071 47671
rect 5153 47648 5239 47671
rect 4985 47608 5010 47648
rect 5010 47608 5050 47648
rect 5050 47608 5071 47648
rect 5153 47608 5174 47648
rect 5174 47608 5214 47648
rect 5214 47608 5239 47648
rect 4985 47585 5071 47608
rect 5153 47585 5239 47608
rect 20105 47648 20191 47671
rect 20273 47648 20359 47671
rect 20105 47608 20130 47648
rect 20130 47608 20170 47648
rect 20170 47608 20191 47648
rect 20273 47608 20294 47648
rect 20294 47608 20334 47648
rect 20334 47608 20359 47648
rect 20105 47585 20191 47608
rect 20273 47585 20359 47608
rect 3745 46892 3831 46915
rect 3913 46892 3999 46915
rect 3745 46852 3770 46892
rect 3770 46852 3810 46892
rect 3810 46852 3831 46892
rect 3913 46852 3934 46892
rect 3934 46852 3974 46892
rect 3974 46852 3999 46892
rect 3745 46829 3831 46852
rect 3913 46829 3999 46852
rect 18865 46892 18951 46915
rect 19033 46892 19119 46915
rect 18865 46852 18890 46892
rect 18890 46852 18930 46892
rect 18930 46852 18951 46892
rect 19033 46852 19054 46892
rect 19054 46852 19094 46892
rect 19094 46852 19119 46892
rect 18865 46829 18951 46852
rect 19033 46829 19119 46852
rect 4985 46136 5071 46159
rect 5153 46136 5239 46159
rect 4985 46096 5010 46136
rect 5010 46096 5050 46136
rect 5050 46096 5071 46136
rect 5153 46096 5174 46136
rect 5174 46096 5214 46136
rect 5214 46096 5239 46136
rect 4985 46073 5071 46096
rect 5153 46073 5239 46096
rect 20105 46136 20191 46159
rect 20273 46136 20359 46159
rect 20105 46096 20130 46136
rect 20130 46096 20170 46136
rect 20170 46096 20191 46136
rect 20273 46096 20294 46136
rect 20294 46096 20334 46136
rect 20334 46096 20359 46136
rect 20105 46073 20191 46096
rect 20273 46073 20359 46096
rect 2109 45905 2195 45991
rect 3745 45380 3831 45403
rect 3913 45380 3999 45403
rect 3745 45340 3770 45380
rect 3770 45340 3810 45380
rect 3810 45340 3831 45380
rect 3913 45340 3934 45380
rect 3934 45340 3974 45380
rect 3974 45340 3999 45380
rect 3745 45317 3831 45340
rect 3913 45317 3999 45340
rect 18865 45380 18951 45403
rect 19033 45380 19119 45403
rect 18865 45340 18890 45380
rect 18890 45340 18930 45380
rect 18930 45340 18951 45380
rect 19033 45340 19054 45380
rect 19054 45340 19094 45380
rect 19094 45340 19119 45380
rect 18865 45317 18951 45340
rect 19033 45317 19119 45340
rect 4985 44624 5071 44647
rect 5153 44624 5239 44647
rect 4985 44584 5010 44624
rect 5010 44584 5050 44624
rect 5050 44584 5071 44624
rect 5153 44584 5174 44624
rect 5174 44584 5214 44624
rect 5214 44584 5239 44624
rect 4985 44561 5071 44584
rect 5153 44561 5239 44584
rect 20105 44624 20191 44647
rect 20273 44624 20359 44647
rect 20105 44584 20130 44624
rect 20130 44584 20170 44624
rect 20170 44584 20191 44624
rect 20273 44584 20294 44624
rect 20294 44584 20334 44624
rect 20334 44584 20359 44624
rect 20105 44561 20191 44584
rect 20273 44561 20359 44584
rect 3745 43868 3831 43891
rect 3913 43868 3999 43891
rect 3745 43828 3770 43868
rect 3770 43828 3810 43868
rect 3810 43828 3831 43868
rect 3913 43828 3934 43868
rect 3934 43828 3974 43868
rect 3974 43828 3999 43868
rect 3745 43805 3831 43828
rect 3913 43805 3999 43828
rect 18865 43868 18951 43891
rect 19033 43868 19119 43891
rect 18865 43828 18890 43868
rect 18890 43828 18930 43868
rect 18930 43828 18951 43868
rect 19033 43828 19054 43868
rect 19054 43828 19094 43868
rect 19094 43828 19119 43868
rect 18865 43805 18951 43828
rect 19033 43805 19119 43828
rect 4985 43112 5071 43135
rect 5153 43112 5239 43135
rect 4985 43072 5010 43112
rect 5010 43072 5050 43112
rect 5050 43072 5071 43112
rect 5153 43072 5174 43112
rect 5174 43072 5214 43112
rect 5214 43072 5239 43112
rect 4985 43049 5071 43072
rect 5153 43049 5239 43072
rect 20105 43112 20191 43135
rect 20273 43112 20359 43135
rect 20105 43072 20130 43112
rect 20130 43072 20170 43112
rect 20170 43072 20191 43112
rect 20273 43072 20294 43112
rect 20294 43072 20334 43112
rect 20334 43072 20359 43112
rect 20105 43049 20191 43072
rect 20273 43049 20359 43072
rect 3745 42356 3831 42379
rect 3913 42356 3999 42379
rect 3745 42316 3770 42356
rect 3770 42316 3810 42356
rect 3810 42316 3831 42356
rect 3913 42316 3934 42356
rect 3934 42316 3974 42356
rect 3974 42316 3999 42356
rect 3745 42293 3831 42316
rect 3913 42293 3999 42316
rect 18865 42356 18951 42379
rect 19033 42356 19119 42379
rect 18865 42316 18890 42356
rect 18890 42316 18930 42356
rect 18930 42316 18951 42356
rect 19033 42316 19054 42356
rect 19054 42316 19094 42356
rect 19094 42316 19119 42356
rect 18865 42293 18951 42316
rect 19033 42293 19119 42316
rect 10317 41873 10403 41959
rect 4985 41600 5071 41623
rect 5153 41600 5239 41623
rect 4985 41560 5010 41600
rect 5010 41560 5050 41600
rect 5050 41560 5071 41600
rect 5153 41560 5174 41600
rect 5174 41560 5214 41600
rect 5214 41560 5239 41600
rect 4985 41537 5071 41560
rect 5153 41537 5239 41560
rect 20105 41600 20191 41623
rect 20273 41600 20359 41623
rect 20105 41560 20130 41600
rect 20130 41560 20170 41600
rect 20170 41560 20191 41600
rect 20273 41560 20294 41600
rect 20294 41560 20334 41600
rect 20334 41560 20359 41600
rect 20105 41537 20191 41560
rect 20273 41537 20359 41560
rect 3745 40844 3831 40867
rect 3913 40844 3999 40867
rect 3745 40804 3770 40844
rect 3770 40804 3810 40844
rect 3810 40804 3831 40844
rect 3913 40804 3934 40844
rect 3934 40804 3974 40844
rect 3974 40804 3999 40844
rect 3745 40781 3831 40804
rect 3913 40781 3999 40804
rect 18865 40844 18951 40867
rect 19033 40844 19119 40867
rect 18865 40804 18890 40844
rect 18890 40804 18930 40844
rect 18930 40804 18951 40844
rect 19033 40804 19054 40844
rect 19054 40804 19094 40844
rect 19094 40804 19119 40844
rect 18865 40781 18951 40804
rect 19033 40781 19119 40804
rect 4985 40088 5071 40111
rect 5153 40088 5239 40111
rect 4985 40048 5010 40088
rect 5010 40048 5050 40088
rect 5050 40048 5071 40088
rect 5153 40048 5174 40088
rect 5174 40048 5214 40088
rect 5214 40048 5239 40088
rect 4985 40025 5071 40048
rect 5153 40025 5239 40048
rect 20105 40088 20191 40111
rect 20273 40088 20359 40111
rect 20105 40048 20130 40088
rect 20130 40048 20170 40088
rect 20170 40048 20191 40088
rect 20273 40048 20294 40088
rect 20294 40048 20334 40088
rect 20334 40048 20359 40088
rect 20105 40025 20191 40048
rect 20273 40025 20359 40048
rect 3745 39332 3831 39355
rect 3913 39332 3999 39355
rect 3745 39292 3770 39332
rect 3770 39292 3810 39332
rect 3810 39292 3831 39332
rect 3913 39292 3934 39332
rect 3934 39292 3974 39332
rect 3974 39292 3999 39332
rect 3745 39269 3831 39292
rect 3913 39269 3999 39292
rect 18865 39332 18951 39355
rect 19033 39332 19119 39355
rect 18865 39292 18890 39332
rect 18890 39292 18930 39332
rect 18930 39292 18951 39332
rect 19033 39292 19054 39332
rect 19054 39292 19094 39332
rect 19094 39292 19119 39332
rect 18865 39269 18951 39292
rect 19033 39269 19119 39292
rect 4985 38576 5071 38599
rect 5153 38576 5239 38599
rect 4985 38536 5010 38576
rect 5010 38536 5050 38576
rect 5050 38536 5071 38576
rect 5153 38536 5174 38576
rect 5174 38536 5214 38576
rect 5214 38536 5239 38576
rect 4985 38513 5071 38536
rect 5153 38513 5239 38536
rect 20105 38576 20191 38599
rect 20273 38576 20359 38599
rect 20105 38536 20130 38576
rect 20130 38536 20170 38576
rect 20170 38536 20191 38576
rect 20273 38536 20294 38576
rect 20294 38536 20334 38576
rect 20334 38536 20359 38576
rect 20105 38513 20191 38536
rect 20273 38513 20359 38536
rect 3745 37820 3831 37843
rect 3913 37820 3999 37843
rect 3745 37780 3770 37820
rect 3770 37780 3810 37820
rect 3810 37780 3831 37820
rect 3913 37780 3934 37820
rect 3934 37780 3974 37820
rect 3974 37780 3999 37820
rect 3745 37757 3831 37780
rect 3913 37757 3999 37780
rect 18865 37820 18951 37843
rect 19033 37820 19119 37843
rect 18865 37780 18890 37820
rect 18890 37780 18930 37820
rect 18930 37780 18951 37820
rect 19033 37780 19054 37820
rect 19054 37780 19094 37820
rect 19094 37780 19119 37820
rect 18865 37757 18951 37780
rect 19033 37757 19119 37780
rect 4985 37064 5071 37087
rect 5153 37064 5239 37087
rect 4985 37024 5010 37064
rect 5010 37024 5050 37064
rect 5050 37024 5071 37064
rect 5153 37024 5174 37064
rect 5174 37024 5214 37064
rect 5214 37024 5239 37064
rect 4985 37001 5071 37024
rect 5153 37001 5239 37024
rect 20105 37064 20191 37087
rect 20273 37064 20359 37087
rect 20105 37024 20130 37064
rect 20130 37024 20170 37064
rect 20170 37024 20191 37064
rect 20273 37024 20294 37064
rect 20294 37024 20334 37064
rect 20334 37024 20359 37064
rect 20105 37001 20191 37024
rect 20273 37001 20359 37024
rect 3745 36308 3831 36331
rect 3913 36308 3999 36331
rect 3745 36268 3770 36308
rect 3770 36268 3810 36308
rect 3810 36268 3831 36308
rect 3913 36268 3934 36308
rect 3934 36268 3974 36308
rect 3974 36268 3999 36308
rect 3745 36245 3831 36268
rect 3913 36245 3999 36268
rect 18865 36308 18951 36331
rect 19033 36308 19119 36331
rect 18865 36268 18890 36308
rect 18890 36268 18930 36308
rect 18930 36268 18951 36308
rect 19033 36268 19054 36308
rect 19054 36268 19094 36308
rect 19094 36268 19119 36308
rect 18865 36245 18951 36268
rect 19033 36245 19119 36268
rect 4985 35552 5071 35575
rect 5153 35552 5239 35575
rect 4985 35512 5010 35552
rect 5010 35512 5050 35552
rect 5050 35512 5071 35552
rect 5153 35512 5174 35552
rect 5174 35512 5214 35552
rect 5214 35512 5239 35552
rect 4985 35489 5071 35512
rect 5153 35489 5239 35512
rect 20105 35552 20191 35575
rect 20273 35552 20359 35575
rect 20105 35512 20130 35552
rect 20130 35512 20170 35552
rect 20170 35512 20191 35552
rect 20273 35512 20294 35552
rect 20294 35512 20334 35552
rect 20334 35512 20359 35552
rect 20105 35489 20191 35512
rect 20273 35489 20359 35512
rect 3745 34796 3831 34819
rect 3913 34796 3999 34819
rect 3745 34756 3770 34796
rect 3770 34756 3810 34796
rect 3810 34756 3831 34796
rect 3913 34756 3934 34796
rect 3934 34756 3974 34796
rect 3974 34756 3999 34796
rect 3745 34733 3831 34756
rect 3913 34733 3999 34756
rect 18865 34796 18951 34819
rect 19033 34796 19119 34819
rect 18865 34756 18890 34796
rect 18890 34756 18930 34796
rect 18930 34756 18951 34796
rect 19033 34756 19054 34796
rect 19054 34756 19094 34796
rect 19094 34756 19119 34796
rect 18865 34733 18951 34756
rect 19033 34733 19119 34756
rect 1197 34313 1283 34399
rect 4985 34040 5071 34063
rect 5153 34040 5239 34063
rect 4985 34000 5010 34040
rect 5010 34000 5050 34040
rect 5050 34000 5071 34040
rect 5153 34000 5174 34040
rect 5174 34000 5214 34040
rect 5214 34000 5239 34040
rect 4985 33977 5071 34000
rect 5153 33977 5239 34000
rect 20105 34040 20191 34063
rect 20273 34040 20359 34063
rect 20105 34000 20130 34040
rect 20130 34000 20170 34040
rect 20170 34000 20191 34040
rect 20273 34000 20294 34040
rect 20294 34000 20334 34040
rect 20334 34000 20359 34040
rect 20105 33977 20191 34000
rect 20273 33977 20359 34000
rect 3745 33284 3831 33307
rect 3913 33284 3999 33307
rect 3745 33244 3770 33284
rect 3770 33244 3810 33284
rect 3810 33244 3831 33284
rect 3913 33244 3934 33284
rect 3934 33244 3974 33284
rect 3974 33244 3999 33284
rect 3745 33221 3831 33244
rect 3913 33221 3999 33244
rect 18865 33284 18951 33307
rect 19033 33284 19119 33307
rect 18865 33244 18890 33284
rect 18890 33244 18930 33284
rect 18930 33244 18951 33284
rect 19033 33244 19054 33284
rect 19054 33244 19094 33284
rect 19094 33244 19119 33284
rect 18865 33221 18951 33244
rect 19033 33221 19119 33244
rect 4985 32528 5071 32551
rect 5153 32528 5239 32551
rect 4985 32488 5010 32528
rect 5010 32488 5050 32528
rect 5050 32488 5071 32528
rect 5153 32488 5174 32528
rect 5174 32488 5214 32528
rect 5214 32488 5239 32528
rect 4985 32465 5071 32488
rect 5153 32465 5239 32488
rect 20105 32528 20191 32551
rect 20273 32528 20359 32551
rect 20105 32488 20130 32528
rect 20130 32488 20170 32528
rect 20170 32488 20191 32528
rect 20273 32488 20294 32528
rect 20294 32488 20334 32528
rect 20334 32488 20359 32528
rect 20105 32465 20191 32488
rect 20273 32465 20359 32488
rect 3745 31772 3831 31795
rect 3913 31772 3999 31795
rect 3745 31732 3770 31772
rect 3770 31732 3810 31772
rect 3810 31732 3831 31772
rect 3913 31732 3934 31772
rect 3934 31732 3974 31772
rect 3974 31732 3999 31772
rect 3745 31709 3831 31732
rect 3913 31709 3999 31732
rect 18865 31772 18951 31795
rect 19033 31772 19119 31795
rect 18865 31732 18890 31772
rect 18890 31732 18930 31772
rect 18930 31732 18951 31772
rect 19033 31732 19054 31772
rect 19054 31732 19094 31772
rect 19094 31732 19119 31772
rect 18865 31709 18951 31732
rect 19033 31709 19119 31732
rect 4985 31016 5071 31039
rect 5153 31016 5239 31039
rect 4985 30976 5010 31016
rect 5010 30976 5050 31016
rect 5050 30976 5071 31016
rect 5153 30976 5174 31016
rect 5174 30976 5214 31016
rect 5214 30976 5239 31016
rect 4985 30953 5071 30976
rect 5153 30953 5239 30976
rect 20105 31016 20191 31039
rect 20273 31016 20359 31039
rect 20105 30976 20130 31016
rect 20130 30976 20170 31016
rect 20170 30976 20191 31016
rect 20273 30976 20294 31016
rect 20294 30976 20334 31016
rect 20334 30976 20359 31016
rect 20105 30953 20191 30976
rect 20273 30953 20359 30976
rect 3745 30260 3831 30283
rect 3913 30260 3999 30283
rect 3745 30220 3770 30260
rect 3770 30220 3810 30260
rect 3810 30220 3831 30260
rect 3913 30220 3934 30260
rect 3934 30220 3974 30260
rect 3974 30220 3999 30260
rect 3745 30197 3831 30220
rect 3913 30197 3999 30220
rect 18865 30260 18951 30283
rect 19033 30260 19119 30283
rect 18865 30220 18890 30260
rect 18890 30220 18930 30260
rect 18930 30220 18951 30260
rect 19033 30220 19054 30260
rect 19054 30220 19094 30260
rect 19094 30220 19119 30260
rect 18865 30197 18951 30220
rect 19033 30197 19119 30220
rect 4985 29504 5071 29527
rect 5153 29504 5239 29527
rect 4985 29464 5010 29504
rect 5010 29464 5050 29504
rect 5050 29464 5071 29504
rect 5153 29464 5174 29504
rect 5174 29464 5214 29504
rect 5214 29464 5239 29504
rect 4985 29441 5071 29464
rect 5153 29441 5239 29464
rect 20105 29504 20191 29527
rect 20273 29504 20359 29527
rect 20105 29464 20130 29504
rect 20130 29464 20170 29504
rect 20170 29464 20191 29504
rect 20273 29464 20294 29504
rect 20294 29464 20334 29504
rect 20334 29464 20359 29504
rect 20105 29441 20191 29464
rect 20273 29441 20359 29464
rect 3745 28748 3831 28771
rect 3913 28748 3999 28771
rect 3745 28708 3770 28748
rect 3770 28708 3810 28748
rect 3810 28708 3831 28748
rect 3913 28708 3934 28748
rect 3934 28708 3974 28748
rect 3974 28708 3999 28748
rect 3745 28685 3831 28708
rect 3913 28685 3999 28708
rect 18865 28748 18951 28771
rect 19033 28748 19119 28771
rect 18865 28708 18890 28748
rect 18890 28708 18930 28748
rect 18930 28708 18951 28748
rect 19033 28708 19054 28748
rect 19054 28708 19094 28748
rect 19094 28708 19119 28748
rect 18865 28685 18951 28708
rect 19033 28685 19119 28708
rect 4985 27992 5071 28015
rect 5153 27992 5239 28015
rect 4985 27952 5010 27992
rect 5010 27952 5050 27992
rect 5050 27952 5071 27992
rect 5153 27952 5174 27992
rect 5174 27952 5214 27992
rect 5214 27952 5239 27992
rect 4985 27929 5071 27952
rect 5153 27929 5239 27952
rect 20105 27992 20191 28015
rect 20273 27992 20359 28015
rect 20105 27952 20130 27992
rect 20130 27952 20170 27992
rect 20170 27952 20191 27992
rect 20273 27952 20294 27992
rect 20294 27952 20334 27992
rect 20334 27952 20359 27992
rect 20105 27929 20191 27952
rect 20273 27929 20359 27952
rect 3745 27236 3831 27259
rect 3913 27236 3999 27259
rect 3745 27196 3770 27236
rect 3770 27196 3810 27236
rect 3810 27196 3831 27236
rect 3913 27196 3934 27236
rect 3934 27196 3974 27236
rect 3974 27196 3999 27236
rect 3745 27173 3831 27196
rect 3913 27173 3999 27196
rect 18865 27236 18951 27259
rect 19033 27236 19119 27259
rect 18865 27196 18890 27236
rect 18890 27196 18930 27236
rect 18930 27196 18951 27236
rect 19033 27196 19054 27236
rect 19054 27196 19094 27236
rect 19094 27196 19119 27236
rect 18865 27173 18951 27196
rect 19033 27173 19119 27196
rect 4985 26480 5071 26503
rect 5153 26480 5239 26503
rect 4985 26440 5010 26480
rect 5010 26440 5050 26480
rect 5050 26440 5071 26480
rect 5153 26440 5174 26480
rect 5174 26440 5214 26480
rect 5214 26440 5239 26480
rect 4985 26417 5071 26440
rect 5153 26417 5239 26440
rect 20105 26480 20191 26503
rect 20273 26480 20359 26503
rect 20105 26440 20130 26480
rect 20130 26440 20170 26480
rect 20170 26440 20191 26480
rect 20273 26440 20294 26480
rect 20294 26440 20334 26480
rect 20334 26440 20359 26480
rect 20105 26417 20191 26440
rect 20273 26417 20359 26440
rect 3745 25724 3831 25747
rect 3913 25724 3999 25747
rect 3745 25684 3770 25724
rect 3770 25684 3810 25724
rect 3810 25684 3831 25724
rect 3913 25684 3934 25724
rect 3934 25684 3974 25724
rect 3974 25684 3999 25724
rect 3745 25661 3831 25684
rect 3913 25661 3999 25684
rect 18865 25724 18951 25747
rect 19033 25724 19119 25747
rect 18865 25684 18890 25724
rect 18890 25684 18930 25724
rect 18930 25684 18951 25724
rect 19033 25684 19054 25724
rect 19054 25684 19094 25724
rect 19094 25684 19119 25724
rect 18865 25661 18951 25684
rect 19033 25661 19119 25684
rect 4985 24968 5071 24991
rect 5153 24968 5239 24991
rect 4985 24928 5010 24968
rect 5010 24928 5050 24968
rect 5050 24928 5071 24968
rect 5153 24928 5174 24968
rect 5174 24928 5214 24968
rect 5214 24928 5239 24968
rect 4985 24905 5071 24928
rect 5153 24905 5239 24928
rect 20105 24968 20191 24991
rect 20273 24968 20359 24991
rect 20105 24928 20130 24968
rect 20130 24928 20170 24968
rect 20170 24928 20191 24968
rect 20273 24928 20294 24968
rect 20294 24928 20334 24968
rect 20334 24928 20359 24968
rect 20105 24905 20191 24928
rect 20273 24905 20359 24928
rect 16245 24569 16331 24655
rect 3745 24212 3831 24235
rect 3913 24212 3999 24235
rect 3745 24172 3770 24212
rect 3770 24172 3810 24212
rect 3810 24172 3831 24212
rect 3913 24172 3934 24212
rect 3934 24172 3974 24212
rect 3974 24172 3999 24212
rect 3745 24149 3831 24172
rect 3913 24149 3999 24172
rect 18865 24212 18951 24235
rect 19033 24212 19119 24235
rect 18865 24172 18890 24212
rect 18890 24172 18930 24212
rect 18930 24172 18951 24212
rect 19033 24172 19054 24212
rect 19054 24172 19094 24212
rect 19094 24172 19119 24212
rect 18865 24149 18951 24172
rect 19033 24149 19119 24172
rect 4985 23456 5071 23479
rect 5153 23456 5239 23479
rect 4985 23416 5010 23456
rect 5010 23416 5050 23456
rect 5050 23416 5071 23456
rect 5153 23416 5174 23456
rect 5174 23416 5214 23456
rect 5214 23416 5239 23456
rect 4985 23393 5071 23416
rect 5153 23393 5239 23416
rect 20105 23456 20191 23479
rect 20273 23456 20359 23479
rect 20105 23416 20130 23456
rect 20130 23416 20170 23456
rect 20170 23416 20191 23456
rect 20273 23416 20294 23456
rect 20294 23416 20334 23456
rect 20334 23416 20359 23456
rect 20105 23393 20191 23416
rect 20273 23393 20359 23416
rect 3745 22700 3831 22723
rect 3913 22700 3999 22723
rect 3745 22660 3770 22700
rect 3770 22660 3810 22700
rect 3810 22660 3831 22700
rect 3913 22660 3934 22700
rect 3934 22660 3974 22700
rect 3974 22660 3999 22700
rect 3745 22637 3831 22660
rect 3913 22637 3999 22660
rect 18865 22700 18951 22723
rect 19033 22700 19119 22723
rect 18865 22660 18890 22700
rect 18890 22660 18930 22700
rect 18930 22660 18951 22700
rect 19033 22660 19054 22700
rect 19054 22660 19094 22700
rect 19094 22660 19119 22700
rect 18865 22637 18951 22660
rect 19033 22637 19119 22660
rect 4985 21944 5071 21967
rect 5153 21944 5239 21967
rect 4985 21904 5010 21944
rect 5010 21904 5050 21944
rect 5050 21904 5071 21944
rect 5153 21904 5174 21944
rect 5174 21904 5214 21944
rect 5214 21904 5239 21944
rect 4985 21881 5071 21904
rect 5153 21881 5239 21904
rect 20105 21944 20191 21967
rect 20273 21944 20359 21967
rect 20105 21904 20130 21944
rect 20130 21904 20170 21944
rect 20170 21904 20191 21944
rect 20273 21904 20294 21944
rect 20294 21904 20334 21944
rect 20334 21904 20359 21944
rect 20105 21881 20191 21904
rect 20273 21881 20359 21904
rect 3745 21188 3831 21211
rect 3913 21188 3999 21211
rect 3745 21148 3770 21188
rect 3770 21148 3810 21188
rect 3810 21148 3831 21188
rect 3913 21148 3934 21188
rect 3934 21148 3974 21188
rect 3974 21148 3999 21188
rect 3745 21125 3831 21148
rect 3913 21125 3999 21148
rect 18865 21188 18951 21211
rect 19033 21188 19119 21211
rect 18865 21148 18890 21188
rect 18890 21148 18930 21188
rect 18930 21148 18951 21188
rect 19033 21148 19054 21188
rect 19054 21148 19094 21188
rect 19094 21148 19119 21188
rect 18865 21125 18951 21148
rect 19033 21125 19119 21148
rect 4985 20432 5071 20455
rect 5153 20432 5239 20455
rect 4985 20392 5010 20432
rect 5010 20392 5050 20432
rect 5050 20392 5071 20432
rect 5153 20392 5174 20432
rect 5174 20392 5214 20432
rect 5214 20392 5239 20432
rect 4985 20369 5071 20392
rect 5153 20369 5239 20392
rect 20105 20432 20191 20455
rect 20273 20432 20359 20455
rect 20105 20392 20130 20432
rect 20130 20392 20170 20432
rect 20170 20392 20191 20432
rect 20273 20392 20294 20432
rect 20294 20392 20334 20432
rect 20334 20392 20359 20432
rect 20105 20369 20191 20392
rect 20273 20369 20359 20392
rect 3745 19676 3831 19699
rect 3913 19676 3999 19699
rect 3745 19636 3770 19676
rect 3770 19636 3810 19676
rect 3810 19636 3831 19676
rect 3913 19636 3934 19676
rect 3934 19636 3974 19676
rect 3974 19636 3999 19676
rect 3745 19613 3831 19636
rect 3913 19613 3999 19636
rect 18865 19676 18951 19699
rect 19033 19676 19119 19699
rect 18865 19636 18890 19676
rect 18890 19636 18930 19676
rect 18930 19636 18951 19676
rect 19033 19636 19054 19676
rect 19054 19636 19094 19676
rect 19094 19636 19119 19676
rect 18865 19613 18951 19636
rect 19033 19613 19119 19636
rect 4985 18920 5071 18943
rect 5153 18920 5239 18943
rect 4985 18880 5010 18920
rect 5010 18880 5050 18920
rect 5050 18880 5071 18920
rect 5153 18880 5174 18920
rect 5174 18880 5214 18920
rect 5214 18880 5239 18920
rect 4985 18857 5071 18880
rect 5153 18857 5239 18880
rect 20105 18920 20191 18943
rect 20273 18920 20359 18943
rect 20105 18880 20130 18920
rect 20130 18880 20170 18920
rect 20170 18880 20191 18920
rect 20273 18880 20294 18920
rect 20294 18880 20334 18920
rect 20334 18880 20359 18920
rect 20105 18857 20191 18880
rect 20273 18857 20359 18880
rect 3745 18164 3831 18187
rect 3913 18164 3999 18187
rect 3745 18124 3770 18164
rect 3770 18124 3810 18164
rect 3810 18124 3831 18164
rect 3913 18124 3934 18164
rect 3934 18124 3974 18164
rect 3974 18124 3999 18164
rect 3745 18101 3831 18124
rect 3913 18101 3999 18124
rect 18865 18164 18951 18187
rect 19033 18164 19119 18187
rect 18865 18124 18890 18164
rect 18890 18124 18930 18164
rect 18930 18124 18951 18164
rect 19033 18124 19054 18164
rect 19054 18124 19094 18164
rect 19094 18124 19119 18164
rect 18865 18101 18951 18124
rect 19033 18101 19119 18124
rect 13509 17597 13595 17683
rect 4985 17408 5071 17431
rect 5153 17408 5239 17431
rect 4985 17368 5010 17408
rect 5010 17368 5050 17408
rect 5050 17368 5071 17408
rect 5153 17368 5174 17408
rect 5174 17368 5214 17408
rect 5214 17368 5239 17408
rect 4985 17345 5071 17368
rect 5153 17345 5239 17368
rect 20105 17408 20191 17431
rect 20273 17408 20359 17431
rect 20105 17368 20130 17408
rect 20130 17368 20170 17408
rect 20170 17368 20191 17408
rect 20273 17368 20294 17408
rect 20294 17368 20334 17408
rect 20334 17368 20359 17408
rect 20105 17345 20191 17368
rect 20273 17345 20359 17368
rect 3745 16652 3831 16675
rect 3913 16652 3999 16675
rect 3745 16612 3770 16652
rect 3770 16612 3810 16652
rect 3810 16612 3831 16652
rect 3913 16612 3934 16652
rect 3934 16612 3974 16652
rect 3974 16612 3999 16652
rect 3745 16589 3831 16612
rect 3913 16589 3999 16612
rect 18865 16652 18951 16675
rect 19033 16652 19119 16675
rect 18865 16612 18890 16652
rect 18890 16612 18930 16652
rect 18930 16612 18951 16652
rect 19033 16612 19054 16652
rect 19054 16612 19094 16652
rect 19094 16612 19119 16652
rect 18865 16589 18951 16612
rect 19033 16589 19119 16612
rect 4985 15896 5071 15919
rect 5153 15896 5239 15919
rect 4985 15856 5010 15896
rect 5010 15856 5050 15896
rect 5050 15856 5071 15896
rect 5153 15856 5174 15896
rect 5174 15856 5214 15896
rect 5214 15856 5239 15896
rect 4985 15833 5071 15856
rect 5153 15833 5239 15856
rect 20105 15896 20191 15919
rect 20273 15896 20359 15919
rect 20105 15856 20130 15896
rect 20130 15856 20170 15896
rect 20170 15856 20191 15896
rect 20273 15856 20294 15896
rect 20294 15856 20334 15896
rect 20334 15856 20359 15896
rect 20105 15833 20191 15856
rect 20273 15833 20359 15856
rect 14877 15665 14963 15751
rect 3745 15140 3831 15163
rect 3913 15140 3999 15163
rect 3745 15100 3770 15140
rect 3770 15100 3810 15140
rect 3810 15100 3831 15140
rect 3913 15100 3934 15140
rect 3934 15100 3974 15140
rect 3974 15100 3999 15140
rect 3745 15077 3831 15100
rect 3913 15077 3999 15100
rect 18865 15140 18951 15163
rect 19033 15140 19119 15163
rect 18865 15100 18890 15140
rect 18890 15100 18930 15140
rect 18930 15100 18951 15140
rect 19033 15100 19054 15140
rect 19054 15100 19094 15140
rect 19094 15100 19119 15140
rect 18865 15077 18951 15100
rect 19033 15077 19119 15100
rect 4985 14384 5071 14407
rect 5153 14384 5239 14407
rect 4985 14344 5010 14384
rect 5010 14344 5050 14384
rect 5050 14344 5071 14384
rect 5153 14344 5174 14384
rect 5174 14344 5214 14384
rect 5214 14344 5239 14384
rect 4985 14321 5071 14344
rect 5153 14321 5239 14344
rect 20105 14384 20191 14407
rect 20273 14384 20359 14407
rect 20105 14344 20130 14384
rect 20130 14344 20170 14384
rect 20170 14344 20191 14384
rect 20273 14344 20294 14384
rect 20294 14344 20334 14384
rect 20334 14344 20359 14384
rect 20105 14321 20191 14344
rect 20273 14321 20359 14344
rect 3745 13628 3831 13651
rect 3913 13628 3999 13651
rect 3745 13588 3770 13628
rect 3770 13588 3810 13628
rect 3810 13588 3831 13628
rect 3913 13588 3934 13628
rect 3934 13588 3974 13628
rect 3974 13588 3999 13628
rect 3745 13565 3831 13588
rect 3913 13565 3999 13588
rect 18865 13628 18951 13651
rect 19033 13628 19119 13651
rect 18865 13588 18890 13628
rect 18890 13588 18930 13628
rect 18930 13588 18951 13628
rect 19033 13588 19054 13628
rect 19054 13588 19094 13628
rect 19094 13588 19119 13628
rect 18865 13565 18951 13588
rect 19033 13565 19119 13588
rect 4985 12872 5071 12895
rect 5153 12872 5239 12895
rect 4985 12832 5010 12872
rect 5010 12832 5050 12872
rect 5050 12832 5071 12872
rect 5153 12832 5174 12872
rect 5174 12832 5214 12872
rect 5214 12832 5239 12872
rect 4985 12809 5071 12832
rect 5153 12809 5239 12832
rect 20105 12872 20191 12895
rect 20273 12872 20359 12895
rect 20105 12832 20130 12872
rect 20130 12832 20170 12872
rect 20170 12832 20191 12872
rect 20273 12832 20294 12872
rect 20294 12832 20334 12872
rect 20334 12832 20359 12872
rect 20105 12809 20191 12832
rect 20273 12809 20359 12832
rect 3745 12116 3831 12139
rect 3913 12116 3999 12139
rect 3745 12076 3770 12116
rect 3770 12076 3810 12116
rect 3810 12076 3831 12116
rect 3913 12076 3934 12116
rect 3934 12076 3974 12116
rect 3974 12076 3999 12116
rect 3745 12053 3831 12076
rect 3913 12053 3999 12076
rect 18865 12116 18951 12139
rect 19033 12116 19119 12139
rect 18865 12076 18890 12116
rect 18890 12076 18930 12116
rect 18930 12076 18951 12116
rect 19033 12076 19054 12116
rect 19054 12076 19094 12116
rect 19094 12076 19119 12116
rect 18865 12053 18951 12076
rect 19033 12053 19119 12076
rect 4985 11360 5071 11383
rect 5153 11360 5239 11383
rect 4985 11320 5010 11360
rect 5010 11320 5050 11360
rect 5050 11320 5071 11360
rect 5153 11320 5174 11360
rect 5174 11320 5214 11360
rect 5214 11320 5239 11360
rect 4985 11297 5071 11320
rect 5153 11297 5239 11320
rect 20105 11360 20191 11383
rect 20273 11360 20359 11383
rect 20105 11320 20130 11360
rect 20130 11320 20170 11360
rect 20170 11320 20191 11360
rect 20273 11320 20294 11360
rect 20294 11320 20334 11360
rect 20334 11320 20359 11360
rect 20105 11297 20191 11320
rect 20273 11297 20359 11320
rect 8493 11045 8579 11131
rect 3745 10604 3831 10627
rect 3913 10604 3999 10627
rect 3745 10564 3770 10604
rect 3770 10564 3810 10604
rect 3810 10564 3831 10604
rect 3913 10564 3934 10604
rect 3934 10564 3974 10604
rect 3974 10564 3999 10604
rect 3745 10541 3831 10564
rect 3913 10541 3999 10564
rect 18865 10604 18951 10627
rect 19033 10604 19119 10627
rect 18865 10564 18890 10604
rect 18890 10564 18930 10604
rect 18930 10564 18951 10604
rect 19033 10564 19054 10604
rect 19054 10564 19094 10604
rect 19094 10564 19119 10604
rect 18865 10541 18951 10564
rect 19033 10541 19119 10564
rect 9405 10205 9491 10291
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 13509 2645 13595 2731
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 2109 2057 2195 2143
rect 7125 2057 7211 2143
rect 12141 2057 12227 2143
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 17157 881 17243 967
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 20105 713 20191 736
rect 20273 713 20359 736
rect 10317 125 10403 211
<< metal6 >>
rect 3652 84715 4092 86016
rect 3652 84629 3745 84715
rect 3831 84629 3913 84715
rect 3999 84629 4092 84715
rect 1988 83539 2316 83660
rect 1988 83453 2109 83539
rect 2195 83453 2316 83539
rect 1076 76567 1404 76688
rect 1076 76481 1197 76567
rect 1283 76481 1404 76567
rect 1076 34399 1404 76481
rect 1988 47923 2316 83453
rect 1988 47837 2109 47923
rect 2195 47837 2316 47923
rect 1988 47716 2316 47837
rect 3652 83203 4092 84629
rect 3652 83117 3745 83203
rect 3831 83117 3913 83203
rect 3999 83117 4092 83203
rect 3652 81691 4092 83117
rect 3652 81605 3745 81691
rect 3831 81605 3913 81691
rect 3999 81605 4092 81691
rect 3652 80179 4092 81605
rect 3652 80093 3745 80179
rect 3831 80093 3913 80179
rect 3999 80093 4092 80179
rect 3652 78667 4092 80093
rect 3652 78581 3745 78667
rect 3831 78581 3913 78667
rect 3999 78581 4092 78667
rect 3652 77155 4092 78581
rect 3652 77069 3745 77155
rect 3831 77069 3913 77155
rect 3999 77069 4092 77155
rect 3652 75643 4092 77069
rect 3652 75557 3745 75643
rect 3831 75557 3913 75643
rect 3999 75557 4092 75643
rect 3652 74131 4092 75557
rect 3652 74045 3745 74131
rect 3831 74045 3913 74131
rect 3999 74045 4092 74131
rect 3652 72619 4092 74045
rect 3652 72533 3745 72619
rect 3831 72533 3913 72619
rect 3999 72533 4092 72619
rect 3652 71107 4092 72533
rect 3652 71021 3745 71107
rect 3831 71021 3913 71107
rect 3999 71021 4092 71107
rect 3652 69595 4092 71021
rect 3652 69509 3745 69595
rect 3831 69509 3913 69595
rect 3999 69509 4092 69595
rect 3652 68083 4092 69509
rect 3652 67997 3745 68083
rect 3831 67997 3913 68083
rect 3999 67997 4092 68083
rect 3652 66571 4092 67997
rect 3652 66485 3745 66571
rect 3831 66485 3913 66571
rect 3999 66485 4092 66571
rect 3652 65059 4092 66485
rect 3652 64973 3745 65059
rect 3831 64973 3913 65059
rect 3999 64973 4092 65059
rect 3652 63547 4092 64973
rect 3652 63461 3745 63547
rect 3831 63461 3913 63547
rect 3999 63461 4092 63547
rect 3652 62035 4092 63461
rect 3652 61949 3745 62035
rect 3831 61949 3913 62035
rect 3999 61949 4092 62035
rect 3652 60523 4092 61949
rect 3652 60437 3745 60523
rect 3831 60437 3913 60523
rect 3999 60437 4092 60523
rect 3652 59011 4092 60437
rect 3652 58925 3745 59011
rect 3831 58925 3913 59011
rect 3999 58925 4092 59011
rect 3652 57499 4092 58925
rect 3652 57413 3745 57499
rect 3831 57413 3913 57499
rect 3999 57413 4092 57499
rect 3652 55987 4092 57413
rect 3652 55901 3745 55987
rect 3831 55901 3913 55987
rect 3999 55901 4092 55987
rect 3652 54475 4092 55901
rect 3652 54389 3745 54475
rect 3831 54389 3913 54475
rect 3999 54389 4092 54475
rect 3652 52963 4092 54389
rect 3652 52877 3745 52963
rect 3831 52877 3913 52963
rect 3999 52877 4092 52963
rect 3652 51451 4092 52877
rect 3652 51365 3745 51451
rect 3831 51365 3913 51451
rect 3999 51365 4092 51451
rect 3652 49939 4092 51365
rect 3652 49853 3745 49939
rect 3831 49853 3913 49939
rect 3999 49853 4092 49939
rect 3652 48427 4092 49853
rect 3652 48341 3745 48427
rect 3831 48341 3913 48427
rect 3999 48341 4092 48427
rect 3652 46915 4092 48341
rect 3652 46829 3745 46915
rect 3831 46829 3913 46915
rect 3999 46829 4092 46915
rect 1076 34313 1197 34399
rect 1283 34313 1404 34399
rect 1076 34192 1404 34313
rect 1988 45991 2316 46112
rect 1988 45905 2109 45991
rect 2195 45905 2316 45991
rect 1988 2143 2316 45905
rect 1988 2057 2109 2143
rect 2195 2057 2316 2143
rect 1988 1936 2316 2057
rect 3652 45403 4092 46829
rect 3652 45317 3745 45403
rect 3831 45317 3913 45403
rect 3999 45317 4092 45403
rect 3652 43891 4092 45317
rect 3652 43805 3745 43891
rect 3831 43805 3913 43891
rect 3999 43805 4092 43891
rect 3652 42379 4092 43805
rect 3652 42293 3745 42379
rect 3831 42293 3913 42379
rect 3999 42293 4092 42379
rect 3652 40867 4092 42293
rect 3652 40781 3745 40867
rect 3831 40781 3913 40867
rect 3999 40781 4092 40867
rect 3652 39355 4092 40781
rect 3652 39269 3745 39355
rect 3831 39269 3913 39355
rect 3999 39269 4092 39355
rect 3652 37843 4092 39269
rect 3652 37757 3745 37843
rect 3831 37757 3913 37843
rect 3999 37757 4092 37843
rect 3652 36331 4092 37757
rect 3652 36245 3745 36331
rect 3831 36245 3913 36331
rect 3999 36245 4092 36331
rect 3652 34819 4092 36245
rect 3652 34733 3745 34819
rect 3831 34733 3913 34819
rect 3999 34733 4092 34819
rect 3652 33307 4092 34733
rect 3652 33221 3745 33307
rect 3831 33221 3913 33307
rect 3999 33221 4092 33307
rect 3652 31795 4092 33221
rect 3652 31709 3745 31795
rect 3831 31709 3913 31795
rect 3999 31709 4092 31795
rect 3652 30283 4092 31709
rect 3652 30197 3745 30283
rect 3831 30197 3913 30283
rect 3999 30197 4092 30283
rect 3652 28771 4092 30197
rect 3652 28685 3745 28771
rect 3831 28685 3913 28771
rect 3999 28685 4092 28771
rect 3652 27259 4092 28685
rect 3652 27173 3745 27259
rect 3831 27173 3913 27259
rect 3999 27173 4092 27259
rect 3652 25747 4092 27173
rect 3652 25661 3745 25747
rect 3831 25661 3913 25747
rect 3999 25661 4092 25747
rect 3652 24235 4092 25661
rect 3652 24149 3745 24235
rect 3831 24149 3913 24235
rect 3999 24149 4092 24235
rect 3652 22723 4092 24149
rect 3652 22637 3745 22723
rect 3831 22637 3913 22723
rect 3999 22637 4092 22723
rect 3652 21211 4092 22637
rect 3652 21125 3745 21211
rect 3831 21125 3913 21211
rect 3999 21125 4092 21211
rect 3652 19699 4092 21125
rect 3652 19613 3745 19699
rect 3831 19613 3913 19699
rect 3999 19613 4092 19699
rect 3652 18187 4092 19613
rect 3652 18101 3745 18187
rect 3831 18101 3913 18187
rect 3999 18101 4092 18187
rect 3652 16675 4092 18101
rect 3652 16589 3745 16675
rect 3831 16589 3913 16675
rect 3999 16589 4092 16675
rect 3652 15163 4092 16589
rect 3652 15077 3745 15163
rect 3831 15077 3913 15163
rect 3999 15077 4092 15163
rect 3652 13651 4092 15077
rect 3652 13565 3745 13651
rect 3831 13565 3913 13651
rect 3999 13565 4092 13651
rect 3652 12139 4092 13565
rect 3652 12053 3745 12139
rect 3831 12053 3913 12139
rect 3999 12053 4092 12139
rect 3652 10627 4092 12053
rect 3652 10541 3745 10627
rect 3831 10541 3913 10627
rect 3999 10541 4092 10627
rect 3652 9115 4092 10541
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 3652 0 4092 1469
rect 4892 83959 5332 86016
rect 12020 85891 12348 86012
rect 12020 85805 12141 85891
rect 12227 85805 12348 85891
rect 4892 83873 4985 83959
rect 5071 83873 5153 83959
rect 5239 83873 5332 83959
rect 4892 82447 5332 83873
rect 4892 82361 4985 82447
rect 5071 82361 5153 82447
rect 5239 82361 5332 82447
rect 4892 80935 5332 82361
rect 4892 80849 4985 80935
rect 5071 80849 5153 80935
rect 5239 80849 5332 80935
rect 4892 79423 5332 80849
rect 4892 79337 4985 79423
rect 5071 79337 5153 79423
rect 5239 79337 5332 79423
rect 4892 77911 5332 79337
rect 4892 77825 4985 77911
rect 5071 77825 5153 77911
rect 5239 77825 5332 77911
rect 4892 76399 5332 77825
rect 4892 76313 4985 76399
rect 5071 76313 5153 76399
rect 5239 76313 5332 76399
rect 4892 74887 5332 76313
rect 4892 74801 4985 74887
rect 5071 74801 5153 74887
rect 5239 74801 5332 74887
rect 4892 73375 5332 74801
rect 4892 73289 4985 73375
rect 5071 73289 5153 73375
rect 5239 73289 5332 73375
rect 4892 71863 5332 73289
rect 4892 71777 4985 71863
rect 5071 71777 5153 71863
rect 5239 71777 5332 71863
rect 4892 70351 5332 71777
rect 4892 70265 4985 70351
rect 5071 70265 5153 70351
rect 5239 70265 5332 70351
rect 4892 68839 5332 70265
rect 4892 68753 4985 68839
rect 5071 68753 5153 68839
rect 5239 68753 5332 68839
rect 4892 67327 5332 68753
rect 4892 67241 4985 67327
rect 5071 67241 5153 67327
rect 5239 67241 5332 67327
rect 4892 65815 5332 67241
rect 4892 65729 4985 65815
rect 5071 65729 5153 65815
rect 5239 65729 5332 65815
rect 4892 64303 5332 65729
rect 4892 64217 4985 64303
rect 5071 64217 5153 64303
rect 5239 64217 5332 64303
rect 4892 62791 5332 64217
rect 4892 62705 4985 62791
rect 5071 62705 5153 62791
rect 5239 62705 5332 62791
rect 4892 61279 5332 62705
rect 4892 61193 4985 61279
rect 5071 61193 5153 61279
rect 5239 61193 5332 61279
rect 4892 59767 5332 61193
rect 4892 59681 4985 59767
rect 5071 59681 5153 59767
rect 5239 59681 5332 59767
rect 4892 58255 5332 59681
rect 4892 58169 4985 58255
rect 5071 58169 5153 58255
rect 5239 58169 5332 58255
rect 4892 56743 5332 58169
rect 4892 56657 4985 56743
rect 5071 56657 5153 56743
rect 5239 56657 5332 56743
rect 4892 55231 5332 56657
rect 4892 55145 4985 55231
rect 5071 55145 5153 55231
rect 5239 55145 5332 55231
rect 4892 53719 5332 55145
rect 4892 53633 4985 53719
rect 5071 53633 5153 53719
rect 5239 53633 5332 53719
rect 4892 52207 5332 53633
rect 4892 52121 4985 52207
rect 5071 52121 5153 52207
rect 5239 52121 5332 52207
rect 4892 50695 5332 52121
rect 4892 50609 4985 50695
rect 5071 50609 5153 50695
rect 5239 50609 5332 50695
rect 4892 49183 5332 50609
rect 4892 49097 4985 49183
rect 5071 49097 5153 49183
rect 5239 49097 5332 49183
rect 4892 47671 5332 49097
rect 4892 47585 4985 47671
rect 5071 47585 5153 47671
rect 5239 47585 5332 47671
rect 4892 46159 5332 47585
rect 4892 46073 4985 46159
rect 5071 46073 5153 46159
rect 5239 46073 5332 46159
rect 4892 44647 5332 46073
rect 4892 44561 4985 44647
rect 5071 44561 5153 44647
rect 5239 44561 5332 44647
rect 4892 43135 5332 44561
rect 4892 43049 4985 43135
rect 5071 43049 5153 43135
rect 5239 43049 5332 43135
rect 4892 41623 5332 43049
rect 4892 41537 4985 41623
rect 5071 41537 5153 41623
rect 5239 41537 5332 41623
rect 4892 40111 5332 41537
rect 4892 40025 4985 40111
rect 5071 40025 5153 40111
rect 5239 40025 5332 40111
rect 4892 38599 5332 40025
rect 4892 38513 4985 38599
rect 5071 38513 5153 38599
rect 5239 38513 5332 38599
rect 4892 37087 5332 38513
rect 4892 37001 4985 37087
rect 5071 37001 5153 37087
rect 5239 37001 5332 37087
rect 4892 35575 5332 37001
rect 4892 35489 4985 35575
rect 5071 35489 5153 35575
rect 5239 35489 5332 35575
rect 4892 34063 5332 35489
rect 4892 33977 4985 34063
rect 5071 33977 5153 34063
rect 5239 33977 5332 34063
rect 4892 32551 5332 33977
rect 4892 32465 4985 32551
rect 5071 32465 5153 32551
rect 5239 32465 5332 32551
rect 4892 31039 5332 32465
rect 4892 30953 4985 31039
rect 5071 30953 5153 31039
rect 5239 30953 5332 31039
rect 4892 29527 5332 30953
rect 4892 29441 4985 29527
rect 5071 29441 5153 29527
rect 5239 29441 5332 29527
rect 4892 28015 5332 29441
rect 4892 27929 4985 28015
rect 5071 27929 5153 28015
rect 5239 27929 5332 28015
rect 4892 26503 5332 27929
rect 4892 26417 4985 26503
rect 5071 26417 5153 26503
rect 5239 26417 5332 26503
rect 4892 24991 5332 26417
rect 4892 24905 4985 24991
rect 5071 24905 5153 24991
rect 5239 24905 5332 24991
rect 4892 23479 5332 24905
rect 4892 23393 4985 23479
rect 5071 23393 5153 23479
rect 5239 23393 5332 23479
rect 4892 21967 5332 23393
rect 4892 21881 4985 21967
rect 5071 21881 5153 21967
rect 5239 21881 5332 21967
rect 4892 20455 5332 21881
rect 4892 20369 4985 20455
rect 5071 20369 5153 20455
rect 5239 20369 5332 20455
rect 4892 18943 5332 20369
rect 4892 18857 4985 18943
rect 5071 18857 5153 18943
rect 5239 18857 5332 18943
rect 4892 17431 5332 18857
rect 4892 17345 4985 17431
rect 5071 17345 5153 17431
rect 5239 17345 5332 17431
rect 4892 15919 5332 17345
rect 4892 15833 4985 15919
rect 5071 15833 5153 15919
rect 5239 15833 5332 15919
rect 4892 14407 5332 15833
rect 4892 14321 4985 14407
rect 5071 14321 5153 14407
rect 5239 14321 5332 14407
rect 4892 12895 5332 14321
rect 4892 12809 4985 12895
rect 5071 12809 5153 12895
rect 5239 12809 5332 12895
rect 4892 11383 5332 12809
rect 4892 11297 4985 11383
rect 5071 11297 5153 11383
rect 5239 11297 5332 11383
rect 4892 9871 5332 11297
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 7004 84463 7332 84584
rect 7004 84377 7125 84463
rect 7211 84377 7332 84463
rect 7004 2143 7332 84377
rect 8372 76735 8700 76856
rect 8372 76649 8493 76735
rect 8579 76649 8700 76735
rect 8372 11131 8700 76649
rect 8372 11045 8493 11131
rect 8579 11045 8700 11131
rect 8372 10924 8700 11045
rect 9284 76735 9612 76856
rect 9284 76649 9405 76735
rect 9491 76649 9612 76735
rect 9284 10291 9612 76649
rect 9284 10205 9405 10291
rect 9491 10205 9612 10291
rect 9284 10084 9612 10205
rect 10196 41959 10524 42080
rect 10196 41873 10317 41959
rect 10403 41873 10524 41959
rect 7004 2057 7125 2143
rect 7211 2057 7332 2143
rect 7004 1936 7332 2057
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 4892 0 5332 713
rect 10196 211 10524 41873
rect 12020 2143 12348 85805
rect 17036 85807 17364 85928
rect 17036 85721 17157 85807
rect 17243 85721 17364 85807
rect 16124 85135 16452 85256
rect 16124 85049 16245 85135
rect 16331 85049 16452 85135
rect 14756 84463 15084 84584
rect 14756 84377 14877 84463
rect 14963 84377 15084 84463
rect 13388 17683 13716 17804
rect 13388 17597 13509 17683
rect 13595 17597 13716 17683
rect 13388 2731 13716 17597
rect 14756 15751 15084 84377
rect 16124 24655 16452 85049
rect 16124 24569 16245 24655
rect 16331 24569 16452 24655
rect 16124 24448 16452 24569
rect 14756 15665 14877 15751
rect 14963 15665 15084 15751
rect 14756 15544 15084 15665
rect 13388 2645 13509 2731
rect 13595 2645 13716 2731
rect 13388 2524 13716 2645
rect 12020 2057 12141 2143
rect 12227 2057 12348 2143
rect 12020 1936 12348 2057
rect 17036 967 17364 85721
rect 17036 881 17157 967
rect 17243 881 17364 967
rect 17036 760 17364 881
rect 18772 84715 19212 86016
rect 18772 84629 18865 84715
rect 18951 84629 19033 84715
rect 19119 84629 19212 84715
rect 18772 83203 19212 84629
rect 18772 83117 18865 83203
rect 18951 83117 19033 83203
rect 19119 83117 19212 83203
rect 18772 81691 19212 83117
rect 18772 81605 18865 81691
rect 18951 81605 19033 81691
rect 19119 81605 19212 81691
rect 18772 80179 19212 81605
rect 18772 80093 18865 80179
rect 18951 80093 19033 80179
rect 19119 80093 19212 80179
rect 18772 78667 19212 80093
rect 18772 78581 18865 78667
rect 18951 78581 19033 78667
rect 19119 78581 19212 78667
rect 18772 77155 19212 78581
rect 18772 77069 18865 77155
rect 18951 77069 19033 77155
rect 19119 77069 19212 77155
rect 18772 75643 19212 77069
rect 18772 75557 18865 75643
rect 18951 75557 19033 75643
rect 19119 75557 19212 75643
rect 18772 74131 19212 75557
rect 18772 74045 18865 74131
rect 18951 74045 19033 74131
rect 19119 74045 19212 74131
rect 18772 72619 19212 74045
rect 18772 72533 18865 72619
rect 18951 72533 19033 72619
rect 19119 72533 19212 72619
rect 18772 71107 19212 72533
rect 18772 71021 18865 71107
rect 18951 71021 19033 71107
rect 19119 71021 19212 71107
rect 18772 69595 19212 71021
rect 18772 69509 18865 69595
rect 18951 69509 19033 69595
rect 19119 69509 19212 69595
rect 18772 68083 19212 69509
rect 18772 67997 18865 68083
rect 18951 67997 19033 68083
rect 19119 67997 19212 68083
rect 18772 66571 19212 67997
rect 18772 66485 18865 66571
rect 18951 66485 19033 66571
rect 19119 66485 19212 66571
rect 18772 65059 19212 66485
rect 18772 64973 18865 65059
rect 18951 64973 19033 65059
rect 19119 64973 19212 65059
rect 18772 63547 19212 64973
rect 18772 63461 18865 63547
rect 18951 63461 19033 63547
rect 19119 63461 19212 63547
rect 18772 62035 19212 63461
rect 18772 61949 18865 62035
rect 18951 61949 19033 62035
rect 19119 61949 19212 62035
rect 18772 60523 19212 61949
rect 18772 60437 18865 60523
rect 18951 60437 19033 60523
rect 19119 60437 19212 60523
rect 18772 59011 19212 60437
rect 18772 58925 18865 59011
rect 18951 58925 19033 59011
rect 19119 58925 19212 59011
rect 18772 57499 19212 58925
rect 18772 57413 18865 57499
rect 18951 57413 19033 57499
rect 19119 57413 19212 57499
rect 18772 55987 19212 57413
rect 18772 55901 18865 55987
rect 18951 55901 19033 55987
rect 19119 55901 19212 55987
rect 18772 54475 19212 55901
rect 18772 54389 18865 54475
rect 18951 54389 19033 54475
rect 19119 54389 19212 54475
rect 18772 52963 19212 54389
rect 18772 52877 18865 52963
rect 18951 52877 19033 52963
rect 19119 52877 19212 52963
rect 18772 51451 19212 52877
rect 18772 51365 18865 51451
rect 18951 51365 19033 51451
rect 19119 51365 19212 51451
rect 18772 49939 19212 51365
rect 18772 49853 18865 49939
rect 18951 49853 19033 49939
rect 19119 49853 19212 49939
rect 18772 48427 19212 49853
rect 18772 48341 18865 48427
rect 18951 48341 19033 48427
rect 19119 48341 19212 48427
rect 18772 46915 19212 48341
rect 18772 46829 18865 46915
rect 18951 46829 19033 46915
rect 19119 46829 19212 46915
rect 18772 45403 19212 46829
rect 18772 45317 18865 45403
rect 18951 45317 19033 45403
rect 19119 45317 19212 45403
rect 18772 43891 19212 45317
rect 18772 43805 18865 43891
rect 18951 43805 19033 43891
rect 19119 43805 19212 43891
rect 18772 42379 19212 43805
rect 18772 42293 18865 42379
rect 18951 42293 19033 42379
rect 19119 42293 19212 42379
rect 18772 40867 19212 42293
rect 18772 40781 18865 40867
rect 18951 40781 19033 40867
rect 19119 40781 19212 40867
rect 18772 39355 19212 40781
rect 18772 39269 18865 39355
rect 18951 39269 19033 39355
rect 19119 39269 19212 39355
rect 18772 37843 19212 39269
rect 18772 37757 18865 37843
rect 18951 37757 19033 37843
rect 19119 37757 19212 37843
rect 18772 36331 19212 37757
rect 18772 36245 18865 36331
rect 18951 36245 19033 36331
rect 19119 36245 19212 36331
rect 18772 34819 19212 36245
rect 18772 34733 18865 34819
rect 18951 34733 19033 34819
rect 19119 34733 19212 34819
rect 18772 33307 19212 34733
rect 18772 33221 18865 33307
rect 18951 33221 19033 33307
rect 19119 33221 19212 33307
rect 18772 31795 19212 33221
rect 18772 31709 18865 31795
rect 18951 31709 19033 31795
rect 19119 31709 19212 31795
rect 18772 30283 19212 31709
rect 18772 30197 18865 30283
rect 18951 30197 19033 30283
rect 19119 30197 19212 30283
rect 18772 28771 19212 30197
rect 18772 28685 18865 28771
rect 18951 28685 19033 28771
rect 19119 28685 19212 28771
rect 18772 27259 19212 28685
rect 18772 27173 18865 27259
rect 18951 27173 19033 27259
rect 19119 27173 19212 27259
rect 18772 25747 19212 27173
rect 18772 25661 18865 25747
rect 18951 25661 19033 25747
rect 19119 25661 19212 25747
rect 18772 24235 19212 25661
rect 18772 24149 18865 24235
rect 18951 24149 19033 24235
rect 19119 24149 19212 24235
rect 18772 22723 19212 24149
rect 18772 22637 18865 22723
rect 18951 22637 19033 22723
rect 19119 22637 19212 22723
rect 18772 21211 19212 22637
rect 18772 21125 18865 21211
rect 18951 21125 19033 21211
rect 19119 21125 19212 21211
rect 18772 19699 19212 21125
rect 18772 19613 18865 19699
rect 18951 19613 19033 19699
rect 19119 19613 19212 19699
rect 18772 18187 19212 19613
rect 18772 18101 18865 18187
rect 18951 18101 19033 18187
rect 19119 18101 19212 18187
rect 18772 16675 19212 18101
rect 18772 16589 18865 16675
rect 18951 16589 19033 16675
rect 19119 16589 19212 16675
rect 18772 15163 19212 16589
rect 18772 15077 18865 15163
rect 18951 15077 19033 15163
rect 19119 15077 19212 15163
rect 18772 13651 19212 15077
rect 18772 13565 18865 13651
rect 18951 13565 19033 13651
rect 19119 13565 19212 13651
rect 18772 12139 19212 13565
rect 18772 12053 18865 12139
rect 18951 12053 19033 12139
rect 19119 12053 19212 12139
rect 18772 10627 19212 12053
rect 18772 10541 18865 10627
rect 18951 10541 19033 10627
rect 19119 10541 19212 10627
rect 18772 9115 19212 10541
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 10196 125 10317 211
rect 10403 125 10524 211
rect 10196 4 10524 125
rect 18772 0 19212 1469
rect 20012 83959 20452 86016
rect 20012 83873 20105 83959
rect 20191 83873 20273 83959
rect 20359 83873 20452 83959
rect 20012 82447 20452 83873
rect 20012 82361 20105 82447
rect 20191 82361 20273 82447
rect 20359 82361 20452 82447
rect 20012 80935 20452 82361
rect 20012 80849 20105 80935
rect 20191 80849 20273 80935
rect 20359 80849 20452 80935
rect 20012 79423 20452 80849
rect 20012 79337 20105 79423
rect 20191 79337 20273 79423
rect 20359 79337 20452 79423
rect 20012 77911 20452 79337
rect 20012 77825 20105 77911
rect 20191 77825 20273 77911
rect 20359 77825 20452 77911
rect 20012 76399 20452 77825
rect 20012 76313 20105 76399
rect 20191 76313 20273 76399
rect 20359 76313 20452 76399
rect 20012 74887 20452 76313
rect 20012 74801 20105 74887
rect 20191 74801 20273 74887
rect 20359 74801 20452 74887
rect 20012 73375 20452 74801
rect 20012 73289 20105 73375
rect 20191 73289 20273 73375
rect 20359 73289 20452 73375
rect 20012 71863 20452 73289
rect 20012 71777 20105 71863
rect 20191 71777 20273 71863
rect 20359 71777 20452 71863
rect 20012 70351 20452 71777
rect 20012 70265 20105 70351
rect 20191 70265 20273 70351
rect 20359 70265 20452 70351
rect 20012 68839 20452 70265
rect 20012 68753 20105 68839
rect 20191 68753 20273 68839
rect 20359 68753 20452 68839
rect 20012 67327 20452 68753
rect 20012 67241 20105 67327
rect 20191 67241 20273 67327
rect 20359 67241 20452 67327
rect 20012 65815 20452 67241
rect 20012 65729 20105 65815
rect 20191 65729 20273 65815
rect 20359 65729 20452 65815
rect 20012 64303 20452 65729
rect 20012 64217 20105 64303
rect 20191 64217 20273 64303
rect 20359 64217 20452 64303
rect 20012 62791 20452 64217
rect 20012 62705 20105 62791
rect 20191 62705 20273 62791
rect 20359 62705 20452 62791
rect 20012 61279 20452 62705
rect 20012 61193 20105 61279
rect 20191 61193 20273 61279
rect 20359 61193 20452 61279
rect 20012 59767 20452 61193
rect 20012 59681 20105 59767
rect 20191 59681 20273 59767
rect 20359 59681 20452 59767
rect 20012 58255 20452 59681
rect 20012 58169 20105 58255
rect 20191 58169 20273 58255
rect 20359 58169 20452 58255
rect 20012 56743 20452 58169
rect 20012 56657 20105 56743
rect 20191 56657 20273 56743
rect 20359 56657 20452 56743
rect 20012 55231 20452 56657
rect 20012 55145 20105 55231
rect 20191 55145 20273 55231
rect 20359 55145 20452 55231
rect 20012 53719 20452 55145
rect 20012 53633 20105 53719
rect 20191 53633 20273 53719
rect 20359 53633 20452 53719
rect 20012 52207 20452 53633
rect 20012 52121 20105 52207
rect 20191 52121 20273 52207
rect 20359 52121 20452 52207
rect 20012 50695 20452 52121
rect 20012 50609 20105 50695
rect 20191 50609 20273 50695
rect 20359 50609 20452 50695
rect 20012 49183 20452 50609
rect 20012 49097 20105 49183
rect 20191 49097 20273 49183
rect 20359 49097 20452 49183
rect 20012 47671 20452 49097
rect 20012 47585 20105 47671
rect 20191 47585 20273 47671
rect 20359 47585 20452 47671
rect 20012 46159 20452 47585
rect 20012 46073 20105 46159
rect 20191 46073 20273 46159
rect 20359 46073 20452 46159
rect 20012 44647 20452 46073
rect 20012 44561 20105 44647
rect 20191 44561 20273 44647
rect 20359 44561 20452 44647
rect 20012 43135 20452 44561
rect 20012 43049 20105 43135
rect 20191 43049 20273 43135
rect 20359 43049 20452 43135
rect 20012 41623 20452 43049
rect 20012 41537 20105 41623
rect 20191 41537 20273 41623
rect 20359 41537 20452 41623
rect 20012 40111 20452 41537
rect 20012 40025 20105 40111
rect 20191 40025 20273 40111
rect 20359 40025 20452 40111
rect 20012 38599 20452 40025
rect 20012 38513 20105 38599
rect 20191 38513 20273 38599
rect 20359 38513 20452 38599
rect 20012 37087 20452 38513
rect 20012 37001 20105 37087
rect 20191 37001 20273 37087
rect 20359 37001 20452 37087
rect 20012 35575 20452 37001
rect 20012 35489 20105 35575
rect 20191 35489 20273 35575
rect 20359 35489 20452 35575
rect 20012 34063 20452 35489
rect 20012 33977 20105 34063
rect 20191 33977 20273 34063
rect 20359 33977 20452 34063
rect 20012 32551 20452 33977
rect 20012 32465 20105 32551
rect 20191 32465 20273 32551
rect 20359 32465 20452 32551
rect 20012 31039 20452 32465
rect 20012 30953 20105 31039
rect 20191 30953 20273 31039
rect 20359 30953 20452 31039
rect 20012 29527 20452 30953
rect 20012 29441 20105 29527
rect 20191 29441 20273 29527
rect 20359 29441 20452 29527
rect 20012 28015 20452 29441
rect 20012 27929 20105 28015
rect 20191 27929 20273 28015
rect 20359 27929 20452 28015
rect 20012 26503 20452 27929
rect 20012 26417 20105 26503
rect 20191 26417 20273 26503
rect 20359 26417 20452 26503
rect 20012 24991 20452 26417
rect 20012 24905 20105 24991
rect 20191 24905 20273 24991
rect 20359 24905 20452 24991
rect 20012 23479 20452 24905
rect 20012 23393 20105 23479
rect 20191 23393 20273 23479
rect 20359 23393 20452 23479
rect 20012 21967 20452 23393
rect 20012 21881 20105 21967
rect 20191 21881 20273 21967
rect 20359 21881 20452 21967
rect 20012 20455 20452 21881
rect 20012 20369 20105 20455
rect 20191 20369 20273 20455
rect 20359 20369 20452 20455
rect 20012 18943 20452 20369
rect 20012 18857 20105 18943
rect 20191 18857 20273 18943
rect 20359 18857 20452 18943
rect 20012 17431 20452 18857
rect 20012 17345 20105 17431
rect 20191 17345 20273 17431
rect 20359 17345 20452 17431
rect 20012 15919 20452 17345
rect 20012 15833 20105 15919
rect 20191 15833 20273 15919
rect 20359 15833 20452 15919
rect 20012 14407 20452 15833
rect 20012 14321 20105 14407
rect 20191 14321 20273 14407
rect 20359 14321 20452 14407
rect 20012 12895 20452 14321
rect 20012 12809 20105 12895
rect 20191 12809 20273 12895
rect 20359 12809 20452 12895
rect 20012 11383 20452 12809
rect 20012 11297 20105 11383
rect 20191 11297 20273 11383
rect 20359 11297 20452 11383
rect 20012 9871 20452 11297
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
use sg13g2_inv_1  _0357_
timestamp 1676382929
transform -1 0 3264 0 -1 55188
box -48 -56 336 834
use sg13g2_inv_1  _0358_
timestamp 1676382929
transform -1 0 5280 0 -1 56700
box -48 -56 336 834
use sg13g2_inv_1  _0359_
timestamp 1676382929
transform -1 0 15840 0 -1 58212
box -48 -56 336 834
use sg13g2_inv_1  _0360_
timestamp 1676382929
transform -1 0 14400 0 1 52164
box -48 -56 336 834
use sg13g2_inv_1  _0361_
timestamp 1676382929
transform -1 0 20352 0 -1 50652
box -48 -56 336 834
use sg13g2_inv_1  _0362_
timestamp 1676382929
transform -1 0 4224 0 -1 50652
box -48 -56 336 834
use sg13g2_inv_1  _0363_
timestamp 1676382929
transform 1 0 5280 0 -1 52164
box -48 -56 336 834
use sg13g2_inv_1  _0364_
timestamp 1676382929
transform -1 0 20352 0 -1 53676
box -48 -56 336 834
use sg13g2_inv_1  _0365_
timestamp 1676382929
transform -1 0 3840 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  _0366_
timestamp 1676382929
transform -1 0 6816 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_1  _0367_
timestamp 1676382929
transform -1 0 15456 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _0368_
timestamp 1676382929
transform -1 0 3072 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0369_
timestamp 1676382929
transform -1 0 5184 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  _0370_
timestamp 1676382929
transform -1 0 15552 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  _0371_
timestamp 1676382929
transform -1 0 17664 0 1 14364
box -48 -56 336 834
use sg13g2_inv_1  _0372_
timestamp 1676382929
transform -1 0 10464 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  _0373_
timestamp 1676382929
transform 1 0 7104 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_1  _0374_
timestamp 1676382929
transform -1 0 14976 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  _0375_
timestamp 1676382929
transform -1 0 6528 0 -1 14364
box -48 -56 336 834
use sg13g2_inv_1  _0376_
timestamp 1676382929
transform 1 0 3264 0 1 11340
box -48 -56 336 834
use sg13g2_inv_1  _0377_
timestamp 1676382929
transform 1 0 2784 0 1 9828
box -48 -56 336 834
use sg13g2_nand2b_1  _0378_
timestamp 1676567195
transform 1 0 3840 0 1 55188
box -48 -56 528 834
use sg13g2_nor3_1  _0379_
timestamp 1676639442
transform 1 0 2880 0 -1 53676
box -48 -56 528 834
use sg13g2_a221oi_1  _0380_
timestamp 1685197497
transform 1 0 3072 0 1 55188
box -48 -56 816 834
use sg13g2_mux4_1  _0381_
timestamp 1677257233
transform 1 0 2784 0 1 46116
box -48 -56 2064 834
use sg13g2_nand2b_1  _0382_
timestamp 1676567195
transform -1 0 3264 0 1 32508
box -48 -56 528 834
use sg13g2_nor3_1  _0383_
timestamp 1676639442
transform -1 0 4896 0 -1 32508
box -48 -56 528 834
use sg13g2_a221oi_1  _0384_
timestamp 1685197497
transform -1 0 4032 0 1 32508
box -48 -56 816 834
use sg13g2_mux4_1  _0385_
timestamp 1677257233
transform -1 0 5184 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0386_
timestamp 1677257233
transform 1 0 2688 0 1 61236
box -48 -56 2064 834
use sg13g2_mux4_1  _0387_
timestamp 1677257233
transform -1 0 4608 0 1 49140
box -48 -56 2064 834
use sg13g2_nand2b_1  _0388_
timestamp 1676567195
transform 1 0 4896 0 1 56700
box -48 -56 528 834
use sg13g2_nor3_1  _0389_
timestamp 1676639442
transform 1 0 3072 0 -1 58212
box -48 -56 528 834
use sg13g2_a221oi_1  _0390_
timestamp 1685197497
transform 1 0 3552 0 -1 58212
box -48 -56 816 834
use sg13g2_mux4_1  _0391_
timestamp 1677257233
transform 1 0 2976 0 1 53676
box -48 -56 2064 834
use sg13g2_nand2b_1  _0392_
timestamp 1676567195
transform -1 0 4320 0 1 15876
box -48 -56 528 834
use sg13g2_nor3_1  _0393_
timestamp 1676639442
transform 1 0 4320 0 1 17388
box -48 -56 528 834
use sg13g2_a221oi_1  _0394_
timestamp 1685197497
transform -1 0 3840 0 -1 17388
box -48 -56 816 834
use sg13g2_mux4_1  _0395_
timestamp 1677257233
transform 1 0 2784 0 1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0396_
timestamp 1677257233
transform 1 0 2592 0 -1 65772
box -48 -56 2064 834
use sg13g2_mux4_1  _0397_
timestamp 1677257233
transform 1 0 2880 0 1 56700
box -48 -56 2064 834
use sg13g2_nand2b_1  _0398_
timestamp 1676567195
transform 1 0 16896 0 1 58212
box -48 -56 528 834
use sg13g2_nor3_1  _0399_
timestamp 1676639442
transform -1 0 15552 0 1 59724
box -48 -56 528 834
use sg13g2_a221oi_1  _0400_
timestamp 1685197497
transform 1 0 15552 0 -1 59724
box -48 -56 816 834
use sg13g2_mux4_1  _0401_
timestamp 1677257233
transform 1 0 13632 0 -1 56700
box -48 -56 2064 834
use sg13g2_nand2b_1  _0402_
timestamp 1676567195
transform 1 0 14976 0 1 21924
box -48 -56 528 834
use sg13g2_nor3_1  _0403_
timestamp 1676639442
transform 1 0 14496 0 1 21924
box -48 -56 528 834
use sg13g2_a221oi_1  _0404_
timestamp 1685197497
transform 1 0 14400 0 -1 21924
box -48 -56 816 834
use sg13g2_mux4_1  _0405_
timestamp 1677257233
transform 1 0 12960 0 -1 23436
box -48 -56 2064 834
use sg13g2_mux4_1  _0406_
timestamp 1677257233
transform 1 0 12864 0 1 76356
box -48 -56 2064 834
use sg13g2_mux4_1  _0407_
timestamp 1677257233
transform 1 0 13536 0 1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0408_
timestamp 1677257233
transform -1 0 14688 0 1 49140
box -48 -56 2064 834
use sg13g2_mux2_1  _0409_
timestamp 1677247768
transform 1 0 8352 0 1 14364
box -48 -56 1008 834
use sg13g2_nor2_1  _0410_
timestamp 1676627187
transform 1 0 9312 0 1 14364
box -48 -56 432 834
use sg13g2_nand2b_1  _0411_
timestamp 1676567195
transform -1 0 7776 0 1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _0412_
timestamp 1676557249
transform -1 0 10848 0 -1 15876
box -48 -56 432 834
use sg13g2_nand3_1  _0413_
timestamp 1683988354
transform 1 0 7776 0 1 12852
box -48 -56 528 834
use sg13g2_nand2b_1  _0414_
timestamp 1676567195
transform 1 0 10176 0 -1 12852
box -48 -56 528 834
use sg13g2_nor2b_1  _0415_
timestamp 1685181386
transform 1 0 9696 0 1 14364
box -54 -56 528 834
use sg13g2_mux4_1  _0416_
timestamp 1677257233
transform 1 0 13248 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0417_
timestamp 1677257233
transform 1 0 8352 0 -1 74844
box -48 -56 2064 834
use sg13g2_mux4_1  _0418_
timestamp 1677257233
transform -1 0 14976 0 1 50652
box -48 -56 2064 834
use sg13g2_mux4_1  _0419_
timestamp 1677257233
transform 1 0 7872 0 1 50652
box -48 -56 2064 834
use sg13g2_mux2_1  _0420_
timestamp 1677247768
transform 1 0 9216 0 1 35532
box -48 -56 1008 834
use sg13g2_nor2_1  _0421_
timestamp 1676627187
transform -1 0 12288 0 1 35532
box -48 -56 432 834
use sg13g2_nand2b_1  _0422_
timestamp 1676567195
transform -1 0 9984 0 -1 37044
box -48 -56 528 834
use sg13g2_nand2_1  _0423_
timestamp 1676557249
transform 1 0 9600 0 -1 38556
box -48 -56 432 834
use sg13g2_nand3_1  _0424_
timestamp 1683988354
transform -1 0 9792 0 1 37044
box -48 -56 528 834
use sg13g2_nand2b_1  _0425_
timestamp 1676567195
transform 1 0 9408 0 -1 34020
box -48 -56 528 834
use sg13g2_nor2b_1  _0426_
timestamp 1685181386
transform 1 0 7680 0 1 34020
box -54 -56 528 834
use sg13g2_mux4_1  _0427_
timestamp 1677257233
transform 1 0 6912 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0428_
timestamp 1677257233
transform 1 0 8352 0 1 73332
box -48 -56 2064 834
use sg13g2_mux4_1  _0429_
timestamp 1677257233
transform -1 0 8544 0 -1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0430_
timestamp 1677257233
transform 1 0 9600 0 -1 49140
box -48 -56 2064 834
use sg13g2_mux2_1  _0431_
timestamp 1677247768
transform 1 0 4416 0 1 15876
box -48 -56 1008 834
use sg13g2_nor2_1  _0432_
timestamp 1676627187
transform 1 0 4896 0 -1 18900
box -48 -56 432 834
use sg13g2_nand2b_1  _0433_
timestamp 1676567195
transform -1 0 5280 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _0434_
timestamp 1676557249
transform -1 0 6624 0 -1 18900
box -48 -56 432 834
use sg13g2_nand3_1  _0435_
timestamp 1683988354
transform 1 0 1728 0 1 17388
box -48 -56 528 834
use sg13g2_nand2b_1  _0436_
timestamp 1676567195
transform 1 0 5760 0 -1 18900
box -48 -56 528 834
use sg13g2_nor2b_1  _0437_
timestamp 1685181386
transform 1 0 5280 0 -1 18900
box -54 -56 528 834
use sg13g2_mux4_1  _0438_
timestamp 1677257233
transform 1 0 3744 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0439_
timestamp 1677257233
transform 1 0 5280 0 1 73332
box -48 -56 2064 834
use sg13g2_mux4_1  _0440_
timestamp 1677257233
transform 1 0 9408 0 1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0441_
timestamp 1677257233
transform 1 0 12960 0 -1 53676
box -48 -56 2064 834
use sg13g2_mux2_1  _0442_
timestamp 1677247768
transform 1 0 9984 0 1 9828
box -48 -56 1008 834
use sg13g2_nor2_1  _0443_
timestamp 1676627187
transform -1 0 11328 0 1 9828
box -48 -56 432 834
use sg13g2_nand2b_1  _0444_
timestamp 1676567195
transform -1 0 10272 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _0445_
timestamp 1676557249
transform 1 0 9120 0 -1 11340
box -48 -56 432 834
use sg13g2_nand3_1  _0446_
timestamp 1683988354
transform 1 0 9408 0 1 9828
box -48 -56 528 834
use sg13g2_nand2b_1  _0447_
timestamp 1676567195
transform 1 0 10656 0 1 8316
box -48 -56 528 834
use sg13g2_nor2b_1  _0448_
timestamp 1685181386
transform 1 0 10272 0 1 11340
box -54 -56 528 834
use sg13g2_mux4_1  _0449_
timestamp 1677257233
transform 1 0 11136 0 -1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0450_
timestamp 1677257233
transform 1 0 8256 0 1 76356
box -48 -56 2064 834
use sg13g2_mux4_1  _0451_
timestamp 1677257233
transform 1 0 12768 0 1 53676
box -48 -56 2064 834
use sg13g2_mux4_1  _0452_
timestamp 1677257233
transform 1 0 18240 0 1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0453_
timestamp 1677257233
transform 1 0 9504 0 1 41580
box -48 -56 2064 834
use sg13g2_mux4_1  _0454_
timestamp 1677257233
transform 1 0 10176 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0455_
timestamp 1677257233
transform 1 0 10272 0 1 76356
box -48 -56 2064 834
use sg13g2_mux4_1  _0456_
timestamp 1677257233
transform -1 0 20352 0 1 50652
box -48 -56 2064 834
use sg13g2_mux4_1  _0457_
timestamp 1677257233
transform 1 0 9984 0 1 46116
box -48 -56 2064 834
use sg13g2_mux4_1  _0458_
timestamp 1677257233
transform 1 0 8352 0 -1 41580
box -48 -56 2064 834
use sg13g2_mux4_1  _0459_
timestamp 1677257233
transform 1 0 7104 0 -1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _0460_
timestamp 1677257233
transform 1 0 8832 0 -1 71820
box -48 -56 2064 834
use sg13g2_mux4_1  _0461_
timestamp 1677257233
transform 1 0 10176 0 1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0462_
timestamp 1677257233
transform 1 0 8448 0 -1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0463_
timestamp 1677257233
transform 1 0 9216 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0464_
timestamp 1677257233
transform 1 0 6816 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _0465_
timestamp 1677257233
transform 1 0 8448 0 -1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0466_
timestamp 1677257233
transform -1 0 10560 0 1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0467_
timestamp 1677257233
transform 1 0 18048 0 -1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0468_
timestamp 1677257233
transform 1 0 9984 0 -1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0469_
timestamp 1677257233
transform 1 0 15264 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0470_
timestamp 1677257233
transform 1 0 10656 0 -1 79380
box -48 -56 2064 834
use sg13g2_mux4_1  _0471_
timestamp 1677257233
transform 1 0 18336 0 1 46116
box -48 -56 2064 834
use sg13g2_nand2b_1  _0472_
timestamp 1676567195
transform -1 0 12672 0 1 52164
box -48 -56 528 834
use sg13g2_nor3_1  _0473_
timestamp 1676639442
transform 1 0 12672 0 1 52164
box -48 -56 528 834
use sg13g2_a221oi_1  _0474_
timestamp 1685197497
transform 1 0 13152 0 1 52164
box -48 -56 816 834
use sg13g2_mux4_1  _0475_
timestamp 1677257233
transform 1 0 12672 0 1 46116
box -48 -56 2064 834
use sg13g2_nand2b_1  _0476_
timestamp 1676567195
transform 1 0 14880 0 1 9828
box -48 -56 528 834
use sg13g2_nor3_1  _0477_
timestamp 1676639442
transform 1 0 13536 0 -1 9828
box -48 -56 528 834
use sg13g2_a221oi_1  _0478_
timestamp 1685197497
transform 1 0 14208 0 -1 9828
box -48 -56 816 834
use sg13g2_mux4_1  _0479_
timestamp 1677257233
transform 1 0 12768 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _0480_
timestamp 1677257233
transform 1 0 11520 0 1 58212
box -48 -56 2064 834
use sg13g2_mux4_1  _0481_
timestamp 1677257233
transform 1 0 5088 0 1 58212
box -48 -56 2064 834
use sg13g2_mux4_1  _0482_
timestamp 1677257233
transform 1 0 2976 0 -1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0483_
timestamp 1677257233
transform 1 0 13056 0 1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0484_
timestamp 1677257233
transform 1 0 17280 0 -1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0485_
timestamp 1677257233
transform 1 0 9408 0 1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0486_
timestamp 1677257233
transform 1 0 10560 0 -1 61236
box -48 -56 2064 834
use sg13g2_mux4_1  _0487_
timestamp 1677257233
transform 1 0 15936 0 -1 61236
box -48 -56 2064 834
use sg13g2_mux4_1  _0488_
timestamp 1677257233
transform 1 0 17952 0 -1 61236
box -48 -56 2064 834
use sg13g2_mux4_1  _0489_
timestamp 1677257233
transform 1 0 10368 0 1 61236
box -48 -56 2064 834
use sg13g2_mux4_1  _0490_
timestamp 1677257233
transform 1 0 7392 0 -1 62748
box -48 -56 2064 834
use sg13g2_mux4_1  _0491_
timestamp 1677257233
transform 1 0 13728 0 -1 62748
box -48 -56 2064 834
use sg13g2_mux4_1  _0492_
timestamp 1677257233
transform 1 0 17376 0 1 62748
box -48 -56 2064 834
use sg13g2_mux4_1  _0493_
timestamp 1677257233
transform 1 0 7392 0 1 58212
box -48 -56 2064 834
use sg13g2_mux4_1  _0494_
timestamp 1677257233
transform 1 0 10656 0 -1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0495_
timestamp 1677257233
transform 1 0 13728 0 -1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0496_
timestamp 1677257233
transform 1 0 17280 0 -1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0497_
timestamp 1677257233
transform 1 0 10656 0 -1 65772
box -48 -56 2064 834
use sg13g2_mux4_1  _0498_
timestamp 1677257233
transform 1 0 7392 0 1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0499_
timestamp 1677257233
transform 1 0 13536 0 -1 65772
box -48 -56 2064 834
use sg13g2_mux4_1  _0500_
timestamp 1677257233
transform 1 0 16416 0 -1 65772
box -48 -56 2064 834
use sg13g2_mux4_1  _0501_
timestamp 1677257233
transform 1 0 9600 0 1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0502_
timestamp 1677257233
transform 1 0 6240 0 -1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0503_
timestamp 1677257233
transform 1 0 11232 0 1 73332
box -48 -56 2064 834
use sg13g2_mux4_1  _0504_
timestamp 1677257233
transform 1 0 13344 0 -1 67284
box -48 -56 2064 834
use sg13g2_mux4_1  _0505_
timestamp 1677257233
transform 1 0 12960 0 -1 79380
box -48 -56 2064 834
use sg13g2_mux4_1  _0506_
timestamp 1677257233
transform 1 0 16032 0 1 67284
box -48 -56 2064 834
use sg13g2_mux4_1  _0507_
timestamp 1677257233
transform 1 0 3264 0 -1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0508_
timestamp 1677257233
transform 1 0 7776 0 -1 67284
box -48 -56 2064 834
use sg13g2_mux4_1  _0509_
timestamp 1677257233
transform 1 0 3264 0 -1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0510_
timestamp 1677257233
transform 1 0 6144 0 -1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0511_
timestamp 1677257233
transform 1 0 12480 0 -1 74844
box -48 -56 2064 834
use sg13g2_mux4_1  _0512_
timestamp 1677257233
transform 1 0 17472 0 -1 70308
box -48 -56 2064 834
use sg13g2_mux4_1  _0513_
timestamp 1677257233
transform 1 0 14880 0 1 76356
box -48 -56 2064 834
use sg13g2_mux4_1  _0514_
timestamp 1677257233
transform 1 0 17472 0 -1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0515_
timestamp 1677257233
transform 1 0 2688 0 1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0516_
timestamp 1677257233
transform 1 0 9408 0 -1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0517_
timestamp 1677257233
transform 1 0 2688 0 1 62748
box -48 -56 2064 834
use sg13g2_mux4_1  _0518_
timestamp 1677257233
transform 1 0 6624 0 1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0519_
timestamp 1677257233
transform 1 0 11904 0 -1 73332
box -48 -56 2064 834
use sg13g2_mux4_1  _0520_
timestamp 1677257233
transform 1 0 15456 0 -1 70308
box -48 -56 2064 834
use sg13g2_mux4_1  _0521_
timestamp 1677257233
transform 1 0 14784 0 1 77868
box -48 -56 2064 834
use sg13g2_mux4_1  _0522_
timestamp 1677257233
transform 1 0 17280 0 1 65772
box -48 -56 2064 834
use sg13g2_mux4_1  _0523_
timestamp 1677257233
transform 1 0 3456 0 1 65772
box -48 -56 2064 834
use sg13g2_mux4_1  _0524_
timestamp 1677257233
transform 1 0 10464 0 -1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0525_
timestamp 1677257233
transform 1 0 2976 0 -1 61236
box -48 -56 2064 834
use sg13g2_mux4_1  _0526_
timestamp 1677257233
transform 1 0 5952 0 1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0527_
timestamp 1677257233
transform 1 0 11808 0 -1 71820
box -48 -56 2064 834
use sg13g2_mux4_1  _0528_
timestamp 1677257233
transform 1 0 13440 0 1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0529_
timestamp 1677257233
transform 1 0 13824 0 -1 71820
box -48 -56 2064 834
use sg13g2_mux4_1  _0530_
timestamp 1677257233
transform 1 0 5664 0 1 65772
box -48 -56 2064 834
use sg13g2_mux4_1  _0531_
timestamp 1677257233
transform 1 0 4416 0 -1 71820
box -48 -56 2064 834
use sg13g2_mux4_1  _0532_
timestamp 1677257233
transform 1 0 15072 0 -1 74844
box -48 -56 2064 834
use sg13g2_mux4_1  _0533_
timestamp 1677257233
transform 1 0 17376 0 -1 74844
box -48 -56 2064 834
use sg13g2_mux4_1  _0534_
timestamp 1677257233
transform 1 0 9504 0 1 67284
box -48 -56 2064 834
use sg13g2_mux4_1  _0535_
timestamp 1677257233
transform 1 0 6432 0 -1 71820
box -48 -56 2064 834
use sg13g2_mux4_1  _0536_
timestamp 1677257233
transform 1 0 16512 0 -1 73332
box -48 -56 2064 834
use sg13g2_mux4_1  _0537_
timestamp 1677257233
transform 1 0 17472 0 -1 76356
box -48 -56 2064 834
use sg13g2_mux4_1  _0538_
timestamp 1677257233
transform 1 0 9984 0 -1 70308
box -48 -56 2064 834
use sg13g2_mux4_1  _0539_
timestamp 1677257233
transform 1 0 7008 0 -1 61236
box -48 -56 2064 834
use sg13g2_mux4_1  _0540_
timestamp 1677257233
transform 1 0 16608 0 1 71820
box -48 -56 2064 834
use sg13g2_nand2b_1  _0541_
timestamp 1676567195
transform 1 0 16320 0 1 47628
box -48 -56 528 834
use sg13g2_o21ai_1  _0542_
timestamp 1685175443
transform -1 0 17760 0 -1 49140
box -48 -56 538 834
use sg13g2_o21ai_1  _0543_
timestamp 1685175443
transform 1 0 15360 0 1 49140
box -48 -56 538 834
use sg13g2_mux2_1  _0544_
timestamp 1677247768
transform 1 0 15840 0 1 49140
box -48 -56 1008 834
use sg13g2_a21oi_1  _0545_
timestamp 1683973020
transform 1 0 17280 0 1 50652
box -48 -56 528 834
use sg13g2_mux4_1  _0546_
timestamp 1677257233
transform 1 0 15264 0 -1 49140
box -48 -56 2064 834
use sg13g2_nor2_1  _0547_
timestamp 1676627187
transform -1 0 17472 0 -1 50652
box -48 -56 432 834
use sg13g2_nor2_1  _0548_
timestamp 1676627187
transform 1 0 14976 0 1 49140
box -48 -56 432 834
use sg13g2_nand2b_1  _0549_
timestamp 1676567195
transform 1 0 6912 0 1 47628
box -48 -56 528 834
use sg13g2_o21ai_1  _0550_
timestamp 1685175443
transform 1 0 7392 0 1 47628
box -48 -56 538 834
use sg13g2_o21ai_1  _0551_
timestamp 1685175443
transform 1 0 7584 0 -1 50652
box -48 -56 538 834
use sg13g2_mux2_1  _0552_
timestamp 1677247768
transform -1 0 8160 0 1 49140
box -48 -56 1008 834
use sg13g2_a21oi_1  _0553_
timestamp 1683973020
transform -1 0 6528 0 -1 52164
box -48 -56 528 834
use sg13g2_mux4_1  _0554_
timestamp 1677257233
transform 1 0 5568 0 -1 49140
box -48 -56 2064 834
use sg13g2_nor2_1  _0555_
timestamp 1676627187
transform -1 0 7968 0 -1 49140
box -48 -56 432 834
use sg13g2_nor2_1  _0556_
timestamp 1676627187
transform -1 0 8544 0 1 49140
box -48 -56 432 834
use sg13g2_nand2b_1  _0557_
timestamp 1676567195
transform 1 0 7296 0 -1 55188
box -48 -56 528 834
use sg13g2_o21ai_1  _0558_
timestamp 1685175443
transform 1 0 7296 0 1 56700
box -48 -56 538 834
use sg13g2_o21ai_1  _0559_
timestamp 1685175443
transform 1 0 8064 0 1 55188
box -48 -56 538 834
use sg13g2_mux2_1  _0560_
timestamp 1677247768
transform 1 0 7392 0 -1 56700
box -48 -56 1008 834
use sg13g2_a21oi_1  _0561_
timestamp 1683973020
transform 1 0 8352 0 -1 56700
box -48 -56 528 834
use sg13g2_mux4_1  _0562_
timestamp 1677257233
transform 1 0 6048 0 1 55188
box -48 -56 2064 834
use sg13g2_nor2_1  _0563_
timestamp 1676627187
transform -1 0 9216 0 -1 56700
box -48 -56 432 834
use sg13g2_nor2_1  _0564_
timestamp 1676627187
transform 1 0 6912 0 1 56700
box -48 -56 432 834
use sg13g2_nand2b_1  _0565_
timestamp 1676567195
transform 1 0 16800 0 -1 56700
box -48 -56 528 834
use sg13g2_o21ai_1  _0566_
timestamp 1685175443
transform 1 0 17472 0 -1 58212
box -48 -56 538 834
use sg13g2_o21ai_1  _0567_
timestamp 1685175443
transform 1 0 18912 0 -1 58212
box -48 -56 538 834
use sg13g2_mux2_1  _0568_
timestamp 1677247768
transform 1 0 17952 0 -1 58212
box -48 -56 1008 834
use sg13g2_a21oi_1  _0569_
timestamp 1683973020
transform 1 0 19872 0 1 56700
box -48 -56 528 834
use sg13g2_mux4_1  _0570_
timestamp 1677257233
transform 1 0 17760 0 -1 56700
box -48 -56 2064 834
use sg13g2_nor2_1  _0571_
timestamp 1676627187
transform 1 0 19392 0 -1 58212
box -48 -56 432 834
use sg13g2_nor2_1  _0572_
timestamp 1676627187
transform 1 0 17856 0 1 56700
box -48 -56 432 834
use sg13g2_nand2b_1  _0573_
timestamp 1676567195
transform -1 0 14880 0 -1 46116
box -48 -56 528 834
use sg13g2_o21ai_1  _0574_
timestamp 1685175443
transform 1 0 13056 0 1 43092
box -48 -56 538 834
use sg13g2_o21ai_1  _0575_
timestamp 1685175443
transform 1 0 14016 0 -1 44604
box -48 -56 538 834
use sg13g2_inv_1  _0576_
timestamp 1676382929
transform -1 0 11904 0 -1 44604
box -48 -56 336 834
use sg13g2_nand2b_1  _0577_
timestamp 1676567195
transform -1 0 14016 0 -1 44604
box -48 -56 528 834
use sg13g2_and2_1  _0578_
timestamp 1676901763
transform 1 0 13536 0 1 43092
box -48 -56 528 834
use sg13g2_o21ai_1  _0579_
timestamp 1685175443
transform 1 0 14016 0 1 43092
box -48 -56 538 834
use sg13g2_mux4_1  _0580_
timestamp 1677257233
transform 1 0 13152 0 1 44604
box -48 -56 2064 834
use sg13g2_nor2_1  _0581_
timestamp 1676627187
transform 1 0 15168 0 1 44604
box -48 -56 432 834
use sg13g2_a21oi_1  _0582_
timestamp 1683973020
transform 1 0 16512 0 1 43092
box -48 -56 528 834
use sg13g2_nand2b_1  _0583_
timestamp 1676567195
transform -1 0 6816 0 -1 47628
box -48 -56 528 834
use sg13g2_o21ai_1  _0584_
timestamp 1685175443
transform 1 0 6048 0 1 46116
box -48 -56 538 834
use sg13g2_o21ai_1  _0585_
timestamp 1685175443
transform 1 0 7008 0 1 46116
box -48 -56 538 834
use sg13g2_inv_1  _0586_
timestamp 1676382929
transform 1 0 8064 0 1 44604
box -48 -56 336 834
use sg13g2_nand2b_1  _0587_
timestamp 1676567195
transform -1 0 7968 0 1 46116
box -48 -56 528 834
use sg13g2_and2_1  _0588_
timestamp 1676901763
transform 1 0 6528 0 1 46116
box -48 -56 528 834
use sg13g2_o21ai_1  _0589_
timestamp 1685175443
transform 1 0 7104 0 1 44604
box -48 -56 538 834
use sg13g2_mux4_1  _0590_
timestamp 1677257233
transform 1 0 5664 0 -1 46116
box -48 -56 2064 834
use sg13g2_nor2_1  _0591_
timestamp 1676627187
transform -1 0 8352 0 1 46116
box -48 -56 432 834
use sg13g2_a21oi_1  _0592_
timestamp 1683973020
transform -1 0 8064 0 1 44604
box -48 -56 528 834
use sg13g2_nand2b_1  _0593_
timestamp 1676567195
transform 1 0 8448 0 -1 53676
box -48 -56 528 834
use sg13g2_o21ai_1  _0594_
timestamp 1685175443
transform -1 0 11040 0 1 52164
box -48 -56 538 834
use sg13g2_o21ai_1  _0595_
timestamp 1685175443
transform 1 0 10080 0 1 52164
box -48 -56 538 834
use sg13g2_inv_1  _0596_
timestamp 1676382929
transform 1 0 10848 0 1 53676
box -48 -56 336 834
use sg13g2_nand2b_1  _0597_
timestamp 1676567195
transform -1 0 8448 0 -1 53676
box -48 -56 528 834
use sg13g2_and2_1  _0598_
timestamp 1676901763
transform 1 0 11040 0 1 52164
box -48 -56 528 834
use sg13g2_o21ai_1  _0599_
timestamp 1685175443
transform 1 0 9984 0 -1 55188
box -48 -56 538 834
use sg13g2_mux4_1  _0600_
timestamp 1677257233
transform 1 0 8832 0 1 53676
box -48 -56 2064 834
use sg13g2_nor2_1  _0601_
timestamp 1676627187
transform -1 0 11904 0 1 52164
box -48 -56 432 834
use sg13g2_a21oi_1  _0602_
timestamp 1683973020
transform -1 0 11232 0 -1 53676
box -48 -56 528 834
use sg13g2_nand2b_1  _0603_
timestamp 1676567195
transform 1 0 17280 0 -1 56700
box -48 -56 528 834
use sg13g2_o21ai_1  _0604_
timestamp 1685175443
transform 1 0 15456 0 1 53676
box -48 -56 538 834
use sg13g2_o21ai_1  _0605_
timestamp 1685175443
transform -1 0 17280 0 -1 53676
box -48 -56 538 834
use sg13g2_inv_1  _0606_
timestamp 1676382929
transform -1 0 16032 0 -1 52164
box -48 -56 336 834
use sg13g2_nand2b_1  _0607_
timestamp 1676567195
transform 1 0 17568 0 1 55188
box -48 -56 528 834
use sg13g2_and2_1  _0608_
timestamp 1676901763
transform 1 0 17760 0 -1 55188
box -48 -56 528 834
use sg13g2_o21ai_1  _0609_
timestamp 1685175443
transform -1 0 17760 0 -1 55188
box -48 -56 538 834
use sg13g2_mux4_1  _0610_
timestamp 1677257233
transform -1 0 17952 0 1 53676
box -48 -56 2064 834
use sg13g2_nor2_1  _0611_
timestamp 1676627187
transform 1 0 15072 0 1 53676
box -48 -56 432 834
use sg13g2_a21oi_1  _0612_
timestamp 1683973020
transform 1 0 16608 0 -1 55188
box -48 -56 528 834
use sg13g2_mux4_1  _0613_
timestamp 1677257233
transform 1 0 12096 0 -1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0614_
timestamp 1677257233
transform 1 0 3552 0 -1 41580
box -48 -56 2064 834
use sg13g2_mux4_1  _0615_
timestamp 1677257233
transform 1 0 2304 0 1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0616_
timestamp 1677257233
transform 1 0 12288 0 -1 40068
box -48 -56 2064 834
use sg13g2_a21oi_1  _0617_
timestamp 1683973020
transform 1 0 19104 0 -1 50652
box -48 -56 528 834
use sg13g2_o21ai_1  _0618_
timestamp 1685175443
transform 1 0 19584 0 -1 50652
box -48 -56 538 834
use sg13g2_mux4_1  _0619_
timestamp 1677257233
transform -1 0 19776 0 -1 49140
box -48 -56 2064 834
use sg13g2_nor2_1  _0620_
timestamp 1676627187
transform -1 0 18144 0 1 52164
box -48 -56 432 834
use sg13g2_a21oi_1  _0621_
timestamp 1683973020
transform 1 0 19776 0 -1 49140
box -48 -56 528 834
use sg13g2_a21oi_1  _0622_
timestamp 1683973020
transform -1 0 3552 0 -1 49140
box -48 -56 528 834
use sg13g2_o21ai_1  _0623_
timestamp 1685175443
transform -1 0 5088 0 1 49140
box -48 -56 538 834
use sg13g2_mux4_1  _0624_
timestamp 1677257233
transform -1 0 5568 0 -1 49140
box -48 -56 2064 834
use sg13g2_nor2_1  _0625_
timestamp 1676627187
transform 1 0 2784 0 1 47628
box -48 -56 432 834
use sg13g2_a21oi_1  _0626_
timestamp 1683973020
transform 1 0 2400 0 -1 47628
box -48 -56 528 834
use sg13g2_a21oi_1  _0627_
timestamp 1683973020
transform 1 0 6144 0 1 52164
box -48 -56 528 834
use sg13g2_o21ai_1  _0628_
timestamp 1685175443
transform 1 0 4992 0 1 53676
box -48 -56 538 834
use sg13g2_mux4_1  _0629_
timestamp 1677257233
transform -1 0 7968 0 -1 53676
box -48 -56 2064 834
use sg13g2_nor2_1  _0630_
timestamp 1676627187
transform 1 0 5760 0 1 52164
box -48 -56 432 834
use sg13g2_a21oi_1  _0631_
timestamp 1683973020
transform -1 0 6048 0 -1 52164
box -48 -56 528 834
use sg13g2_a21oi_1  _0632_
timestamp 1683973020
transform 1 0 19776 0 -1 56700
box -48 -56 528 834
use sg13g2_o21ai_1  _0633_
timestamp 1685175443
transform -1 0 20256 0 1 52164
box -48 -56 538 834
use sg13g2_mux4_1  _0634_
timestamp 1677257233
transform -1 0 20160 0 1 53676
box -48 -56 2064 834
use sg13g2_nor2_1  _0635_
timestamp 1676627187
transform 1 0 16416 0 1 52164
box -48 -56 432 834
use sg13g2_a21oi_1  _0636_
timestamp 1683973020
transform 1 0 19584 0 -1 53676
box -48 -56 528 834
use sg13g2_nor2b_1  _0637_
timestamp 1685181386
transform 1 0 17376 0 -1 46116
box -54 -56 528 834
use sg13g2_o21ai_1  _0638_
timestamp 1685175443
transform 1 0 16896 0 1 46116
box -48 -56 538 834
use sg13g2_mux4_1  _0639_
timestamp 1677257233
transform 1 0 15360 0 -1 46116
box -48 -56 2064 834
use sg13g2_nor2b_1  _0640_
timestamp 1685181386
transform -1 0 17568 0 -1 44604
box -54 -56 528 834
use sg13g2_nor3_1  _0641_
timestamp 1676639442
transform -1 0 18336 0 -1 46116
box -48 -56 528 834
use sg13g2_or2_1  _0642_
timestamp 1684236171
transform -1 0 16992 0 -1 44604
box -48 -56 528 834
use sg13g2_nor2b_1  _0643_
timestamp 1685181386
transform -1 0 4992 0 -1 47628
box -54 -56 528 834
use sg13g2_o21ai_1  _0644_
timestamp 1685175443
transform -1 0 5280 0 1 46116
box -48 -56 538 834
use sg13g2_mux4_1  _0645_
timestamp 1677257233
transform -1 0 5280 0 -1 46116
box -48 -56 2064 834
use sg13g2_nor2b_1  _0646_
timestamp 1685181386
transform 1 0 4608 0 1 44604
box -54 -56 528 834
use sg13g2_nor3_1  _0647_
timestamp 1676639442
transform 1 0 3648 0 1 44604
box -48 -56 528 834
use sg13g2_or2_1  _0648_
timestamp 1684236171
transform -1 0 4608 0 1 44604
box -48 -56 528 834
use sg13g2_nor2b_1  _0649_
timestamp 1685181386
transform 1 0 3264 0 1 50652
box -54 -56 528 834
use sg13g2_o21ai_1  _0650_
timestamp 1685175443
transform -1 0 4224 0 1 50652
box -48 -56 538 834
use sg13g2_mux4_1  _0651_
timestamp 1677257233
transform -1 0 4992 0 -1 52164
box -48 -56 2064 834
use sg13g2_nor2b_1  _0652_
timestamp 1685181386
transform 1 0 2976 0 1 52164
box -54 -56 528 834
use sg13g2_nor3_1  _0653_
timestamp 1676639442
transform 1 0 3456 0 1 52164
box -48 -56 528 834
use sg13g2_or2_1  _0654_
timestamp 1684236171
transform -1 0 3264 0 1 50652
box -48 -56 528 834
use sg13g2_nor2b_1  _0655_
timestamp 1685181386
transform 1 0 16800 0 1 52164
box -54 -56 528 834
use sg13g2_o21ai_1  _0656_
timestamp 1685175443
transform 1 0 17472 0 -1 53676
box -48 -56 538 834
use sg13g2_mux4_1  _0657_
timestamp 1677257233
transform 1 0 16032 0 -1 52164
box -48 -56 2064 834
use sg13g2_nor2b_1  _0658_
timestamp 1685181386
transform -1 0 18528 0 -1 52164
box -54 -56 528 834
use sg13g2_nor3_1  _0659_
timestamp 1676639442
transform 1 0 17280 0 1 52164
box -48 -56 528 834
use sg13g2_or2_1  _0660_
timestamp 1684236171
transform -1 0 18240 0 1 50652
box -48 -56 528 834
use sg13g2_mux4_1  _0661_
timestamp 1677257233
transform 1 0 12384 0 1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0662_
timestamp 1677257233
transform 1 0 13152 0 -1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0663_
timestamp 1677257233
transform 1 0 5664 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0664_
timestamp 1677257233
transform 1 0 4416 0 -1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0665_
timestamp 1677257233
transform 1 0 12480 0 1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0666_
timestamp 1677257233
transform 1 0 13248 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0667_
timestamp 1677257233
transform 1 0 7392 0 -1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0668_
timestamp 1677257233
transform 1 0 6720 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0669_
timestamp 1677257233
transform 1 0 10656 0 -1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _0670_
timestamp 1677257233
transform 1 0 10848 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0671_
timestamp 1677257233
transform 1 0 8064 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0672_
timestamp 1677257233
transform 1 0 8544 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0673_
timestamp 1677257233
transform 1 0 12480 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0674_
timestamp 1677257233
transform 1 0 12864 0 -1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0675_
timestamp 1677257233
transform 1 0 2208 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0676_
timestamp 1677257233
transform 1 0 2208 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0677_
timestamp 1677257233
transform 1 0 14784 0 -1 18900
box -48 -56 2064 834
use sg13g2_nand2b_1  _0678_
timestamp 1676567195
transform 1 0 19680 0 1 15876
box -48 -56 528 834
use sg13g2_nor3_1  _0679_
timestamp 1676639442
transform 1 0 18432 0 1 15876
box -48 -56 528 834
use sg13g2_a221oi_1  _0680_
timestamp 1685197497
transform 1 0 18912 0 1 15876
box -48 -56 816 834
use sg13g2_nand2b_1  _0681_
timestamp 1676567195
transform 1 0 9600 0 1 17388
box -48 -56 528 834
use sg13g2_nor3_1  _0682_
timestamp 1676639442
transform 1 0 9120 0 1 17388
box -48 -56 528 834
use sg13g2_a221oi_1  _0683_
timestamp 1685197497
transform 1 0 10560 0 1 17388
box -48 -56 816 834
use sg13g2_nand2b_1  _0684_
timestamp 1676567195
transform 1 0 12768 0 1 15876
box -48 -56 528 834
use sg13g2_nor3_1  _0685_
timestamp 1676639442
transform -1 0 14208 0 1 17388
box -48 -56 528 834
use sg13g2_a221oi_1  _0686_
timestamp 1685197497
transform -1 0 13728 0 1 17388
box -48 -56 816 834
use sg13g2_nand2b_1  _0687_
timestamp 1676567195
transform -1 0 19872 0 1 5292
box -48 -56 528 834
use sg13g2_nor3_1  _0688_
timestamp 1676639442
transform 1 0 18912 0 1 6804
box -48 -56 528 834
use sg13g2_a221oi_1  _0689_
timestamp 1685197497
transform 1 0 19200 0 1 8316
box -48 -56 816 834
use sg13g2_nand2b_1  _0690_
timestamp 1676567195
transform -1 0 19968 0 1 6804
box -48 -56 528 834
use sg13g2_nor3_1  _0691_
timestamp 1676639442
transform -1 0 20352 0 -1 8316
box -48 -56 528 834
use sg13g2_a221oi_1  _0692_
timestamp 1685197497
transform -1 0 19968 0 -1 9828
box -48 -56 816 834
use sg13g2_nand2b_1  _0693_
timestamp 1676567195
transform 1 0 9024 0 -1 20412
box -48 -56 528 834
use sg13g2_nor3_1  _0694_
timestamp 1676639442
transform 1 0 7776 0 -1 20412
box -48 -56 528 834
use sg13g2_a221oi_1  _0695_
timestamp 1685197497
transform 1 0 8256 0 -1 20412
box -48 -56 816 834
use sg13g2_nand2b_1  _0696_
timestamp 1676567195
transform 1 0 11904 0 1 20412
box -48 -56 528 834
use sg13g2_nor3_1  _0697_
timestamp 1676639442
transform -1 0 11712 0 -1 20412
box -48 -56 528 834
use sg13g2_a221oi_1  _0698_
timestamp 1685197497
transform 1 0 11136 0 1 20412
box -48 -56 816 834
use sg13g2_nand2b_1  _0699_
timestamp 1676567195
transform 1 0 19008 0 -1 18900
box -48 -56 528 834
use sg13g2_nor3_1  _0700_
timestamp 1676639442
transform -1 0 20064 0 1 18900
box -48 -56 528 834
use sg13g2_a221oi_1  _0701_
timestamp 1685197497
transform -1 0 19776 0 -1 20412
box -48 -56 816 834
use sg13g2_nand2b_1  _0702_
timestamp 1676567195
transform 1 0 19680 0 1 17388
box -48 -56 528 834
use sg13g2_nor3_1  _0703_
timestamp 1676639442
transform -1 0 19968 0 -1 18900
box -48 -56 528 834
use sg13g2_a221oi_1  _0704_
timestamp 1685197497
transform -1 0 19680 0 1 17388
box -48 -56 816 834
use sg13g2_nand2b_1  _0705_
timestamp 1676567195
transform 1 0 10464 0 -1 18900
box -48 -56 528 834
use sg13g2_nor3_1  _0706_
timestamp 1676639442
transform 1 0 10080 0 1 17388
box -48 -56 528 834
use sg13g2_a221oi_1  _0707_
timestamp 1685197497
transform 1 0 10464 0 1 18900
box -48 -56 816 834
use sg13g2_nand2b_1  _0708_
timestamp 1676567195
transform 1 0 14016 0 1 18900
box -48 -56 528 834
use sg13g2_nor3_1  _0709_
timestamp 1676639442
transform 1 0 12576 0 1 20412
box -48 -56 528 834
use sg13g2_a221oi_1  _0710_
timestamp 1685197497
transform 1 0 13248 0 1 18900
box -48 -56 816 834
use sg13g2_nand2b_1  _0711_
timestamp 1676567195
transform -1 0 15552 0 1 20412
box -48 -56 528 834
use sg13g2_nor3_1  _0712_
timestamp 1676639442
transform -1 0 17568 0 -1 21924
box -48 -56 528 834
use sg13g2_a221oi_1  _0713_
timestamp 1685197497
transform -1 0 16608 0 1 21924
box -48 -56 816 834
use sg13g2_nand2b_1  _0714_
timestamp 1676567195
transform -1 0 19680 0 -1 21924
box -48 -56 528 834
use sg13g2_nor3_1  _0715_
timestamp 1676639442
transform -1 0 20256 0 -1 21924
box -48 -56 528 834
use sg13g2_a221oi_1  _0716_
timestamp 1685197497
transform -1 0 19776 0 -1 23436
box -48 -56 816 834
use sg13g2_nand2b_1  _0717_
timestamp 1676567195
transform 1 0 9600 0 -1 21924
box -48 -56 528 834
use sg13g2_nor3_1  _0718_
timestamp 1676639442
transform 1 0 8640 0 -1 23436
box -48 -56 528 834
use sg13g2_a221oi_1  _0719_
timestamp 1685197497
transform 1 0 9696 0 1 21924
box -48 -56 816 834
use sg13g2_nand2b_1  _0720_
timestamp 1676567195
transform 1 0 10944 0 -1 21924
box -48 -56 528 834
use sg13g2_nor3_1  _0721_
timestamp 1676639442
transform 1 0 9120 0 -1 23436
box -48 -56 528 834
use sg13g2_a221oi_1  _0722_
timestamp 1685197497
transform 1 0 11136 0 1 23436
box -48 -56 816 834
use sg13g2_nand2b_1  _0723_
timestamp 1676567195
transform -1 0 17376 0 -1 18900
box -48 -56 528 834
use sg13g2_nor3_1  _0724_
timestamp 1676639442
transform -1 0 20256 0 -1 20412
box -48 -56 528 834
use sg13g2_a221oi_1  _0725_
timestamp 1685197497
transform -1 0 18624 0 1 20412
box -48 -56 816 834
use sg13g2_mux4_1  _0726_
timestamp 1677257233
transform 1 0 17376 0 1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0727_
timestamp 1677257233
transform 1 0 7680 0 -1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0728_
timestamp 1677257233
transform 1 0 10080 0 -1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0729_
timestamp 1677257233
transform 1 0 17088 0 1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0730_
timestamp 1677257233
transform 1 0 12096 0 1 41580
box -48 -56 2064 834
use sg13g2_mux4_1  _0731_
timestamp 1677257233
transform 1 0 14112 0 1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0732_
timestamp 1677257233
transform 1 0 2784 0 -1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0733_
timestamp 1677257233
transform 1 0 6816 0 1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0734_
timestamp 1677257233
transform 1 0 4032 0 1 41580
box -48 -56 2064 834
use sg13g2_mux4_1  _0735_
timestamp 1677257233
transform 1 0 10464 0 -1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0736_
timestamp 1677257233
transform 1 0 14208 0 1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0737_
timestamp 1677257233
transform 1 0 16320 0 -1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0738_
timestamp 1677257233
transform 1 0 14208 0 -1 41580
box -48 -56 2064 834
use sg13g2_mux4_1  _0739_
timestamp 1677257233
transform -1 0 19392 0 -1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0740_
timestamp 1677257233
transform 1 0 2400 0 -1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _0741_
timestamp 1677257233
transform 1 0 7584 0 1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0742_
timestamp 1677257233
transform 1 0 2976 0 -1 43092
box -48 -56 2064 834
use sg13g2_mux4_1  _0743_
timestamp 1677257233
transform 1 0 9984 0 -1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0744_
timestamp 1677257233
transform 1 0 13056 0 -1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0745_
timestamp 1677257233
transform 1 0 17472 0 1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0746_
timestamp 1677257233
transform 1 0 14208 0 1 41580
box -48 -56 2064 834
use sg13g2_mux4_1  _0747_
timestamp 1677257233
transform 1 0 13056 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0748_
timestamp 1677257233
transform 1 0 2784 0 1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _0749_
timestamp 1677257233
transform 1 0 6624 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0750_
timestamp 1677257233
transform 1 0 3648 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0751_
timestamp 1677257233
transform 1 0 10464 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0752_
timestamp 1677257233
transform 1 0 15072 0 -1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0753_
timestamp 1677257233
transform 1 0 17088 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0754_
timestamp 1677257233
transform 1 0 15168 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0755_
timestamp 1677257233
transform 1 0 6240 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0756_
timestamp 1677257233
transform 1 0 6048 0 -1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0757_
timestamp 1677257233
transform 1 0 14208 0 1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0758_
timestamp 1677257233
transform 1 0 16512 0 1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0759_
timestamp 1677257233
transform 1 0 7008 0 -1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0760_
timestamp 1677257233
transform 1 0 7488 0 -1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0761_
timestamp 1677257233
transform 1 0 15072 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0762_
timestamp 1677257233
transform 1 0 14304 0 1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0763_
timestamp 1677257233
transform 1 0 7296 0 1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0764_
timestamp 1677257233
transform 1 0 9888 0 1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0765_
timestamp 1677257233
transform 1 0 17472 0 1 35532
box -48 -56 2064 834
use sg13g2_mux2_1  _0766_
timestamp 1677247768
transform 1 0 15744 0 -1 11340
box -48 -56 1008 834
use sg13g2_nand2b_1  _0767_
timestamp 1676567195
transform 1 0 17568 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _0768_
timestamp 1685175443
transform 1 0 17088 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _0769_
timestamp 1683973020
transform -1 0 17184 0 -1 11340
box -48 -56 528 834
use sg13g2_nor2b_1  _0770_
timestamp 1685181386
transform -1 0 18336 0 1 11340
box -54 -56 528 834
use sg13g2_mux4_1  _0771_
timestamp 1677257233
transform -1 0 17280 0 -1 12852
box -48 -56 2064 834
use sg13g2_nor2_1  _0772_
timestamp 1676627187
transform -1 0 15744 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _0773_
timestamp 1683973020
transform -1 0 15264 0 -1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _0774_
timestamp 1677247768
transform 1 0 7680 0 -1 35532
box -48 -56 1008 834
use sg13g2_nand2b_1  _0775_
timestamp 1676567195
transform 1 0 7680 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _0776_
timestamp 1685175443
transform -1 0 5664 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  _0777_
timestamp 1683973020
transform 1 0 5184 0 -1 35532
box -48 -56 528 834
use sg13g2_nor2b_1  _0778_
timestamp 1685181386
transform 1 0 4704 0 -1 35532
box -54 -56 528 834
use sg13g2_mux4_1  _0779_
timestamp 1677257233
transform 1 0 5664 0 -1 35532
box -48 -56 2064 834
use sg13g2_nor2_1  _0780_
timestamp 1676627187
transform -1 0 8448 0 -1 38556
box -48 -56 432 834
use sg13g2_a21oi_1  _0781_
timestamp 1683973020
transform -1 0 7296 0 1 35532
box -48 -56 528 834
use sg13g2_mux2_1  _0782_
timestamp 1677247768
transform 1 0 5280 0 -1 27972
box -48 -56 1008 834
use sg13g2_nand2b_1  _0783_
timestamp 1676567195
transform 1 0 5760 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _0784_
timestamp 1685175443
transform -1 0 1632 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _0785_
timestamp 1683973020
transform 1 0 4512 0 1 23436
box -48 -56 528 834
use sg13g2_nor2b_1  _0786_
timestamp 1685181386
transform 1 0 5280 0 1 26460
box -54 -56 528 834
use sg13g2_mux4_1  _0787_
timestamp 1677257233
transform -1 0 5760 0 1 24948
box -48 -56 2064 834
use sg13g2_nor2_1  _0788_
timestamp 1676627187
transform 1 0 3264 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _0789_
timestamp 1683973020
transform -1 0 6720 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _0790_
timestamp 1677247768
transform 1 0 14304 0 -1 29484
box -48 -56 1008 834
use sg13g2_nand2b_1  _0791_
timestamp 1676567195
transform 1 0 14688 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _0792_
timestamp 1685175443
transform -1 0 14208 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _0793_
timestamp 1683973020
transform 1 0 16416 0 -1 27972
box -48 -56 528 834
use sg13g2_nor2b_1  _0794_
timestamp 1685181386
transform 1 0 11808 0 1 27972
box -54 -56 528 834
use sg13g2_mux4_1  _0795_
timestamp 1677257233
transform 1 0 12672 0 1 26460
box -48 -56 2064 834
use sg13g2_nor2_1  _0796_
timestamp 1676627187
transform -1 0 16224 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _0797_
timestamp 1683973020
transform -1 0 14112 0 1 29484
box -48 -56 528 834
use sg13g2_mux2_1  _0798_
timestamp 1677247768
transform 1 0 15072 0 1 12852
box -48 -56 1008 834
use sg13g2_nand2b_1  _0799_
timestamp 1676567195
transform 1 0 17664 0 -1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _0800_
timestamp 1677247768
transform 1 0 16032 0 1 12852
box -48 -56 1008 834
use sg13g2_a21oi_1  _0801_
timestamp 1683973020
transform -1 0 17376 0 1 14364
box -48 -56 528 834
use sg13g2_mux4_1  _0802_
timestamp 1677257233
transform 1 0 15648 0 -1 14364
box -48 -56 2064 834
use sg13g2_nor2_1  _0803_
timestamp 1676627187
transform -1 0 18336 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _0804_
timestamp 1683973020
transform -1 0 17568 0 -1 15876
box -48 -56 528 834
use sg13g2_mux2_1  _0805_
timestamp 1677247768
transform 1 0 9216 0 -1 35532
box -48 -56 1008 834
use sg13g2_nand2b_1  _0806_
timestamp 1676567195
transform 1 0 12384 0 -1 32508
box -48 -56 528 834
use sg13g2_mux2_1  _0807_
timestamp 1677247768
transform 1 0 10464 0 -1 37044
box -48 -56 1008 834
use sg13g2_a21oi_1  _0808_
timestamp 1683973020
transform 1 0 12096 0 -1 35532
box -48 -56 528 834
use sg13g2_mux4_1  _0809_
timestamp 1677257233
transform 1 0 10080 0 1 34020
box -48 -56 2064 834
use sg13g2_nor2_1  _0810_
timestamp 1676627187
transform -1 0 12768 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _0811_
timestamp 1683973020
transform -1 0 12576 0 1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _0812_
timestamp 1677247768
transform 1 0 6336 0 -1 23436
box -48 -56 1008 834
use sg13g2_nand2b_1  _0813_
timestamp 1676567195
transform -1 0 8064 0 1 21924
box -48 -56 528 834
use sg13g2_mux2_1  _0814_
timestamp 1677247768
transform 1 0 7008 0 -1 21924
box -48 -56 1008 834
use sg13g2_a21oi_1  _0815_
timestamp 1683973020
transform 1 0 7872 0 -1 23436
box -48 -56 528 834
use sg13g2_mux4_1  _0816_
timestamp 1677257233
transform -1 0 7584 0 1 21924
box -48 -56 2064 834
use sg13g2_nor2_1  _0817_
timestamp 1676627187
transform 1 0 5184 0 1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _0818_
timestamp 1683973020
transform 1 0 7392 0 -1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _0819_
timestamp 1677247768
transform 1 0 16128 0 1 26460
box -48 -56 1008 834
use sg13g2_nand2b_1  _0820_
timestamp 1676567195
transform 1 0 18816 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _0821_
timestamp 1677247768
transform 1 0 16416 0 -1 23436
box -48 -56 1008 834
use sg13g2_a21oi_1  _0822_
timestamp 1683973020
transform 1 0 17856 0 -1 24948
box -48 -56 528 834
use sg13g2_mux4_1  _0823_
timestamp 1677257233
transform 1 0 15840 0 -1 24948
box -48 -56 2064 834
use sg13g2_nor2_1  _0824_
timestamp 1676627187
transform 1 0 17472 0 1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _0825_
timestamp 1683973020
transform -1 0 16320 0 -1 23436
box -48 -56 528 834
use sg13g2_nor2_1  _0826_
timestamp 1676627187
transform -1 0 20352 0 -1 9828
box -48 -56 432 834
use sg13g2_nor2b_1  _0827_
timestamp 1685181386
transform -1 0 18624 0 1 9828
box -54 -56 528 834
use sg13g2_mux4_1  _0828_
timestamp 1677257233
transform 1 0 18336 0 -1 12852
box -48 -56 2064 834
use sg13g2_nor3_1  _0829_
timestamp 1676639442
transform -1 0 19776 0 1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _0830_
timestamp 1677247768
transform -1 0 19968 0 1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  _0831_
timestamp 1677247768
transform 1 0 4608 0 1 30996
box -48 -56 1008 834
use sg13g2_nand3b_1  _0832_
timestamp 1676573470
transform 1 0 5664 0 1 29484
box -48 -56 720 834
use sg13g2_mux4_1  _0833_
timestamp 1677257233
transform 1 0 4896 0 -1 30996
box -48 -56 2064 834
use sg13g2_inv_1  _0834_
timestamp 1676382929
transform -1 0 6624 0 1 29484
box -48 -56 336 834
use sg13g2_o21ai_1  _0835_
timestamp 1685175443
transform 1 0 6912 0 -1 30996
box -48 -56 538 834
use sg13g2_nor2b_1  _0836_
timestamp 1685181386
transform 1 0 3744 0 -1 23436
box -54 -56 528 834
use sg13g2_nor2_1  _0837_
timestamp 1676627187
transform 1 0 1248 0 -1 24948
box -48 -56 432 834
use sg13g2_mux4_1  _0838_
timestamp 1677257233
transform -1 0 5664 0 -1 24948
box -48 -56 2064 834
use sg13g2_nor3_1  _0839_
timestamp 1676639442
transform 1 0 1152 0 1 24948
box -48 -56 528 834
use sg13g2_mux2_1  _0840_
timestamp 1677247768
transform -1 0 4512 0 1 23436
box -48 -56 1008 834
use sg13g2_nor2_1  _0841_
timestamp 1676627187
transform 1 0 13344 0 -1 26460
box -48 -56 432 834
use sg13g2_nor2b_1  _0842_
timestamp 1685181386
transform 1 0 14208 0 -1 24948
box -54 -56 528 834
use sg13g2_mux4_1  _0843_
timestamp 1677257233
transform -1 0 13728 0 1 24948
box -48 -56 2064 834
use sg13g2_nor3_1  _0844_
timestamp 1676639442
transform 1 0 13152 0 -1 24948
box -48 -56 528 834
use sg13g2_mux2_1  _0845_
timestamp 1677247768
transform -1 0 13344 0 -1 26460
box -48 -56 1008 834
use sg13g2_mux4_1  _0846_
timestamp 1677257233
transform 1 0 18240 0 -1 11340
box -48 -56 2064 834
use sg13g2_nand2b_1  _0847_
timestamp 1676567195
transform 1 0 19392 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2b_1  _0848_
timestamp 1676567195
transform -1 0 18144 0 -1 11340
box -48 -56 528 834
use sg13g2_nand2b_1  _0849_
timestamp 1676567195
transform 1 0 16800 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _0850_
timestamp 1685175443
transform -1 0 18144 0 1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _0851_
timestamp 1685175443
transform -1 0 17664 0 -1 11340
box -48 -56 538 834
use sg13g2_mux4_1  _0852_
timestamp 1677257233
transform 1 0 2880 0 1 27972
box -48 -56 2064 834
use sg13g2_nand2b_1  _0853_
timestamp 1676567195
transform 1 0 4416 0 -1 29484
box -48 -56 528 834
use sg13g2_nand2b_1  _0854_
timestamp 1676567195
transform -1 0 2400 0 -1 29484
box -48 -56 528 834
use sg13g2_nand2b_1  _0855_
timestamp 1676567195
transform -1 0 5376 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _0856_
timestamp 1685175443
transform -1 0 4032 0 1 29484
box -48 -56 538 834
use sg13g2_o21ai_1  _0857_
timestamp 1685175443
transform -1 0 1632 0 1 26460
box -48 -56 538 834
use sg13g2_nand2b_1  _0858_
timestamp 1676567195
transform 1 0 4320 0 -1 21924
box -48 -56 528 834
use sg13g2_nand2b_1  _0859_
timestamp 1676567195
transform -1 0 3840 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _0860_
timestamp 1685175443
transform 1 0 3264 0 -1 23436
box -48 -56 538 834
use sg13g2_mux4_1  _0861_
timestamp 1677257233
transform 1 0 2880 0 1 21924
box -48 -56 2064 834
use sg13g2_nand2b_1  _0862_
timestamp 1676567195
transform 1 0 4992 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _0863_
timestamp 1685175443
transform -1 0 4320 0 -1 21924
box -48 -56 538 834
use sg13g2_mux4_1  _0864_
timestamp 1677257233
transform 1 0 18336 0 -1 24948
box -48 -56 2064 834
use sg13g2_nand2b_1  _0865_
timestamp 1676567195
transform -1 0 20160 0 1 23436
box -48 -56 528 834
use sg13g2_nand2b_1  _0866_
timestamp 1676567195
transform 1 0 19776 0 -1 23436
box -48 -56 528 834
use sg13g2_nand2b_1  _0867_
timestamp 1676567195
transform 1 0 19680 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _0868_
timestamp 1685175443
transform 1 0 19200 0 1 24948
box -48 -56 538 834
use sg13g2_o21ai_1  _0869_
timestamp 1685175443
transform -1 0 20160 0 -1 26460
box -48 -56 538 834
use sg13g2_nor2b_1  _0870_
timestamp 1685181386
transform -1 0 6528 0 -1 12852
box -54 -56 528 834
use sg13g2_nor2_1  _0871_
timestamp 1676627187
transform -1 0 7200 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _0872_
timestamp 1683973020
transform -1 0 6048 0 -1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _0873_
timestamp 1677247768
transform -1 0 4512 0 1 12852
box -48 -56 1008 834
use sg13g2_nor3_1  _0874_
timestamp 1676639442
transform -1 0 4032 0 1 11340
box -48 -56 528 834
use sg13g2_mux4_1  _0875_
timestamp 1677257233
transform 1 0 4992 0 1 12852
box -48 -56 2064 834
use sg13g2_inv_1  _0876_
timestamp 1676382929
transform 1 0 7008 0 1 12852
box -48 -56 336 834
use sg13g2_a221oi_1  _0877_
timestamp 1685197497
transform 1 0 4800 0 -1 14364
box -48 -56 816 834
use sg13g2_nor3_1  _0878_
timestamp 1676639442
transform 1 0 5568 0 1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _0879_
timestamp 1677247768
transform -1 0 5472 0 -1 12852
box -48 -56 1008 834
use sg13g2_o21ai_1  _0880_
timestamp 1685175443
transform 1 0 3264 0 -1 12852
box -48 -56 538 834
use sg13g2_nand2b_1  _0881_
timestamp 1676567195
transform -1 0 6240 0 -1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _0882_
timestamp 1685173987
transform 1 0 3936 0 -1 14364
box -48 -56 624 834
use sg13g2_nor3_1  _0883_
timestamp 1676639442
transform 1 0 3456 0 1 14364
box -48 -56 528 834
use sg13g2_nor3_1  _0884_
timestamp 1676639442
transform -1 0 4512 0 1 11340
box -48 -56 528 834
use sg13g2_nor2b_1  _0885_
timestamp 1685181386
transform 1 0 2976 0 1 14364
box -54 -56 528 834
use sg13g2_o21ai_1  _0886_
timestamp 1685175443
transform -1 0 3936 0 -1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _0887_
timestamp 1685175443
transform -1 0 4224 0 -1 12852
box -48 -56 538 834
use sg13g2_inv_1  _0888_
timestamp 1676382929
transform -1 0 3072 0 -1 34020
box -48 -56 336 834
use sg13g2_nor2b_1  _0889_
timestamp 1685181386
transform 1 0 4128 0 1 6804
box -54 -56 528 834
use sg13g2_nor2b_1  _0890_
timestamp 1685181386
transform -1 0 5952 0 -1 9828
box -54 -56 528 834
use sg13g2_nor2b_1  _0891_
timestamp 1685181386
transform -1 0 4800 0 1 8316
box -54 -56 528 834
use sg13g2_nand2_1  _0892_
timestamp 1676557249
transform 1 0 4128 0 1 9828
box -48 -56 432 834
use sg13g2_nand3_1  _0893_
timestamp 1683988354
transform -1 0 4320 0 1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _0894_
timestamp 1677247768
transform 1 0 3840 0 -1 9828
box -48 -56 1008 834
use sg13g2_nor3_1  _0895_
timestamp 1676639442
transform -1 0 7392 0 1 9828
box -48 -56 528 834
use sg13g2_nor2b_1  _0896_
timestamp 1685181386
transform -1 0 6432 0 1 9828
box -54 -56 528 834
use sg13g2_a21oi_1  _0897_
timestamp 1683973020
transform 1 0 5952 0 -1 9828
box -48 -56 528 834
use sg13g2_nor2b_1  _0898_
timestamp 1685181386
transform 1 0 5088 0 -1 11340
box -54 -56 528 834
use sg13g2_a21oi_1  _0899_
timestamp 1683973020
transform 1 0 5568 0 -1 11340
box -48 -56 528 834
use sg13g2_a221oi_1  _0900_
timestamp 1685197497
transform -1 0 5760 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _0901_
timestamp 1685175443
transform 1 0 4800 0 -1 9828
box -48 -56 538 834
use sg13g2_nand2b_1  _0902_
timestamp 1676567195
transform -1 0 6528 0 -1 11340
box -48 -56 528 834
use sg13g2_nor3_1  _0903_
timestamp 1676639442
transform -1 0 5088 0 -1 8316
box -48 -56 528 834
use sg13g2_a21oi_1  _0904_
timestamp 1683973020
transform 1 0 4512 0 1 9828
box -48 -56 528 834
use sg13g2_nand3_1  _0905_
timestamp 1683988354
transform -1 0 4320 0 -1 8316
box -48 -56 528 834
use sg13g2_nor3_1  _0906_
timestamp 1676639442
transform 1 0 1152 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _0907_
timestamp 1685175443
transform -1 0 3360 0 -1 8316
box -48 -56 538 834
use sg13g2_nor2b_1  _0908_
timestamp 1685181386
transform 1 0 3072 0 1 9828
box -54 -56 528 834
use sg13g2_nor3_1  _0909_
timestamp 1676639442
transform 1 0 1152 0 1 11340
box -48 -56 528 834
use sg13g2_a21oi_1  _0910_
timestamp 1683973020
transform -1 0 3840 0 -1 8316
box -48 -56 528 834
use sg13g2_a22oi_1  _0911_
timestamp 1685173987
transform 1 0 3552 0 1 9828
box -48 -56 624 834
use sg13g2_dlhq_1  _0912_
timestamp 1678805552
transform 1 0 13920 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _0913_
timestamp 1678805552
transform -1 0 16896 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _0914_
timestamp 1678805552
transform 1 0 1248 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _0915_
timestamp 1678805552
transform 1 0 1536 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _0916_
timestamp 1678805552
transform 1 0 1344 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _0917_
timestamp 1678805552
transform 1 0 1248 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _0918_
timestamp 1678805552
transform 1 0 11424 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _0919_
timestamp 1678805552
transform 1 0 11232 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _0920_
timestamp 1678805552
transform 1 0 9024 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _0921_
timestamp 1678805552
transform 1 0 10944 0 1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _0922_
timestamp 1678805552
transform 1 0 6816 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _0923_
timestamp 1678805552
transform 1 0 8544 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _0924_
timestamp 1678805552
transform 1 0 7488 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0925_
timestamp 1678805552
transform 1 0 7200 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0926_
timestamp 1678805552
transform 1 0 8736 0 -1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _0927_
timestamp 1678805552
transform 1 0 10560 0 -1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _0928_
timestamp 1678805552
transform 1 0 6624 0 1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0929_
timestamp 1678805552
transform 1 0 8640 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0930_
timestamp 1678805552
transform 1 0 3648 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0931_
timestamp 1678805552
transform 1 0 5088 0 -1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0932_
timestamp 1678805552
transform 1 0 6720 0 -1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0933_
timestamp 1678805552
transform 1 0 7008 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0934_
timestamp 1678805552
transform 1 0 6624 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0935_
timestamp 1678805552
transform 1 0 6624 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0936_
timestamp 1678805552
transform 1 0 12960 0 -1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _0937_
timestamp 1678805552
transform 1 0 11424 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0938_
timestamp 1678805552
transform 1 0 1248 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0939_
timestamp 1678805552
transform 1 0 1152 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0940_
timestamp 1678805552
transform 1 0 1344 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _0941_
timestamp 1678805552
transform 1 0 1152 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _0942_
timestamp 1678805552
transform 1 0 10848 0 -1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0943_
timestamp 1678805552
transform 1 0 9120 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0944_
timestamp 1678805552
transform 1 0 13152 0 -1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0945_
timestamp 1678805552
transform 1 0 11616 0 1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _0946_
timestamp 1678805552
transform 1 0 2880 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0947_
timestamp 1678805552
transform 1 0 1440 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0948_
timestamp 1678805552
transform 1 0 2496 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _0949_
timestamp 1678805552
transform 1 0 1344 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0950_
timestamp 1678805552
transform 1 0 12960 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0951_
timestamp 1678805552
transform 1 0 10752 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0952_
timestamp 1678805552
transform 1 0 14976 0 -1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _0953_
timestamp 1678805552
transform 1 0 13248 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0954_
timestamp 1678805552
transform 1 0 2304 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0955_
timestamp 1678805552
transform 1 0 1152 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0956_
timestamp 1678805552
transform 1 0 1632 0 -1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _0957_
timestamp 1678805552
transform 1 0 1152 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0958_
timestamp 1678805552
transform 1 0 10272 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0959_
timestamp 1678805552
transform 1 0 8640 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0960_
timestamp 1678805552
transform 1 0 15264 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _0961_
timestamp 1678805552
transform 1 0 13344 0 1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _0962_
timestamp 1678805552
transform 1 0 2880 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0963_
timestamp 1678805552
transform 1 0 1440 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0964_
timestamp 1678805552
transform 1 0 2880 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _0965_
timestamp 1678805552
transform 1 0 1152 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _0966_
timestamp 1678805552
transform 1 0 11904 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0967_
timestamp 1678805552
transform 1 0 10272 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0968_
timestamp 1678805552
transform 1 0 15456 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _0969_
timestamp 1678805552
transform 1 0 15456 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _0970_
timestamp 1678805552
transform 1 0 14592 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _0971_
timestamp 1678805552
transform 1 0 1344 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _0972_
timestamp 1678805552
transform 1 0 1344 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _0973_
timestamp 1678805552
transform 1 0 1152 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0974_
timestamp 1678805552
transform 1 0 1920 0 1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _0975_
timestamp 1678805552
transform 1 0 3072 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _0976_
timestamp 1678805552
transform 1 0 1344 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _0977_
timestamp 1678805552
transform 1 0 15264 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _0978_
timestamp 1678805552
transform 1 0 14592 0 1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _0979_
timestamp 1678805552
transform 1 0 14592 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _0980_
timestamp 1678805552
transform -1 0 20064 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _0981_
timestamp 1678805552
transform -1 0 19776 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _0982_
timestamp 1678805552
transform 1 0 17952 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0983_
timestamp 1678805552
transform -1 0 7104 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0984_
timestamp 1678805552
transform 1 0 4128 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _0985_
timestamp 1678805552
transform 1 0 4320 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0986_
timestamp 1678805552
transform -1 0 4800 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _0987_
timestamp 1678805552
transform 1 0 1152 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _0988_
timestamp 1678805552
transform 1 0 1248 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _0989_
timestamp 1678805552
transform 1 0 16896 0 1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _0990_
timestamp 1678805552
transform 1 0 18528 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _0991_
timestamp 1678805552
transform 1 0 16896 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _0992_
timestamp 1678805552
transform 1 0 14880 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0993_
timestamp 1678805552
transform 1 0 17088 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0994_
timestamp 1678805552
transform 1 0 5280 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _0995_
timestamp 1678805552
transform 1 0 7104 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _0996_
timestamp 1678805552
transform 1 0 8352 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0997_
timestamp 1678805552
transform 1 0 10272 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0998_
timestamp 1678805552
transform -1 0 18528 0 1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0999_
timestamp 1678805552
transform 1 0 17664 0 -1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _1000_
timestamp 1678805552
transform 1 0 16896 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _1001_
timestamp 1678805552
transform 1 0 14976 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1002_
timestamp 1678805552
transform 1 0 5856 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1003_
timestamp 1678805552
transform 1 0 4224 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1004_
timestamp 1678805552
transform 1 0 8160 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1005_
timestamp 1678805552
transform 1 0 9984 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1006_
timestamp 1678805552
transform 1 0 15552 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _1007_
timestamp 1678805552
transform -1 0 20160 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _1008_
timestamp 1678805552
transform 1 0 15264 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _1009_
timestamp 1678805552
transform 1 0 13344 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1010_
timestamp 1678805552
transform 1 0 3936 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1011_
timestamp 1678805552
transform 1 0 3840 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1012_
timestamp 1678805552
transform 1 0 4512 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1013_
timestamp 1678805552
transform 1 0 3264 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1014_
timestamp 1678805552
transform 1 0 13824 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1015_
timestamp 1678805552
transform 1 0 11904 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1016_
timestamp 1678805552
transform 1 0 13440 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1017_
timestamp 1678805552
transform 1 0 11808 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1018_
timestamp 1678805552
transform 1 0 5376 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1019_
timestamp 1678805552
transform 1 0 4512 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1020_
timestamp 1678805552
transform -1 0 13152 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1021_
timestamp 1678805552
transform 1 0 8832 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1022_
timestamp 1678805552
transform 1 0 18048 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1023_
timestamp 1678805552
transform 1 0 15648 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1024_
timestamp 1678805552
transform -1 0 19296 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1025_
timestamp 1678805552
transform 1 0 13824 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1026_
timestamp 1678805552
transform 1 0 5568 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1027_
timestamp 1678805552
transform 1 0 4512 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1028_
timestamp 1678805552
transform 1 0 9696 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1029_
timestamp 1678805552
transform 1 0 7776 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1030_
timestamp 1678805552
transform 1 0 18048 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1031_
timestamp 1678805552
transform 1 0 16032 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1032_
timestamp 1678805552
transform 1 0 17664 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1033_
timestamp 1678805552
transform 1 0 15840 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1034_
timestamp 1678805552
transform 1 0 6144 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1035_
timestamp 1678805552
transform 1 0 4704 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1036_
timestamp 1678805552
transform 1 0 7776 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1037_
timestamp 1678805552
transform 1 0 6144 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1038_
timestamp 1678805552
transform 1 0 16032 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1039_
timestamp 1678805552
transform 1 0 14016 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1040_
timestamp 1678805552
transform 1 0 13344 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1041_
timestamp 1678805552
transform 1 0 11712 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1042_
timestamp 1678805552
transform 1 0 5760 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1043_
timestamp 1678805552
transform 1 0 4896 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1044_
timestamp 1678805552
transform 1 0 9024 0 -1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1045_
timestamp 1678805552
transform 1 0 5760 0 -1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1046_
timestamp 1678805552
transform 1 0 17184 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1047_
timestamp 1678805552
transform 1 0 15552 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1048_
timestamp 1678805552
transform 1 0 13920 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1049_
timestamp 1678805552
transform 1 0 12288 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1050_
timestamp 1678805552
transform 1 0 7392 0 -1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1051_
timestamp 1678805552
transform 1 0 4128 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1052_
timestamp 1678805552
transform 1 0 10656 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1053_
timestamp 1678805552
transform 1 0 9024 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1054_
timestamp 1678805552
transform 1 0 17664 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1055_
timestamp 1678805552
transform 1 0 15648 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1056_
timestamp 1678805552
transform 1 0 13920 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1057_
timestamp 1678805552
transform 1 0 12288 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1058_
timestamp 1678805552
transform 1 0 9024 0 -1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1059_
timestamp 1678805552
transform 1 0 8928 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1060_
timestamp 1678805552
transform 1 0 7488 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1061_
timestamp 1678805552
transform 1 0 5952 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1062_
timestamp 1678805552
transform 1 0 17952 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1063_
timestamp 1678805552
transform 1 0 15456 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1064_
timestamp 1678805552
transform 1 0 13728 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1065_
timestamp 1678805552
transform 1 0 12384 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1066_
timestamp 1678805552
transform 1 0 7296 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1067_
timestamp 1678805552
transform 1 0 5568 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1068_
timestamp 1678805552
transform 1 0 10560 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1069_
timestamp 1678805552
transform 1 0 8736 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1070_
timestamp 1678805552
transform 1 0 18048 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1071_
timestamp 1678805552
transform 1 0 15936 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1072_
timestamp 1678805552
transform 1 0 16128 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1073_
timestamp 1678805552
transform 1 0 14496 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1074_
timestamp 1678805552
transform 1 0 10848 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1075_
timestamp 1678805552
transform 1 0 9120 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1076_
timestamp 1678805552
transform 1 0 9600 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1077_
timestamp 1678805552
transform 1 0 7776 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1078_
timestamp 1678805552
transform 1 0 17568 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1079_
timestamp 1678805552
transform 1 0 15840 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1080_
timestamp 1678805552
transform 1 0 11424 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1081_
timestamp 1678805552
transform 1 0 13248 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1082_
timestamp 1678805552
transform 1 0 1344 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1083_
timestamp 1678805552
transform 1 0 2976 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1084_
timestamp 1678805552
transform 1 0 3456 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1085_
timestamp 1678805552
transform 1 0 5280 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1086_
timestamp 1678805552
transform 1 0 9888 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1087_
timestamp 1678805552
transform 1 0 11808 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1088_
timestamp 1678805552
transform 1 0 15648 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1089_
timestamp 1678805552
transform -1 0 16800 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1090_
timestamp 1678805552
transform 1 0 14784 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1091_
timestamp 1678805552
transform 1 0 8160 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1092_
timestamp 1678805552
transform 1 0 8928 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1093_
timestamp 1678805552
transform 1 0 7200 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1094_
timestamp 1678805552
transform 1 0 5472 0 1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1095_
timestamp 1678805552
transform 1 0 5184 0 1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1096_
timestamp 1678805552
transform 1 0 4800 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1097_
timestamp 1678805552
transform 1 0 11328 0 1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1098_
timestamp 1678805552
transform 1 0 11904 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1099_
timestamp 1678805552
transform 1 0 11232 0 1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1100_
timestamp 1678805552
transform 1 0 18336 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1101_
timestamp 1678805552
transform 1 0 16608 0 1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1102_
timestamp 1678805552
transform 1 0 8640 0 1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1103_
timestamp 1678805552
transform 1 0 6816 0 1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1104_
timestamp 1678805552
transform 1 0 9504 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1105_
timestamp 1678805552
transform 1 0 8352 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1106_
timestamp 1678805552
transform 1 0 17088 0 1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1107_
timestamp 1678805552
transform 1 0 18528 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1108_
timestamp 1678805552
transform 1 0 13152 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1109_
timestamp 1678805552
transform 1 0 11136 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1110_
timestamp 1678805552
transform 1 0 9792 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1111_
timestamp 1678805552
transform 1 0 8160 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1112_
timestamp 1678805552
transform 1 0 8256 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1113_
timestamp 1678805552
transform 1 0 6240 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1114_
timestamp 1678805552
transform -1 0 14400 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1115_
timestamp 1678805552
transform 1 0 11616 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1116_
timestamp 1678805552
transform 1 0 13920 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1117_
timestamp 1678805552
transform 1 0 11904 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1118_
timestamp 1678805552
transform 1 0 3264 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1119_
timestamp 1678805552
transform 1 0 1344 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1120_
timestamp 1678805552
transform 1 0 2880 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1121_
timestamp 1678805552
transform 1 0 1152 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1122_
timestamp 1678805552
transform 1 0 11136 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1123_
timestamp 1678805552
transform 1 0 12768 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1124_
timestamp 1678805552
transform 1 0 18336 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1125_
timestamp 1678805552
transform 1 0 18240 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1126_
timestamp 1678805552
transform 1 0 16224 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1127_
timestamp 1678805552
transform 1 0 5472 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1128_
timestamp 1678805552
transform 1 0 5760 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1129_
timestamp 1678805552
transform 1 0 4416 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1130_
timestamp 1678805552
transform 1 0 5280 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1131_
timestamp 1678805552
transform 1 0 5568 0 1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1132_
timestamp 1678805552
transform 1 0 4512 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1133_
timestamp 1678805552
transform 1 0 14880 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1134_
timestamp 1678805552
transform 1 0 14688 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1135_
timestamp 1678805552
transform 1 0 13632 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1136_
timestamp 1678805552
transform 1 0 18528 0 1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1137_
timestamp 1678805552
transform 1 0 16704 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1138_
timestamp 1678805552
transform 1 0 7872 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1139_
timestamp 1678805552
transform 1 0 6816 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1140_
timestamp 1678805552
transform 1 0 10464 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1141_
timestamp 1678805552
transform 1 0 8544 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1142_
timestamp 1678805552
transform 1 0 18624 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1143_
timestamp 1678805552
transform 1 0 17472 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1144_
timestamp 1678805552
transform 1 0 12864 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1145_
timestamp 1678805552
transform 1 0 11232 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1146_
timestamp 1678805552
transform 1 0 10176 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1147_
timestamp 1678805552
transform 1 0 7968 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1148_
timestamp 1678805552
transform -1 0 8256 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1149_
timestamp 1678805552
transform 1 0 4608 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1150_
timestamp 1678805552
transform -1 0 14880 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1151_
timestamp 1678805552
transform 1 0 11136 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1152_
timestamp 1678805552
transform 1 0 13632 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1153_
timestamp 1678805552
transform 1 0 11904 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1154_
timestamp 1678805552
transform 1 0 3360 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1155_
timestamp 1678805552
transform 1 0 1248 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1156_
timestamp 1678805552
transform -1 0 3936 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1157_
timestamp 1678805552
transform 1 0 1152 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1158_
timestamp 1678805552
transform 1 0 10848 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1159_
timestamp 1678805552
transform 1 0 12480 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1160_
timestamp 1678805552
transform 1 0 13344 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1161_
timestamp 1678805552
transform 1 0 13440 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1162_
timestamp 1678805552
transform 1 0 3264 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1163_
timestamp 1678805552
transform 1 0 1152 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1164_
timestamp 1678805552
transform 1 0 1920 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1165_
timestamp 1678805552
transform 1 0 1920 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1166_
timestamp 1678805552
transform 1 0 13344 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1167_
timestamp 1678805552
transform 1 0 13248 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1168_
timestamp 1678805552
transform 1 0 8928 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1169_
timestamp 1678805552
transform 1 0 7296 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1170_
timestamp 1678805552
transform 1 0 7296 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1171_
timestamp 1678805552
transform 1 0 5088 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1172_
timestamp 1678805552
transform 1 0 6720 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1173_
timestamp 1678805552
transform 1 0 6720 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1174_
timestamp 1678805552
transform 1 0 6720 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1175_
timestamp 1678805552
transform 1 0 7296 0 1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1176_
timestamp 1678805552
transform 1 0 7488 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1177_
timestamp 1678805552
transform 1 0 7104 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1178_
timestamp 1678805552
transform -1 0 5472 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1179_
timestamp 1678805552
transform 1 0 2208 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1180_
timestamp 1678805552
transform 1 0 7296 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1181_
timestamp 1678805552
transform 1 0 7296 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1182_
timestamp 1678805552
transform -1 0 9792 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1183_
timestamp 1678805552
transform 1 0 6528 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1184_
timestamp 1678805552
transform 1 0 10944 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1185_
timestamp 1678805552
transform 1 0 10656 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1186_
timestamp 1678805552
transform 1 0 1152 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1187_
timestamp 1678805552
transform 1 0 1152 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1188_
timestamp 1678805552
transform 1 0 3552 0 1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1189_
timestamp 1678805552
transform 1 0 1344 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1190_
timestamp 1678805552
transform 1 0 12192 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1191_
timestamp 1678805552
transform 1 0 10560 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1192_
timestamp 1678805552
transform 1 0 11904 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1193_
timestamp 1678805552
transform 1 0 10656 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1194_
timestamp 1678805552
transform 1 0 2400 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1195_
timestamp 1678805552
transform 1 0 1152 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1196_
timestamp 1678805552
transform -1 0 6720 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1197_
timestamp 1678805552
transform 1 0 1728 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1198_
timestamp 1678805552
transform 1 0 14592 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1199_
timestamp 1678805552
transform 1 0 12576 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1200_
timestamp 1678805552
transform -1 0 17856 0 1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1201_
timestamp 1678805552
transform 1 0 12576 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1202_
timestamp 1678805552
transform 1 0 1152 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1203_
timestamp 1678805552
transform 1 0 1152 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1204_
timestamp 1678805552
transform 1 0 2400 0 1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1205_
timestamp 1678805552
transform 1 0 1152 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1206_
timestamp 1678805552
transform 1 0 13056 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1207_
timestamp 1678805552
transform 1 0 11424 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1208_
timestamp 1678805552
transform 1 0 14592 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1209_
timestamp 1678805552
transform 1 0 12672 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1210_
timestamp 1678805552
transform 1 0 3264 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1211_
timestamp 1678805552
transform 1 0 1152 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1212_
timestamp 1678805552
transform 1 0 1824 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1213_
timestamp 1678805552
transform 1 0 1152 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1214_
timestamp 1678805552
transform 1 0 14880 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1215_
timestamp 1678805552
transform 1 0 12768 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1216_
timestamp 1678805552
transform 1 0 1152 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1217_
timestamp 1678805552
transform 1 0 1536 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1218_
timestamp 1678805552
transform 1 0 2784 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1219_
timestamp 1678805552
transform 1 0 1824 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1220_
timestamp 1678805552
transform 1 0 1632 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1221_
timestamp 1678805552
transform 1 0 1632 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1222_
timestamp 1678805552
transform 1 0 1632 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1223_
timestamp 1678805552
transform 1 0 1152 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1224_
timestamp 1678805552
transform 1 0 18528 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1225_
timestamp 1678805552
transform 1 0 16608 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1226_
timestamp 1678805552
transform 1 0 18720 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1227_
timestamp 1678805552
transform 1 0 1152 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1228_
timestamp 1678805552
transform 1 0 1152 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1229_
timestamp 1678805552
transform 1 0 1152 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1230_
timestamp 1678805552
transform 1 0 1920 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1231_
timestamp 1678805552
transform -1 0 5184 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1232_
timestamp 1678805552
transform 1 0 1632 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1233_
timestamp 1678805552
transform 1 0 17568 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1234_
timestamp 1678805552
transform 1 0 15648 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1235_
timestamp 1678805552
transform 1 0 18624 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1236_
timestamp 1678805552
transform 1 0 10080 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1237_
timestamp 1678805552
transform 1 0 11520 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1238_
timestamp 1678805552
transform 1 0 9888 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1239_
timestamp 1678805552
transform 1 0 1152 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1240_
timestamp 1678805552
transform 1 0 1440 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1241_
timestamp 1678805552
transform 1 0 1632 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1242_
timestamp 1678805552
transform 1 0 3264 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1243_
timestamp 1678805552
transform 1 0 4032 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1244_
timestamp 1678805552
transform 1 0 2400 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1245_
timestamp 1678805552
transform 1 0 18336 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1246_
timestamp 1678805552
transform 1 0 18624 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1247_
timestamp 1678805552
transform 1 0 17280 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1248_
timestamp 1678805552
transform 1 0 17088 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1249_
timestamp 1678805552
transform 1 0 18720 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1250_
timestamp 1678805552
transform 1 0 8352 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1251_
timestamp 1678805552
transform 1 0 10080 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1252_
timestamp 1678805552
transform 1 0 5664 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1253_
timestamp 1678805552
transform 1 0 7680 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1254_
timestamp 1678805552
transform 1 0 12672 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1255_
timestamp 1678805552
transform 1 0 14400 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1256_
timestamp 1678805552
transform 1 0 13248 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1257_
timestamp 1678805552
transform 1 0 14880 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1258_
timestamp 1678805552
transform 1 0 5568 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1259_
timestamp 1678805552
transform 1 0 7200 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1260_
timestamp 1678805552
transform 1 0 5376 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1261_
timestamp 1678805552
transform 1 0 7200 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1262_
timestamp 1678805552
transform 1 0 15456 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1263_
timestamp 1678805552
transform 1 0 12768 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1264_
timestamp 1678805552
transform -1 0 18816 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1265_
timestamp 1678805552
transform -1 0 16224 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1266_
timestamp 1678805552
transform 1 0 5664 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1267_
timestamp 1678805552
transform 1 0 4032 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1268_
timestamp 1678805552
transform 1 0 5664 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1269_
timestamp 1678805552
transform 1 0 3456 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1270_
timestamp 1678805552
transform -1 0 19104 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1271_
timestamp 1678805552
transform -1 0 16704 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1272_
timestamp 1678805552
transform 1 0 13248 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1273_
timestamp 1678805552
transform 1 0 17472 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1274_
timestamp 1678805552
transform 1 0 10752 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1275_
timestamp 1678805552
transform 1 0 8832 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1276_
timestamp 1678805552
transform 1 0 4992 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1277_
timestamp 1678805552
transform 1 0 6720 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1278_
timestamp 1678805552
transform 1 0 13536 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1279_
timestamp 1678805552
transform 1 0 11904 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1280_
timestamp 1678805552
transform 1 0 15936 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1281_
timestamp 1678805552
transform 1 0 18336 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1282_
timestamp 1678805552
transform 1 0 9984 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1283_
timestamp 1678805552
transform 1 0 8640 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1284_
timestamp 1678805552
transform 1 0 5952 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1285_
timestamp 1678805552
transform 1 0 7008 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1286_
timestamp 1678805552
transform -1 0 19680 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1287_
timestamp 1678805552
transform 1 0 17184 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1288_
timestamp 1678805552
transform -1 0 17472 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1289_
timestamp 1678805552
transform 1 0 17568 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1290_
timestamp 1678805552
transform 1 0 10944 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1291_
timestamp 1678805552
transform 1 0 9024 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1292_
timestamp 1678805552
transform 1 0 5376 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1293_
timestamp 1678805552
transform 1 0 6048 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1294_
timestamp 1678805552
transform 1 0 13920 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1295_
timestamp 1678805552
transform 1 0 12672 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1296_
timestamp 1678805552
transform 1 0 15552 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1297_
timestamp 1678805552
transform 1 0 17376 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1298_
timestamp 1678805552
transform 1 0 10176 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1299_
timestamp 1678805552
transform 1 0 8352 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1300_
timestamp 1678805552
transform 1 0 5952 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1301_
timestamp 1678805552
transform 1 0 7872 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1302_
timestamp 1678805552
transform 1 0 17760 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1303_
timestamp 1678805552
transform -1 0 18720 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1304_
timestamp 1678805552
transform 1 0 15744 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1305_
timestamp 1678805552
transform 1 0 15744 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1306_
timestamp 1678805552
transform -1 0 11232 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1307_
timestamp 1678805552
transform -1 0 11136 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1308_
timestamp 1678805552
transform 1 0 7968 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1309_
timestamp 1678805552
transform 1 0 8064 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1310_
timestamp 1678805552
transform 1 0 17376 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1311_
timestamp 1678805552
transform 1 0 17568 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1312_
timestamp 1678805552
transform 1 0 15552 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1313_
timestamp 1678805552
transform 1 0 15456 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1314_
timestamp 1678805552
transform 1 0 11616 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1315_
timestamp 1678805552
transform 1 0 11712 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1316_
timestamp 1678805552
transform 1 0 8736 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1317_
timestamp 1678805552
transform 1 0 8640 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1318_
timestamp 1678805552
transform 1 0 17280 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1319_
timestamp 1678805552
transform 1 0 17568 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1320_
timestamp 1678805552
transform 1 0 17760 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1321_
timestamp 1678805552
transform 1 0 17376 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1322_
timestamp 1678805552
transform 1 0 9600 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1323_
timestamp 1678805552
transform 1 0 9504 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1324_
timestamp 1678805552
transform 1 0 6720 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1325_
timestamp 1678805552
transform 1 0 6720 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1326_
timestamp 1678805552
transform 1 0 17568 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1327_
timestamp 1678805552
transform 1 0 17568 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1328_
timestamp 1678805552
transform 1 0 17280 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1329_
timestamp 1678805552
transform 1 0 18624 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1330_
timestamp 1678805552
transform 1 0 11328 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1331_
timestamp 1678805552
transform 1 0 11328 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1332_
timestamp 1678805552
transform -1 0 11040 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1333_
timestamp 1678805552
transform -1 0 10944 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1334_
timestamp 1678805552
transform 1 0 17568 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1335_
timestamp 1678805552
transform 1 0 17664 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1336_
timestamp 1678805552
transform 1 0 13152 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1337_
timestamp 1678805552
transform 1 0 15072 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1338_
timestamp 1678805552
transform 1 0 1152 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1339_
timestamp 1678805552
transform 1 0 1536 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1340_
timestamp 1678805552
transform -1 0 3552 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1341_
timestamp 1678805552
transform 1 0 1920 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1342_
timestamp 1678805552
transform 1 0 11232 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1343_
timestamp 1678805552
transform 1 0 13344 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1344_
timestamp 1678805552
transform 1 0 15840 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1345_
timestamp 1678805552
transform 1 0 13920 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1346_
timestamp 1678805552
transform 1 0 13728 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1347_
timestamp 1678805552
transform 1 0 5376 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1348_
timestamp 1678805552
transform 1 0 5376 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1349_
timestamp 1678805552
transform 1 0 4416 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1350_
timestamp 1678805552
transform -1 0 11904 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1351_
timestamp 1678805552
transform 1 0 10464 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1352_
timestamp 1678805552
transform 1 0 8448 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1353_
timestamp 1678805552
transform 1 0 15456 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1354_
timestamp 1678805552
transform 1 0 15552 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1355_
timestamp 1678805552
transform 1 0 14208 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1356_
timestamp 1678805552
transform 1 0 10848 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1357_
timestamp 1678805552
transform 1 0 12672 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1358_
timestamp 1678805552
transform 1 0 7104 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1359_
timestamp 1678805552
transform 1 0 8832 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1360_
timestamp 1678805552
transform 1 0 6432 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1361_
timestamp 1678805552
transform 1 0 8352 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1362_
timestamp 1678805552
transform 1 0 9600 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1363_
timestamp 1678805552
transform 1 0 11136 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1364_
timestamp 1678805552
transform 1 0 10752 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1365_
timestamp 1678805552
transform 1 0 8256 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1366_
timestamp 1678805552
transform 1 0 6624 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1367_
timestamp 1678805552
transform 1 0 5472 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1368_
timestamp 1678805552
transform 1 0 7584 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1369_
timestamp 1678805552
transform 1 0 5760 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1370_
timestamp 1678805552
transform 1 0 13632 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1371_
timestamp 1678805552
transform 1 0 11520 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1372_
timestamp 1678805552
transform 1 0 12480 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1373_
timestamp 1678805552
transform 1 0 10848 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1374_
timestamp 1678805552
transform 1 0 4704 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1375_
timestamp 1678805552
transform 1 0 2976 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1376_
timestamp 1678805552
transform 1 0 6048 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1377_
timestamp 1678805552
transform 1 0 4032 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1378_
timestamp 1678805552
transform 1 0 13248 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1379_
timestamp 1678805552
transform 1 0 11616 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1380_
timestamp 1678805552
transform -1 0 13920 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1381_
timestamp 1678805552
transform 1 0 12000 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1382_
timestamp 1678805552
transform 1 0 13920 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1383_
timestamp 1678805552
transform 1 0 3648 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1384_
timestamp 1678805552
transform 1 0 1920 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1385_
timestamp 1678805552
transform 1 0 3552 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1386_
timestamp 1678805552
transform 1 0 5472 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1387_
timestamp 1678805552
transform 1 0 4416 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1388_
timestamp 1678805552
transform 1 0 5184 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1389_
timestamp 1678805552
transform -1 0 17088 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1390_
timestamp 1678805552
transform 1 0 13824 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1391_
timestamp 1678805552
transform 1 0 15264 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1392_
timestamp 1678805552
transform 1 0 14976 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1393_
timestamp 1678805552
transform 1 0 13344 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1394_
timestamp 1678805552
transform 1 0 6816 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1395_
timestamp 1678805552
transform 1 0 4800 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1396_
timestamp 1678805552
transform 1 0 7488 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1397_
timestamp 1678805552
transform 1 0 4896 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1398_
timestamp 1678805552
transform 1 0 9888 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1399_
timestamp 1678805552
transform 1 0 8832 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1400_
timestamp 1678805552
transform 1 0 11328 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1401_
timestamp 1678805552
transform 1 0 9504 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1402_
timestamp 1678805552
transform 1 0 3936 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1403_
timestamp 1678805552
transform 1 0 1632 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1404_
timestamp 1678805552
transform 1 0 7008 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1405_
timestamp 1678805552
transform 1 0 5280 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1406_
timestamp 1678805552
transform -1 0 16896 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1407_
timestamp 1678805552
transform 1 0 11520 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1408_
timestamp 1678805552
transform 1 0 11328 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1409_
timestamp 1678805552
transform 1 0 13152 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1410_
timestamp 1678805552
transform 1 0 1152 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1411_
timestamp 1678805552
transform 1 0 2784 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1412_
timestamp 1678805552
transform 1 0 2784 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1413_
timestamp 1678805552
transform -1 0 4416 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1414_
timestamp 1678805552
transform 1 0 9888 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1415_
timestamp 1678805552
transform 1 0 12960 0 -1 12852
box -50 -56 1692 834
use sg13g2_buf_1  _1416_
timestamp 1676381911
transform -1 0 2208 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1417_
timestamp 1676381911
transform 1 0 19680 0 1 58212
box -48 -56 432 834
use sg13g2_buf_1  _1418_
timestamp 1676381911
transform 1 0 19680 0 -1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1419_
timestamp 1676381911
transform 1 0 19680 0 1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1420_
timestamp 1676381911
transform 1 0 19968 0 -1 61236
box -48 -56 432 834
use sg13g2_buf_1  _1421_
timestamp 1676381911
transform 1 0 19776 0 -1 58212
box -48 -56 432 834
use sg13g2_buf_1  _1422_
timestamp 1676381911
transform 1 0 19296 0 1 58212
box -48 -56 432 834
use sg13g2_buf_1  _1423_
timestamp 1676381911
transform 1 0 19296 0 1 61236
box -48 -56 432 834
use sg13g2_buf_1  _1424_
timestamp 1676381911
transform 1 0 18912 0 1 61236
box -48 -56 432 834
use sg13g2_buf_1  _1425_
timestamp 1676381911
transform 1 0 19680 0 1 61236
box -48 -56 432 834
use sg13g2_buf_1  _1426_
timestamp 1676381911
transform 1 0 18528 0 1 61236
box -48 -56 432 834
use sg13g2_buf_1  _1427_
timestamp 1676381911
transform 1 0 19584 0 -1 62748
box -48 -56 432 834
use sg13g2_buf_1  _1428_
timestamp 1676381911
transform 1 0 19968 0 -1 62748
box -48 -56 432 834
use sg13g2_buf_1  _1429_
timestamp 1676381911
transform 1 0 19392 0 1 62748
box -48 -56 432 834
use sg13g2_buf_1  _1430_
timestamp 1676381911
transform 1 0 19296 0 -1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1431_
timestamp 1676381911
transform 1 0 19296 0 -1 64260
box -48 -56 432 834
use sg13g2_buf_1  _1432_
timestamp 1676381911
transform 1 0 19680 0 -1 64260
box -48 -56 432 834
use sg13g2_buf_1  _1433_
timestamp 1676381911
transform 1 0 19296 0 1 64260
box -48 -56 432 834
use sg13g2_buf_1  _1434_
timestamp 1676381911
transform 1 0 18912 0 -1 65772
box -48 -56 432 834
use sg13g2_buf_1  _1435_
timestamp 1676381911
transform 1 0 19680 0 1 64260
box -48 -56 432 834
use sg13g2_buf_1  _1436_
timestamp 1676381911
transform 1 0 19680 0 -1 65772
box -48 -56 432 834
use sg13g2_buf_1  _1437_
timestamp 1676381911
transform 1 0 19296 0 -1 73332
box -48 -56 432 834
use sg13g2_buf_1  _1438_
timestamp 1676381911
transform 1 0 19680 0 -1 73332
box -48 -56 432 834
use sg13g2_buf_1  _1439_
timestamp 1676381911
transform 1 0 8448 0 -1 71820
box -48 -56 432 834
use sg13g2_buf_1  _1440_
timestamp 1676381911
transform 1 0 19776 0 -1 74844
box -48 -56 432 834
use sg13g2_buf_1  _1441_
timestamp 1676381911
transform 1 0 19392 0 -1 74844
box -48 -56 432 834
use sg13g2_buf_1  _1442_
timestamp 1676381911
transform 1 0 19296 0 1 73332
box -48 -56 432 834
use sg13g2_buf_1  _1443_
timestamp 1676381911
transform 1 0 18528 0 -1 73332
box -48 -56 432 834
use sg13g2_buf_1  _1444_
timestamp 1676381911
transform 1 0 18912 0 1 73332
box -48 -56 432 834
use sg13g2_buf_1  _1445_
timestamp 1676381911
transform 1 0 19680 0 -1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1446_
timestamp 1676381911
transform 1 0 19488 0 -1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1447_
timestamp 1676381911
transform 1 0 19872 0 -1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1448_
timestamp 1676381911
transform 1 0 19488 0 1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1449_
timestamp 1676381911
transform 1 0 19296 0 1 65772
box -48 -56 432 834
use sg13g2_buf_1  _1450_
timestamp 1676381911
transform 1 0 19680 0 1 65772
box -48 -56 432 834
use sg13g2_buf_1  _1451_
timestamp 1676381911
transform 1 0 19296 0 -1 65772
box -48 -56 432 834
use sg13g2_buf_1  _1452_
timestamp 1676381911
transform 1 0 19680 0 1 67284
box -48 -56 432 834
use sg13g2_buf_1  _1453_
timestamp 1676381911
transform 1 0 19872 0 -1 68796
box -48 -56 432 834
use sg13g2_buf_1  _1454_
timestamp 1676381911
transform 1 0 19488 0 -1 68796
box -48 -56 432 834
use sg13g2_buf_1  _1455_
timestamp 1676381911
transform 1 0 19872 0 -1 70308
box -48 -56 432 834
use sg13g2_buf_1  _1456_
timestamp 1676381911
transform 1 0 19680 0 1 68796
box -48 -56 432 834
use sg13g2_buf_1  _1457_
timestamp 1676381911
transform 1 0 19488 0 -1 70308
box -48 -56 432 834
use sg13g2_buf_1  _1458_
timestamp 1676381911
transform 1 0 19680 0 1 70308
box -48 -56 432 834
use sg13g2_buf_1  _1459_
timestamp 1676381911
transform 1 0 19296 0 1 70308
box -48 -56 432 834
use sg13g2_buf_1  _1460_
timestamp 1676381911
transform 1 0 19296 0 -1 71820
box -48 -56 432 834
use sg13g2_buf_1  _1461_
timestamp 1676381911
transform 1 0 17664 0 1 68796
box -48 -56 432 834
use sg13g2_buf_1  _1462_
timestamp 1676381911
transform 1 0 19872 0 -1 71820
box -48 -56 432 834
use sg13g2_buf_1  _1463_
timestamp 1676381911
transform 1 0 19680 0 1 71820
box -48 -56 432 834
use sg13g2_buf_1  _1464_
timestamp 1676381911
transform 1 0 19296 0 1 71820
box -48 -56 432 834
use sg13g2_buf_1  _1465_
timestamp 1676381911
transform 1 0 19872 0 1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1466_
timestamp 1676381911
transform 1 0 19296 0 -1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1467_
timestamp 1676381911
transform 1 0 18912 0 1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1468_
timestamp 1676381911
transform 1 0 19296 0 1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1469_
timestamp 1676381911
transform 1 0 18528 0 1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1470_
timestamp 1676381911
transform 1 0 19680 0 1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1471_
timestamp 1676381911
transform 1 0 15168 0 -1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1472_
timestamp 1676381911
transform 1 0 19296 0 -1 79380
box -48 -56 432 834
use sg13g2_buf_1  _1473_
timestamp 1676381911
transform 1 0 19680 0 -1 79380
box -48 -56 432 834
use sg13g2_buf_1  _1474_
timestamp 1676381911
transform 1 0 18912 0 1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1475_
timestamp 1676381911
transform 1 0 19296 0 1 79380
box -48 -56 432 834
use sg13g2_buf_1  _1476_
timestamp 1676381911
transform 1 0 18528 0 1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1477_
timestamp 1676381911
transform 1 0 18912 0 -1 79380
box -48 -56 432 834
use sg13g2_buf_1  _1478_
timestamp 1676381911
transform 1 0 19680 0 1 79380
box -48 -56 432 834
use sg13g2_buf_1  _1479_
timestamp 1676381911
transform 1 0 19296 0 -1 80892
box -48 -56 432 834
use sg13g2_buf_1  _1480_
timestamp 1676381911
transform 1 0 16416 0 1 79380
box -48 -56 432 834
use sg13g2_buf_1  _1481_
timestamp 1676381911
transform 1 0 18912 0 1 79380
box -48 -56 432 834
use sg13g2_buf_1  _1482_
timestamp 1676381911
transform 1 0 18624 0 -1 80892
box -48 -56 432 834
use sg13g2_buf_1  _1483_
timestamp 1676381911
transform 1 0 19680 0 -1 80892
box -48 -56 432 834
use sg13g2_buf_1  _1484_
timestamp 1676381911
transform 1 0 19296 0 1 80892
box -48 -56 432 834
use sg13g2_buf_1  _1485_
timestamp 1676381911
transform 1 0 18912 0 -1 73332
box -48 -56 432 834
use sg13g2_buf_1  _1486_
timestamp 1676381911
transform 1 0 18912 0 1 80892
box -48 -56 432 834
use sg13g2_buf_1  _1487_
timestamp 1676381911
transform 1 0 14016 0 -1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1488_
timestamp 1676381911
transform 1 0 15456 0 -1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1489_
timestamp 1676381911
transform 1 0 19296 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1490_
timestamp 1676381911
transform 1 0 18912 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1491_
timestamp 1676381911
transform 1 0 19584 0 -1 67284
box -48 -56 432 834
use sg13g2_buf_1  _1492_
timestamp 1676381911
transform 1 0 19968 0 -1 67284
box -48 -56 432 834
use sg13g2_buf_1  _1493_
timestamp 1676381911
transform 1 0 18912 0 1 71820
box -48 -56 432 834
use sg13g2_buf_1  _1494_
timestamp 1676381911
transform 1 0 19680 0 1 73332
box -48 -56 432 834
use sg13g2_buf_1  _1495_
timestamp 1676381911
transform 1 0 19296 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1496_
timestamp 1676381911
transform 1 0 18912 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1497_
timestamp 1676381911
transform 1 0 15456 0 1 79380
box -48 -56 432 834
use sg13g2_buf_1  _1498_
timestamp 1676381911
transform -1 0 16224 0 1 79380
box -48 -56 432 834
use sg13g2_buf_1  _1499_
timestamp 1676381911
transform -1 0 17376 0 -1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1500_
timestamp 1676381911
transform -1 0 16992 0 -1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1501_
timestamp 1676381911
transform 1 0 15648 0 1 67284
box -48 -56 432 834
use sg13g2_buf_1  _1502_
timestamp 1676381911
transform 1 0 16512 0 -1 62748
box -48 -56 432 834
use sg13g2_buf_1  _1503_
timestamp 1676381911
transform 1 0 16608 0 -1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1504_
timestamp 1676381911
transform 1 0 16416 0 -1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1505_
timestamp 1676381911
transform -1 0 17568 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1506_
timestamp 1676381911
transform -1 0 17952 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1507_
timestamp 1676381911
transform -1 0 18336 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1508_
timestamp 1676381911
transform -1 0 18720 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1509_
timestamp 1676381911
transform -1 0 18336 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1510_
timestamp 1676381911
transform -1 0 19104 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1511_
timestamp 1676381911
transform -1 0 18720 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1512_
timestamp 1676381911
transform -1 0 19488 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1513_
timestamp 1676381911
transform -1 0 19104 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1514_
timestamp 1676381911
transform -1 0 19872 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1515_
timestamp 1676381911
transform -1 0 19488 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1516_
timestamp 1676381911
transform -1 0 20256 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1517_
timestamp 1676381911
transform 1 0 1440 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1518_
timestamp 1676381911
transform -1 0 2208 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1519_
timestamp 1676381911
transform -1 0 2976 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1520_
timestamp 1676381911
transform -1 0 2592 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1521_
timestamp 1676381911
transform -1 0 3360 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1522_
timestamp 1676381911
transform -1 0 2976 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1523_
timestamp 1676381911
transform -1 0 3744 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1524_
timestamp 1676381911
transform -1 0 3360 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1525_
timestamp 1676381911
transform -1 0 4224 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1526_
timestamp 1676381911
transform -1 0 3744 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1527_
timestamp 1676381911
transform -1 0 4608 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1528_
timestamp 1676381911
transform -1 0 4128 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1529_
timestamp 1676381911
transform -1 0 4896 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1530_
timestamp 1676381911
transform -1 0 4512 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1531_
timestamp 1676381911
transform -1 0 4896 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1532_
timestamp 1676381911
transform -1 0 5280 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1533_
timestamp 1676381911
transform -1 0 5664 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1534_
timestamp 1676381911
transform -1 0 8832 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1535_
timestamp 1676381911
transform -1 0 8064 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1536_
timestamp 1676381911
transform -1 0 6240 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1537_
timestamp 1676381911
transform -1 0 6048 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1538_
timestamp 1676381911
transform -1 0 6816 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1539_
timestamp 1676381911
transform -1 0 6432 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1540_
timestamp 1676381911
transform -1 0 7200 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1541_
timestamp 1676381911
transform -1 0 6816 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1542_
timestamp 1676381911
transform -1 0 7200 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1543_
timestamp 1676381911
transform -1 0 7584 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1544_
timestamp 1676381911
transform -1 0 7968 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1545_
timestamp 1676381911
transform -1 0 16032 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1546_
timestamp 1676381911
transform 1 0 6912 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1547_
timestamp 1676381911
transform 1 0 6432 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1548_
timestamp 1676381911
transform -1 0 13632 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1549_
timestamp 1676381911
transform -1 0 15264 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1550_
timestamp 1676381911
transform 1 0 7296 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1551_
timestamp 1676381911
transform 1 0 8064 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1552_
timestamp 1676381911
transform -1 0 18432 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1553_
timestamp 1676381911
transform 1 0 15264 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1554_
timestamp 1676381911
transform 1 0 19200 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _1555_
timestamp 1676381911
transform 1 0 4224 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1556_
timestamp 1676381911
transform 1 0 3360 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1557_
timestamp 1676381911
transform 1 0 16128 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _1558_
timestamp 1676381911
transform 1 0 17568 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1559_
timestamp 1676381911
transform 1 0 17184 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1560_
timestamp 1676381911
transform 1 0 16512 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _1561_
timestamp 1676381911
transform 1 0 19968 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1562_
timestamp 1676381911
transform 1 0 19968 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1563_
timestamp 1676381911
transform 1 0 16896 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _1564_
timestamp 1676381911
transform 1 0 19968 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1565_
timestamp 1676381911
transform 1 0 19968 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1566_
timestamp 1676381911
transform 1 0 15168 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1567_
timestamp 1676381911
transform 1 0 19200 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1568_
timestamp 1676381911
transform 1 0 19776 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1569_
timestamp 1676381911
transform 1 0 19584 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1570_
timestamp 1676381911
transform 1 0 19584 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _1571_
timestamp 1676381911
transform 1 0 19968 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _1572_
timestamp 1676381911
transform 1 0 15168 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1573_
timestamp 1676381911
transform 1 0 19968 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1574_
timestamp 1676381911
transform 1 0 19584 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1575_
timestamp 1676381911
transform 1 0 19584 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1576_
timestamp 1676381911
transform 1 0 19200 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1577_
timestamp 1676381911
transform 1 0 19968 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1578_
timestamp 1676381911
transform 1 0 19776 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1579_
timestamp 1676381911
transform 1 0 19776 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1580_
timestamp 1676381911
transform 1 0 19488 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1581_
timestamp 1676381911
transform 1 0 19872 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1582_
timestamp 1676381911
transform 1 0 19296 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1583_
timestamp 1676381911
transform 1 0 17088 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1584_
timestamp 1676381911
transform 1 0 19968 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1585_
timestamp 1676381911
transform 1 0 19776 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1586_
timestamp 1676381911
transform 1 0 19968 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1587_
timestamp 1676381911
transform 1 0 16896 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _1588_
timestamp 1676381911
transform 1 0 17088 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1589_
timestamp 1676381911
transform 1 0 19296 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1590_
timestamp 1676381911
transform 1 0 19680 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1591_
timestamp 1676381911
transform 1 0 17184 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  _1592_
timestamp 1676381911
transform 1 0 19296 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1593_
timestamp 1676381911
transform 1 0 16992 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1594_
timestamp 1676381911
transform 1 0 16704 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1595_
timestamp 1676381911
transform 1 0 19968 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  _1596_
timestamp 1676381911
transform 1 0 15168 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1597_
timestamp 1676381911
transform 1 0 19104 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1598_
timestamp 1676381911
transform 1 0 19968 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1599_
timestamp 1676381911
transform 1 0 15168 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1600_
timestamp 1676381911
transform 1 0 16704 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1601_
timestamp 1676381911
transform 1 0 19392 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1602_
timestamp 1676381911
transform 1 0 19584 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1603_
timestamp 1676381911
transform 1 0 19392 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1604_
timestamp 1676381911
transform 1 0 19680 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1605_
timestamp 1676381911
transform 1 0 18528 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1606_
timestamp 1676381911
transform 1 0 12384 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1607_
timestamp 1676381911
transform 1 0 18912 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1608_
timestamp 1676381911
transform 1 0 19296 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1609_
timestamp 1676381911
transform 1 0 16608 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1610_
timestamp 1676381911
transform 1 0 19680 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1611_
timestamp 1676381911
transform 1 0 19296 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1612_
timestamp 1676381911
transform 1 0 19392 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1613_
timestamp 1676381911
transform 1 0 19776 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1614_
timestamp 1676381911
transform 1 0 19392 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1615_
timestamp 1676381911
transform 1 0 19872 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1616_
timestamp 1676381911
transform 1 0 19488 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1617_
timestamp 1676381911
transform 1 0 19968 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1618_
timestamp 1676381911
transform 1 0 18528 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1619_
timestamp 1676381911
transform 1 0 19968 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1620_
timestamp 1676381911
transform 1 0 19200 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1621_
timestamp 1676381911
transform 1 0 19200 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1622_
timestamp 1676381911
transform 1 0 19584 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1623_
timestamp 1676381911
transform 1 0 19200 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1624_
timestamp 1676381911
transform 1 0 19584 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1625_
timestamp 1676381911
transform 1 0 18912 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1626_
timestamp 1676381911
transform 1 0 17760 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1627_
timestamp 1676381911
transform 1 0 19296 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1628_
timestamp 1676381911
transform 1 0 19200 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1629_
timestamp 1676381911
transform 1 0 19584 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1630_
timestamp 1676381911
transform 1 0 19200 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1631_
timestamp 1676381911
transform 1 0 19584 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1632_
timestamp 1676381911
transform 1 0 17856 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1633_
timestamp 1676381911
transform 1 0 19968 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1634_
timestamp 1676381911
transform -1 0 9504 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1635_
timestamp 1676381911
transform 1 0 8064 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1636_
timestamp 1676381911
transform 1 0 6816 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1637_
timestamp 1676381911
transform -1 0 9696 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1638_
timestamp 1676381911
transform -1 0 15840 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1639_
timestamp 1676381911
transform 1 0 8928 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1640_
timestamp 1676381911
transform 1 0 8544 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1641_
timestamp 1676381911
transform -1 0 11616 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1642_
timestamp 1676381911
transform -1 0 11808 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1643_
timestamp 1676381911
transform 1 0 10080 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1644_
timestamp 1676381911
transform 1 0 9696 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1645_
timestamp 1676381911
transform -1 0 13440 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1646_
timestamp 1676381911
transform 1 0 10080 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1647_
timestamp 1676381911
transform 1 0 10272 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1648_
timestamp 1676381911
transform 1 0 11040 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1649_
timestamp 1676381911
transform 1 0 11328 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1650_
timestamp 1676381911
transform 1 0 11520 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1651_
timestamp 1676381911
transform 1 0 10848 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1652_
timestamp 1676381911
transform 1 0 10464 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1653_
timestamp 1676381911
transform 1 0 12000 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1654_
timestamp 1676381911
transform -1 0 14400 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1655_
timestamp 1676381911
transform -1 0 14784 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1656_
timestamp 1676381911
transform -1 0 15072 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1657_
timestamp 1676381911
transform -1 0 14688 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1658_
timestamp 1676381911
transform -1 0 15456 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1659_
timestamp 1676381911
transform 1 0 12960 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1660_
timestamp 1676381911
transform -1 0 15744 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1661_
timestamp 1676381911
transform -1 0 16128 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1662_
timestamp 1676381911
transform 1 0 13728 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1663_
timestamp 1676381911
transform 1 0 13344 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1664_
timestamp 1676381911
transform 1 0 11616 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1665_
timestamp 1676381911
transform -1 0 16224 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1666_
timestamp 1676381911
transform -1 0 16512 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1667_
timestamp 1676381911
transform 1 0 12672 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1668_
timestamp 1676381911
transform 1 0 14304 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1669_
timestamp 1676381911
transform -1 0 16896 0 -1 2268
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 8928 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 16224 0 -1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform 1 0 1632 0 1 26460
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 17184 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 15552 0 1 24948
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform 1 0 17280 0 -1 6804
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform 1 0 6432 0 -1 6804
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform 1 0 14976 0 1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform 1 0 18912 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform 1 0 8928 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform 1 0 16224 0 -1 43092
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform 1 0 1632 0 1 27972
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform 1 0 17184 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 15840 0 1 26460
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform 1 0 17280 0 -1 8316
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform 1 0 6144 0 -1 8316
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 14976 0 1 6804
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform 1 0 18912 0 -1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform 1 0 8928 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform 1 0 16224 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform 1 0 1632 0 -1 26460
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform 1 0 17184 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform 1 0 15552 0 -1 24948
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform 1 0 17280 0 1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform 1 0 6432 0 1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_26
timestamp 1679999689
transform 1 0 14976 0 -1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_27
timestamp 1679999689
transform 1 0 18912 0 1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_28
timestamp 1679999689
transform 1 0 8928 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_29
timestamp 1679999689
transform 1 0 16224 0 1 43092
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_30
timestamp 1679999689
transform 1 0 1632 0 -1 29484
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_31
timestamp 1679999689
transform 1 0 17184 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_32
timestamp 1679999689
transform 1 0 15552 0 1 26460
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_33
timestamp 1679999689
transform 1 0 17280 0 1 8316
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_34
timestamp 1679999689
transform 1 0 6432 0 -1 8316
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_35
timestamp 1679999689
transform 1 0 14976 0 -1 8316
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_36
timestamp 1679999689
transform 1 0 18912 0 1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_37
timestamp 1679999689
transform 1 0 8928 0 -1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_38
timestamp 1679999689
transform 1 0 16224 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_39
timestamp 1679999689
transform 1 0 1632 0 1 24948
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_40
timestamp 1679999689
transform 1 0 17184 0 -1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_41
timestamp 1679999689
transform 1 0 15552 0 1 23436
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_42
timestamp 1679999689
transform 1 0 17280 0 -1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_43
timestamp 1679999689
transform 1 0 6432 0 -1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_44
timestamp 1679999689
transform 1 0 14976 0 1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_45
timestamp 1679999689
transform 1 0 18912 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_46
timestamp 1679999689
transform 1 0 8928 0 1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_47
timestamp 1679999689
transform 1 0 16224 0 -1 44604
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_48
timestamp 1679999689
transform 1 0 1632 0 1 29484
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_49
timestamp 1679999689
transform 1 0 17184 0 -1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_50
timestamp 1679999689
transform 1 0 15552 0 -1 27972
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_51
timestamp 1679999689
transform 1 0 17280 0 -1 9828
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_52
timestamp 1679999689
transform 1 0 6432 0 1 8316
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_53
timestamp 1679999689
transform 1 0 14976 0 1 8316
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_54
timestamp 1679999689
transform 1 0 18912 0 -1 43092
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_55
timestamp 1679999689
transform 1 0 8928 0 1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_56
timestamp 1679999689
transform 1 0 16224 0 1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_57
timestamp 1679999689
transform 1 0 1632 0 -1 24948
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_58
timestamp 1679999689
transform 1 0 17184 0 1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_59
timestamp 1679999689
transform 1 0 15552 0 -1 23436
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_60
timestamp 1679999689
transform 1 0 17280 0 1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_61
timestamp 1679999689
transform 1 0 6432 0 1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_62
timestamp 1679999689
transform 1 0 14976 0 -1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_63
timestamp 1679999689
transform 1 0 18912 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_64
timestamp 1679999689
transform 1 0 8928 0 -1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_65
timestamp 1679999689
transform 1 0 16224 0 1 44604
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_66
timestamp 1679999689
transform 1 0 1632 0 -1 30996
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_67
timestamp 1679999689
transform 1 0 17184 0 -1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_68
timestamp 1679999689
transform 1 0 15552 0 -1 29484
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_69
timestamp 1679999689
transform 1 0 17280 0 1 9828
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_70
timestamp 1679999689
transform 1 0 6816 0 -1 11340
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_71
timestamp 1679999689
transform 1 0 14976 0 -1 9828
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_72
timestamp 1679999689
transform 1 0 18912 0 1 43092
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_73
timestamp 1679999689
transform 1 0 8928 0 -1 43092
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_74
timestamp 1679999689
transform 1 0 16224 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_75
timestamp 1679999689
transform 1 0 1344 0 1 23436
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_76
timestamp 1679999689
transform 1 0 17184 0 -1 43092
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_77
timestamp 1679999689
transform 1 0 15552 0 1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_78
timestamp 1679999689
transform 1 0 17280 0 -1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_79
timestamp 1679999689
transform 1 0 6432 0 -1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_80
timestamp 1679999689
transform -1 0 15264 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_81
timestamp 1679999689
transform 1 0 18912 0 -1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_82
timestamp 1679999689
transform -1 0 7104 0 -1 12852
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_83
timestamp 1679999689
transform 1 0 12768 0 -1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_84
timestamp 1679999689
transform -1 0 17568 0 -1 12852
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_85
timestamp 1679999689
transform 1 0 11904 0 -1 32508
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_86
timestamp 1679999689
transform 1 0 17568 0 1 20412
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_87
timestamp 1679999689
transform 1 0 13344 0 -1 15876
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_88
timestamp 1679999689
transform 1 0 2976 0 -1 18900
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_89
timestamp 1679999689
transform 1 0 11520 0 1 12852
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_90
timestamp 1679999689
transform 1 0 19680 0 1 32508
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_91
timestamp 1679999689
transform 1 0 9504 0 -1 43092
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_92
timestamp 1679999689
transform 1 0 10272 0 -1 76356
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_93
timestamp 1679999689
transform 1 0 8352 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_94
timestamp 1679999689
transform 1 0 8832 0 1 70308
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_95
timestamp 1679999689
transform 1 0 9984 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_96
timestamp 1679999689
transform 1 0 10656 0 1 77868
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_97
timestamp 1679999689
transform 1 0 9984 0 -1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_98
timestamp 1679999689
transform -1 0 10944 0 1 79380
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_99
timestamp 1679999689
transform 1 0 2976 0 1 58212
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_100
timestamp 1679999689
transform 1 0 2688 0 -1 59724
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_101
timestamp 1679999689
transform 1 0 16992 0 -1 59724
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_102
timestamp 1679999689
transform 1 0 17088 0 1 62748
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_103
timestamp 1679999689
transform 1 0 16128 0 -1 65772
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_104
timestamp 1679999689
transform 1 0 16992 0 1 65772
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_105
timestamp 1679999689
transform 1 0 17184 0 -1 76356
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_106
timestamp 1679999689
transform 1 0 6528 0 1 9828
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_107
timestamp 1679999689
transform 1 0 9120 0 1 9828
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_108
timestamp 1679999689
transform 1 0 8256 0 -1 76356
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_109
timestamp 1679999689
transform -1 0 4800 0 1 11340
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_110
timestamp 1679999689
transform 1 0 6528 0 1 11340
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_111
timestamp 1679999689
transform 1 0 9120 0 1 11340
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_112
timestamp 1679999689
transform 1 0 8256 0 -1 77868
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_113
timestamp 1679999689
transform -1 0 4800 0 1 12852
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_114
timestamp 1679999689
transform -1 0 6816 0 -1 9828
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_115
timestamp 1679999689
transform -1 0 9408 0 -1 9828
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_116
timestamp 1679999689
transform 1 0 8256 0 1 74844
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_117
timestamp 1679999689
transform -1 0 4800 0 -1 11340
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_118
timestamp 1679999689
transform 1 0 6528 0 -1 12852
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_119
timestamp 1679999689
transform 1 0 9120 0 -1 12852
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_120
timestamp 1679999689
transform 1 0 8256 0 1 77868
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_121
timestamp 1679999689
transform -1 0 4800 0 -1 14364
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_122
timestamp 1679999689
transform -1 0 14016 0 -1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_123
timestamp 1679999689
transform -1 0 14016 0 1 756
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_124
timestamp 1679999689
transform 1 0 13056 0 1 20412
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_125
timestamp 1679999689
transform 1 0 11616 0 -1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_126
timestamp 1679999689
transform 1 0 18240 0 1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_127
timestamp 1679999689
transform 1 0 12960 0 1 30996
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_128
timestamp 1679999689
transform 1 0 15552 0 1 27972
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_129
timestamp 1679999689
transform -1 0 17760 0 1 18900
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_130
timestamp 1679999689
transform 1 0 8160 0 1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_131
timestamp 1679999689
transform 1 0 1632 0 1 23436
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_132
timestamp 1679999689
transform 1 0 19680 0 -1 43092
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_133
timestamp 1679999689
transform 1 0 14016 0 1 756
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_134
timestamp 1679999689
transform 1 0 15072 0 -1 2268
box -48 -56 336 834
use sg13g2_buf_8  clkbuf_0_Tile_X0Y1_UserCLK
timestamp 1676451365
transform -1 0 10272 0 -1 61236
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_Tile_X0Y1_UserCLK
timestamp 1676451365
transform -1 0 7584 0 -1 50652
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_1__f_Tile_X0Y1_UserCLK
timestamp 1676451365
transform 1 0 10560 0 1 68796
box -48 -56 1296 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 2496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 3168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 4512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 5184 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_49
timestamp 1679577901
transform 1 0 5856 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_53
timestamp 1677580104
transform 1 0 6240 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 7200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7872 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_77
timestamp 1679577901
transform 1 0 8544 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_81
timestamp 1677580104
transform 1 0 8928 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_87
timestamp 1679581782
transform 1 0 9504 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_94
timestamp 1677579658
transform 1 0 10176 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_99
timestamp 1679577901
transform 1 0 10656 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_107
timestamp 1677579658
transform 1 0 11424 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11904 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_119
timestamp 1679577901
transform 1 0 12576 0 1 756
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_157
timestamp 1679581782
transform 1 0 16224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_164
timestamp 1679581782
transform 1 0 16896 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_171
timestamp 1679577901
transform 1 0 17568 0 1 756
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_191
timestamp 1679581782
transform 1 0 19488 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_198
timestamp 1677580104
transform 1 0 20160 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 2496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 3168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 4512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_42
timestamp 1679577901
transform 1 0 5184 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_46
timestamp 1677579658
transform 1 0 5568 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_71
timestamp 1677579658
transform 1 0 7968 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_76
timestamp 1677579658
transform 1 0 8448 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_117
timestamp 1677580104
transform 1 0 12384 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_119
timestamp 1677579658
transform 1 0 12576 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_128
timestamp 1677580104
transform 1 0 13440 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_130
timestamp 1677579658
transform 1 0 13632 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_142
timestamp 1677580104
transform 1 0 14784 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_144
timestamp 1677579658
transform 1 0 14976 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_164
timestamp 1677580104
transform 1 0 16896 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_166
timestamp 1677579658
transform 1 0 17088 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_199
timestamp 1677579658
transform 1 0 20256 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 1824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679581782
transform 1 0 2496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679581782
transform 1 0 3168 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 4512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 5184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 5856 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_56
timestamp 1677580104
transform 1 0 6528 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_58
timestamp 1677579658
transform 1 0 6720 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679581782
transform 1 0 7200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 7872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1679581782
transform 1 0 8544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1679581782
transform 1 0 9216 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1679581782
transform 1 0 9888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1679581782
transform 1 0 10560 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_105
timestamp 1677579658
transform 1 0 11232 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_110
timestamp 1679581782
transform 1 0 11712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_117
timestamp 1679581782
transform 1 0 12384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_124
timestamp 1679581782
transform 1 0 13056 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_135
timestamp 1677580104
transform 1 0 14112 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_141
timestamp 1677580104
transform 1 0 14688 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_143
timestamp 1677579658
transform 1 0 14880 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_147
timestamp 1679581782
transform 1 0 15264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_154
timestamp 1679581782
transform 1 0 15936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_161
timestamp 1679581782
transform 1 0 16608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1679581782
transform 1 0 17280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_175
timestamp 1679581782
transform 1 0 17952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_182
timestamp 1679581782
transform 1 0 18624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_189
timestamp 1679581782
transform 1 0 19296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_196
timestamp 1679577901
transform 1 0 19968 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 1824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 2496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679581782
transform 1 0 3168 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1679581782
transform 1 0 3840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1679581782
transform 1 0 4512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679581782
transform 1 0 5184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_49
timestamp 1679577901
transform 1 0 5856 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_53
timestamp 1677580104
transform 1 0 6240 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_58
timestamp 1679581782
transform 1 0 6720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_65
timestamp 1679581782
transform 1 0 7392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_72
timestamp 1679581782
transform 1 0 8064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_79
timestamp 1679581782
transform 1 0 8736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_86
timestamp 1679581782
transform 1 0 9408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_93
timestamp 1679581782
transform 1 0 10080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_100
timestamp 1679581782
transform 1 0 10752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_107
timestamp 1679581782
transform 1 0 11424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_114
timestamp 1679581782
transform 1 0 12096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_121
timestamp 1679581782
transform 1 0 12768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_128
timestamp 1679581782
transform 1 0 13440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_135
timestamp 1679581782
transform 1 0 14112 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_142
timestamp 1677580104
transform 1 0 14784 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_147
timestamp 1679581782
transform 1 0 15264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_154
timestamp 1679581782
transform 1 0 15936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_161
timestamp 1679581782
transform 1 0 16608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_171
timestamp 1679581782
transform 1 0 17568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_178
timestamp 1679581782
transform 1 0 18240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_185
timestamp 1679581782
transform 1 0 18912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_192
timestamp 1679581782
transform 1 0 19584 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_199
timestamp 1677579658
transform 1 0 20256 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 2496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 3168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 3840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679581782
transform 1 0 4512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1679581782
transform 1 0 5184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_49
timestamp 1679577901
transform 1 0 5856 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_53
timestamp 1677580104
transform 1 0 6240 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_58
timestamp 1679581782
transform 1 0 6720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_65
timestamp 1679581782
transform 1 0 7392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_72
timestamp 1679581782
transform 1 0 8064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_79
timestamp 1679581782
transform 1 0 8736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_86
timestamp 1679581782
transform 1 0 9408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_93
timestamp 1679581782
transform 1 0 10080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_100
timestamp 1679581782
transform 1 0 10752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_107
timestamp 1679581782
transform 1 0 11424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_114
timestamp 1679581782
transform 1 0 12096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_121
timestamp 1679581782
transform 1 0 12768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_128
timestamp 1679581782
transform 1 0 13440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_135
timestamp 1679581782
transform 1 0 14112 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_142
timestamp 1677580104
transform 1 0 14784 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_147
timestamp 1679581782
transform 1 0 15264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_154
timestamp 1679581782
transform 1 0 15936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_161
timestamp 1679581782
transform 1 0 16608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_171
timestamp 1679581782
transform 1 0 17568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_178
timestamp 1679581782
transform 1 0 18240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_185
timestamp 1679581782
transform 1 0 18912 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_192
timestamp 1679581782
transform 1 0 19584 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_199
timestamp 1677579658
transform 1 0 20256 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679581782
transform 1 0 1824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1679581782
transform 1 0 2496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1679581782
transform 1 0 3168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1679581782
transform 1 0 3840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1679581782
transform 1 0 4512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_42
timestamp 1679581782
transform 1 0 5184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_49
timestamp 1679577901
transform 1 0 5856 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_53
timestamp 1677580104
transform 1 0 6240 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_58
timestamp 1679581782
transform 1 0 6720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_65
timestamp 1679581782
transform 1 0 7392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_72
timestamp 1679581782
transform 1 0 8064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_79
timestamp 1679581782
transform 1 0 8736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_86
timestamp 1679581782
transform 1 0 9408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_93
timestamp 1679581782
transform 1 0 10080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_100
timestamp 1679581782
transform 1 0 10752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_107
timestamp 1679581782
transform 1 0 11424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_114
timestamp 1679581782
transform 1 0 12096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_121
timestamp 1679581782
transform 1 0 12768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_128
timestamp 1679581782
transform 1 0 13440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_135
timestamp 1679581782
transform 1 0 14112 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_142
timestamp 1677580104
transform 1 0 14784 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_147
timestamp 1679581782
transform 1 0 15264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_154
timestamp 1679581782
transform 1 0 15936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_161
timestamp 1679581782
transform 1 0 16608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_171
timestamp 1679581782
transform 1 0 17568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_178
timestamp 1679581782
transform 1 0 18240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_185
timestamp 1679581782
transform 1 0 18912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_192
timestamp 1679581782
transform 1 0 19584 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_199
timestamp 1677579658
transform 1 0 20256 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 2496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 3168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 3840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 4512 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679581782
transform 1 0 5184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_49
timestamp 1679577901
transform 1 0 5856 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_53
timestamp 1677580104
transform 1 0 6240 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_58
timestamp 1679581782
transform 1 0 6720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_65
timestamp 1679581782
transform 1 0 7392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_72
timestamp 1679581782
transform 1 0 8064 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_79
timestamp 1679581782
transform 1 0 8736 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_86
timestamp 1679581782
transform 1 0 9408 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_93
timestamp 1679581782
transform 1 0 10080 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_100
timestamp 1679581782
transform 1 0 10752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_107
timestamp 1679581782
transform 1 0 11424 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_114
timestamp 1679581782
transform 1 0 12096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_121
timestamp 1679577901
transform 1 0 12768 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_125
timestamp 1677580104
transform 1 0 13152 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_147
timestamp 1679581782
transform 1 0 15264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_154
timestamp 1679581782
transform 1 0 15936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_161
timestamp 1679581782
transform 1 0 16608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_171
timestamp 1679581782
transform 1 0 17568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_178
timestamp 1679581782
transform 1 0 18240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_185
timestamp 1679577901
transform 1 0 18912 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_189
timestamp 1677579658
transform 1 0 19296 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_195
timestamp 1679577901
transform 1 0 19872 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_199
timestamp 1677579658
transform 1 0 20256 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 2496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 3168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 4512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 5184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_49
timestamp 1679577901
transform 1 0 5856 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_53
timestamp 1677580104
transform 1 0 6240 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_58
timestamp 1679581782
transform 1 0 6720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_65
timestamp 1679581782
transform 1 0 7392 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_72
timestamp 1677580104
transform 1 0 8064 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_74
timestamp 1677579658
transform 1 0 8256 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_92
timestamp 1677579658
transform 1 0 9984 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_97
timestamp 1679581782
transform 1 0 10464 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_104
timestamp 1677580104
transform 1 0 11136 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_106
timestamp 1677579658
transform 1 0 11328 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_111
timestamp 1679581782
transform 1 0 11808 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_118
timestamp 1677580104
transform 1 0 12480 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_137
timestamp 1679581782
transform 1 0 14304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679581782
transform 1 0 16608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_171
timestamp 1679581782
transform 1 0 17568 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_178
timestamp 1679577901
transform 1 0 18240 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_199
timestamp 1677579658
transform 1 0 20256 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 1824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679581782
transform 1 0 2496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_21
timestamp 1679581782
transform 1 0 3168 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_28
timestamp 1677580104
transform 1 0 3840 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_30
timestamp 1677579658
transform 1 0 4032 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_36
timestamp 1679581782
transform 1 0 4608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_43
timestamp 1679581782
transform 1 0 5280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_50
timestamp 1679577901
transform 1 0 5952 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_54
timestamp 1677579658
transform 1 0 6336 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_93
timestamp 1679581782
transform 1 0 10080 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_100
timestamp 1677579658
transform 1 0 10752 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_139
timestamp 1679577901
transform 1 0 14496 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_143
timestamp 1677579658
transform 1 0 14880 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_190
timestamp 1677579658
transform 1 0 19392 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_7
timestamp 1679581782
transform 1 0 1824 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_14
timestamp 1679577901
transform 1 0 2496 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_33
timestamp 1677580104
transform 1 0 4320 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_35
timestamp 1677579658
transform 1 0 4512 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_41
timestamp 1679581782
transform 1 0 5088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_48
timestamp 1679577901
transform 1 0 5760 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_9_58
timestamp 1679577901
transform 1 0 6720 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_79
timestamp 1677579658
transform 1 0 8736 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_97
timestamp 1679577901
transform 1 0 10464 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_9_122
timestamp 1679577901
transform 1 0 12864 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_126
timestamp 1677579658
transform 1 0 13248 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_147
timestamp 1679581782
transform 1 0 15264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_154
timestamp 1679581782
transform 1 0 15936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_161
timestamp 1679581782
transform 1 0 16608 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_188
timestamp 1677580104
transform 1 0 19200 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 1152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_24
timestamp 1679577901
transform 1 0 3456 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_58
timestamp 1677579658
transform 1 0 6720 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_76
timestamp 1677579658
transform 1 0 8448 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_98
timestamp 1677579658
transform 1 0 10560 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_121
timestamp 1679577901
transform 1 0 12768 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_125
timestamp 1677579658
transform 1 0 13152 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_143
timestamp 1677579658
transform 1 0 14880 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_150
timestamp 1679581782
transform 1 0 15552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_157
timestamp 1679577901
transform 1 0 16224 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_161
timestamp 1677580104
transform 1 0 16608 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_0
timestamp 1679577901
transform 1 0 1152 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_4  FILLER_11_21
timestamp 1679577901
transform 1 0 3168 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_43
timestamp 1677580104
transform 1 0 5280 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_55
timestamp 1677579658
transform 1 0 6432 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_80
timestamp 1677580104
transform 1 0 8832 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_82
timestamp 1677579658
transform 1 0 9024 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_86
timestamp 1677580104
transform 1 0 9408 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_105
timestamp 1679577901
transform 1 0 11232 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_126
timestamp 1677580104
transform 1 0 13248 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_128
timestamp 1677579658
transform 1 0 13440 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_134
timestamp 1677580104
transform 1 0 14016 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_164
timestamp 1679577901
transform 1 0 16896 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_48
timestamp 1677580104
transform 1 0 5760 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_55
timestamp 1677579658
transform 1 0 6432 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_59
timestamp 1677579658
transform 1 0 6816 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_65
timestamp 1677579658
transform 1 0 7392 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_91
timestamp 1677579658
transform 1 0 9888 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_123
timestamp 1677580104
transform 1 0 12960 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_125
timestamp 1677579658
transform 1 0 13152 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_148
timestamp 1677580104
transform 1 0 15360 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_150
timestamp 1677579658
transform 1 0 15552 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_171
timestamp 1677579658
transform 1 0 17568 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_199
timestamp 1677579658
transform 1 0 20256 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_34
timestamp 1677579658
transform 1 0 4416 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_38
timestamp 1677580104
transform 1 0 4800 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_40
timestamp 1677579658
transform 1 0 4992 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_79
timestamp 1679577901
transform 1 0 8736 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_146
timestamp 1677580104
transform 1 0 15168 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_177
timestamp 1677579658
transform 1 0 18144 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_199
timestamp 1677579658
transform 1 0 20256 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_38
timestamp 1677579658
transform 1 0 4800 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_63
timestamp 1677580104
transform 1 0 7200 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_65
timestamp 1677579658
transform 1 0 7392 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_86
timestamp 1679577901
transform 1 0 9408 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_117
timestamp 1679581782
transform 1 0 12384 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_124
timestamp 1679581782
transform 1 0 13056 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_131
timestamp 1677579658
transform 1 0 13728 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_171
timestamp 1677580104
transform 1 0 17568 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_173
timestamp 1677579658
transform 1 0 17760 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_179
timestamp 1677580104
transform 1 0 18336 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_181
timestamp 1677579658
transform 1 0 18528 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_199
timestamp 1677579658
transform 1 0 20256 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_32
timestamp 1677580104
transform 1 0 4224 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_34
timestamp 1677579658
transform 1 0 4416 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_45
timestamp 1677579658
transform 1 0 5472 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_86
timestamp 1679581782
transform 1 0 9408 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_93
timestamp 1677579658
transform 1 0 10080 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_120
timestamp 1677580104
transform 1 0 12672 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_122
timestamp 1677579658
transform 1 0 12864 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_140
timestamp 1677580104
transform 1 0 14592 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_176
timestamp 1677580104
transform 1 0 18048 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_178
timestamp 1677579658
transform 1 0 18240 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_0
timestamp 1679577901
transform 1 0 1152 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_4
timestamp 1677579658
transform 1 0 1536 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_22
timestamp 1677580104
transform 1 0 3264 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_24
timestamp 1677579658
transform 1 0 3456 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_38
timestamp 1677580104
transform 1 0 4800 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_111
timestamp 1679581782
transform 1 0 11808 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_118
timestamp 1677580104
transform 1 0 12480 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_120
timestamp 1677579658
transform 1 0 12672 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_142
timestamp 1677580104
transform 1 0 14784 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_144
timestamp 1677579658
transform 1 0 14976 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_165
timestamp 1677580104
transform 1 0 16992 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_167
timestamp 1677579658
transform 1 0 17184 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_185
timestamp 1677579658
transform 1 0 18912 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_0
timestamp 1679577901
transform 1 0 1152 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_4
timestamp 1677579658
transform 1 0 1536 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_22
timestamp 1677580104
transform 1 0 3264 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_46
timestamp 1677580104
transform 1 0 5568 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_90
timestamp 1677579658
transform 1 0 9792 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_125
timestamp 1677579658
transform 1 0 13152 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_147
timestamp 1679577901
transform 1 0 15264 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_177
timestamp 1677580104
transform 1 0 18144 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_17
timestamp 1677580104
transform 1 0 2784 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_51
timestamp 1679577901
transform 1 0 6048 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_55
timestamp 1677580104
transform 1 0 6432 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_74
timestamp 1677579658
transform 1 0 8256 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_115
timestamp 1679581782
transform 1 0 12192 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_122
timestamp 1679577901
transform 1 0 12864 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_198
timestamp 1677580104
transform 1 0 20160 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_19_0
timestamp 1679577901
transform 1 0 1152 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_21
timestamp 1677580104
transform 1 0 3168 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_48
timestamp 1679581782
transform 1 0 5760 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_55
timestamp 1677580104
transform 1 0 6432 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_57
timestamp 1677579658
transform 1 0 6624 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_79
timestamp 1677579658
transform 1 0 8736 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_101
timestamp 1679581782
transform 1 0 10848 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_125
timestamp 1677580104
transform 1 0 13152 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_147
timestamp 1677580104
transform 1 0 15264 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_0
timestamp 1679581782
transform 1 0 1152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_7
timestamp 1679577901
transform 1 0 1824 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_33
timestamp 1677579658
transform 1 0 4320 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_44
timestamp 1677579658
transform 1 0 5376 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_62
timestamp 1679577901
transform 1 0 7104 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_66
timestamp 1677579658
transform 1 0 7488 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_84
timestamp 1677579658
transform 1 0 9216 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_102
timestamp 1679581782
transform 1 0 10944 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_109
timestamp 1679581782
transform 1 0 11616 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_116
timestamp 1679577901
transform 1 0 12288 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_120
timestamp 1677579658
transform 1 0 12672 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_126
timestamp 1677579658
transform 1 0 13248 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_144
timestamp 1677580104
transform 1 0 14976 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_179
timestamp 1677579658
transform 1 0 18336 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_198
timestamp 1677580104
transform 1 0 20160 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_45
timestamp 1677580104
transform 1 0 5472 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_47
timestamp 1677579658
transform 1 0 5664 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_103
timestamp 1677580104
transform 1 0 11040 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_143
timestamp 1677580104
transform 1 0 14880 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_162
timestamp 1677580104
transform 1 0 16704 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_168
timestamp 1677580104
transform 1 0 17280 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_170
timestamp 1677579658
transform 1 0 17472 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_0
timestamp 1679577901
transform 1 0 1152 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_4
timestamp 1677580104
transform 1 0 1536 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_32
timestamp 1677579658
transform 1 0 4224 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_81
timestamp 1677580104
transform 1 0 8928 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_153
timestamp 1677580104
transform 1 0 15840 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_155
timestamp 1677579658
transform 1 0 16032 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_198
timestamp 1677580104
transform 1 0 20160 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_17
timestamp 1677580104
transform 1 0 2784 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_57
timestamp 1677579658
transform 1 0 6624 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_75
timestamp 1677580104
transform 1 0 8352 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_77
timestamp 1677579658
transform 1 0 8544 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_95
timestamp 1677580104
transform 1 0 10272 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_23_102
timestamp 1679577901
transform 1 0 10944 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_123
timestamp 1677580104
transform 1 0 12960 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_163
timestamp 1677579658
transform 1 0 16800 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_17
timestamp 1677580104
transform 1 0 2784 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_36
timestamp 1677579658
transform 1 0 4608 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_54
timestamp 1679577901
transform 1 0 6336 0 1 18900
box -48 -56 432 834
use sg13g2_decap_4  FILLER_24_75
timestamp 1679577901
transform 1 0 8352 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_96
timestamp 1677579658
transform 1 0 10368 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_105
timestamp 1679577901
transform 1 0 11232 0 1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_24_139
timestamp 1679581782
transform 1 0 14496 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_146
timestamp 1679577901
transform 1 0 15168 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_150
timestamp 1677580104
transform 1 0 15552 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_169
timestamp 1677579658
transform 1 0 17376 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_190
timestamp 1677580104
transform 1 0 19392 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_197
timestamp 1677580104
transform 1 0 20064 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_199
timestamp 1677579658
transform 1 0 20256 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_55
timestamp 1679581782
transform 1 0 6432 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_65
timestamp 1679577901
transform 1 0 7392 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_87
timestamp 1677579658
transform 1 0 9504 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_127
timestamp 1677579658
transform 1 0 13344 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_145
timestamp 1679581782
transform 1 0 15072 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_199
timestamp 1677579658
transform 1 0 20256 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_26_38
timestamp 1679577901
transform 1 0 4800 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_42
timestamp 1677580104
transform 1 0 5184 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_78
timestamp 1679581782
transform 1 0 8640 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_85
timestamp 1677580104
transform 1 0 9312 0 1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_117
timestamp 1677580104
transform 1 0 12384 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_144
timestamp 1677579658
transform 1 0 14976 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_182
timestamp 1677579658
transform 1 0 18624 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_0
timestamp 1677580104
transform 1 0 1152 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_2
timestamp 1677579658
transform 1 0 1344 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_20
timestamp 1677580104
transform 1 0 3072 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_22
timestamp 1677579658
transform 1 0 3264 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_38
timestamp 1679577901
transform 1 0 4800 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_42
timestamp 1677580104
transform 1 0 5184 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_93
timestamp 1679581782
transform 1 0 10080 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_100
timestamp 1677580104
transform 1 0 10752 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_107
timestamp 1679581782
transform 1 0 11424 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_114
timestamp 1679577901
transform 1 0 12096 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_135
timestamp 1677580104
transform 1 0 14112 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_137
timestamp 1677579658
transform 1 0 14304 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_193
timestamp 1677579658
transform 1 0 19680 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_199
timestamp 1677579658
transform 1 0 20256 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_17
timestamp 1677579658
transform 1 0 2784 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_39
timestamp 1677580104
transform 1 0 4896 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_41
timestamp 1677579658
transform 1 0 5088 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_97
timestamp 1679577901
transform 1 0 10464 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_149
timestamp 1677579658
transform 1 0 15456 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_198
timestamp 1677580104
transform 1 0 20160 0 1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_29_0
timestamp 1679577901
transform 1 0 1152 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_4
timestamp 1677579658
transform 1 0 1536 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_32
timestamp 1677580104
transform 1 0 4224 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_51
timestamp 1677580104
transform 1 0 6048 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_53
timestamp 1677579658
transform 1 0 6240 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_64
timestamp 1677579658
transform 1 0 7296 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_75
timestamp 1677580104
transform 1 0 8352 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_77
timestamp 1677579658
transform 1 0 8544 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_105
timestamp 1677579658
transform 1 0 11232 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_144
timestamp 1677580104
transform 1 0 14976 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_158
timestamp 1677579658
transform 1 0 16320 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_199
timestamp 1677579658
transform 1 0 20256 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_0
timestamp 1677580104
transform 1 0 1152 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_30_45
timestamp 1679577901
transform 1 0 5472 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_49
timestamp 1677579658
transform 1 0 5856 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_67
timestamp 1677580104
transform 1 0 7584 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_69
timestamp 1677579658
transform 1 0 7776 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_112
timestamp 1679581782
transform 1 0 11904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_119
timestamp 1679577901
transform 1 0 12576 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_123
timestamp 1677580104
transform 1 0 12960 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_142
timestamp 1679581782
transform 1 0 14784 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_149
timestamp 1677579658
transform 1 0 15456 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_174
timestamp 1677580104
transform 1 0 17856 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_198
timestamp 1677580104
transform 1 0 20160 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_0
timestamp 1677579658
transform 1 0 1152 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_25
timestamp 1677579658
transform 1 0 3552 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_47
timestamp 1679577901
transform 1 0 5664 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_89
timestamp 1677580104
transform 1 0 9696 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_130
timestamp 1677579658
transform 1 0 13632 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_144
timestamp 1677580104
transform 1 0 14976 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_25
timestamp 1677580104
transform 1 0 3552 0 1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_32_53
timestamp 1679577901
transform 1 0 6240 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_57
timestamp 1677580104
transform 1 0 6624 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_80
timestamp 1679581782
transform 1 0 8832 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_87
timestamp 1679577901
transform 1 0 9504 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_91
timestamp 1677580104
transform 1 0 9888 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_131
timestamp 1677580104
transform 1 0 13728 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_153
timestamp 1677579658
transform 1 0 15840 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_198
timestamp 1677580104
transform 1 0 20160 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_42
timestamp 1677580104
transform 1 0 5184 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_95
timestamp 1679581782
transform 1 0 10272 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_102
timestamp 1679581782
transform 1 0 10944 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_109
timestamp 1679581782
transform 1 0 11616 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_116
timestamp 1677579658
transform 1 0 12288 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_148
timestamp 1677580104
transform 1 0 15360 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_198
timestamp 1677580104
transform 1 0 20160 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_42
timestamp 1677579658
transform 1 0 5184 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_48
timestamp 1677580104
transform 1 0 5760 0 1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_34_88
timestamp 1679577901
transform 1 0 9600 0 1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_34_109
timestamp 1679581782
transform 1 0 11616 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_116
timestamp 1679577901
transform 1 0 12288 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_187
timestamp 1677580104
transform 1 0 19104 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_197
timestamp 1677580104
transform 1 0 20064 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_199
timestamp 1677579658
transform 1 0 20256 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_0
timestamp 1679577901
transform 1 0 1152 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_4
timestamp 1677579658
transform 1 0 1536 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_130
timestamp 1677580104
transform 1 0 13632 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_132
timestamp 1677579658
transform 1 0 13824 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_157
timestamp 1677580104
transform 1 0 16224 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_164
timestamp 1677579658
transform 1 0 16896 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_198
timestamp 1677580104
transform 1 0 20160 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_36_0
timestamp 1679577901
transform 1 0 1152 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_4
timestamp 1677579658
transform 1 0 1536 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_8
timestamp 1679581782
transform 1 0 1920 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_15
timestamp 1677580104
transform 1 0 2592 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_17
timestamp 1677579658
transform 1 0 2784 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_39
timestamp 1677579658
transform 1 0 4896 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_78
timestamp 1679581782
transform 1 0 8640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_85
timestamp 1679581782
transform 1 0 9312 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_92
timestamp 1677580104
transform 1 0 9984 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_199
timestamp 1677579658
transform 1 0 20256 0 1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_37_0
timestamp 1679577901
transform 1 0 1152 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_4
timestamp 1677579658
transform 1 0 1536 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_37_30
timestamp 1679577901
transform 1 0 4032 0 -1 29484
box -48 -56 432 834
use sg13g2_decap_8  FILLER_37_82
timestamp 1679581782
transform 1 0 9024 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_89
timestamp 1679577901
transform 1 0 9696 0 -1 29484
box -48 -56 432 834
use sg13g2_decap_4  FILLER_37_114
timestamp 1679577901
transform 1 0 12096 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_118
timestamp 1677580104
transform 1 0 12480 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_147
timestamp 1677580104
transform 1 0 15264 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_149
timestamp 1677579658
transform 1 0 15456 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_37_153
timestamp 1679577901
transform 1 0 15840 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_157
timestamp 1677579658
transform 1 0 16224 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_38_0
timestamp 1679577901
transform 1 0 1152 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_4
timestamp 1677579658
transform 1 0 1536 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_38_57
timestamp 1679577901
transform 1 0 6624 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_61
timestamp 1677580104
transform 1 0 7008 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_80
timestamp 1677580104
transform 1 0 8832 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_99
timestamp 1677580104
transform 1 0 10656 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_101
timestamp 1677579658
transform 1 0 10848 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_119
timestamp 1679581782
transform 1 0 12576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_126
timestamp 1679577901
transform 1 0 13248 0 1 29484
box -48 -56 432 834
use sg13g2_decap_4  FILLER_38_156
timestamp 1679577901
transform 1 0 16128 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_160
timestamp 1677580104
transform 1 0 16512 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_191
timestamp 1677579658
transform 1 0 19488 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_39_0
timestamp 1679577901
transform 1 0 1152 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_4
timestamp 1677579658
transform 1 0 1536 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_8
timestamp 1679581782
transform 1 0 1920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_15
timestamp 1679581782
transform 1 0 2592 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_65
timestamp 1677579658
transform 1 0 7392 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_87
timestamp 1679581782
transform 1 0 9504 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_94
timestamp 1677580104
transform 1 0 10176 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_96
timestamp 1677579658
transform 1 0 10368 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_118
timestamp 1679581782
transform 1 0 12480 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_125
timestamp 1677579658
transform 1 0 13152 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_160
timestamp 1677580104
transform 1 0 16512 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_170
timestamp 1677580104
transform 1 0 17472 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_172
timestamp 1677579658
transform 1 0 17664 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_198
timestamp 1677580104
transform 1 0 20160 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 1152 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_7
timestamp 1679577901
transform 1 0 1824 0 1 30996
box -48 -56 432 834
use sg13g2_decap_4  FILLER_40_118
timestamp 1679577901
transform 1 0 12480 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_122
timestamp 1677579658
transform 1 0 12864 0 1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_40_143
timestamp 1679577901
transform 1 0 14880 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_147
timestamp 1677580104
transform 1 0 15264 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_187
timestamp 1677580104
transform 1 0 19104 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_197
timestamp 1677580104
transform 1 0 20064 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_199
timestamp 1677579658
transform 1 0 20256 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_42
timestamp 1679581782
transform 1 0 5184 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_49
timestamp 1679581782
transform 1 0 5856 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_56
timestamp 1679581782
transform 1 0 6528 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_63
timestamp 1679577901
transform 1 0 7200 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_41_67
timestamp 1677579658
transform 1 0 7584 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_73
timestamp 1677580104
transform 1 0 8160 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_92
timestamp 1677579658
transform 1 0 9984 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_110
timestamp 1677580104
transform 1 0 11712 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_115
timestamp 1677580104
transform 1 0 12192 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_122
timestamp 1677580104
transform 1 0 12864 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_42_85
timestamp 1679577901
transform 1 0 9312 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_89
timestamp 1677580104
transform 1 0 9696 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_146
timestamp 1679581782
transform 1 0 15168 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_153
timestamp 1679581782
transform 1 0 15840 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_20
timestamp 1677579658
transform 1 0 3072 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_85
timestamp 1677579658
transform 1 0 9312 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_91
timestamp 1679581782
transform 1 0 9888 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_98
timestamp 1677580104
transform 1 0 10560 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_155
timestamp 1679581782
transform 1 0 16032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_162
timestamp 1679577901
transform 1 0 16704 0 -1 34020
box -48 -56 432 834
use sg13g2_decap_4  FILLER_43_183
timestamp 1679577901
transform 1 0 18720 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_187
timestamp 1677580104
transform 1 0 19104 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_197
timestamp 1677580104
transform 1 0 20064 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_199
timestamp 1677579658
transform 1 0 20256 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_119
timestamp 1677579658
transform 1 0 12576 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_158
timestamp 1677580104
transform 1 0 16320 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_160
timestamp 1677579658
transform 1 0 16512 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_165
timestamp 1679577901
transform 1 0 16992 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_198
timestamp 1677580104
transform 1 0 20160 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 1152 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_11
timestamp 1677580104
transform 1 0 2208 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_34
timestamp 1677580104
transform 1 0 4416 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_36
timestamp 1677579658
transform 1 0 4608 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_78
timestamp 1677580104
transform 1 0 8640 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_80
timestamp 1677579658
transform 1 0 8832 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_119
timestamp 1677580104
transform 1 0 12576 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_141
timestamp 1677580104
transform 1 0 14688 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_160
timestamp 1679581782
transform 1 0 16512 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_187
timestamp 1677580104
transform 1 0 19104 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_189
timestamp 1677579658
transform 1 0 19296 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_198
timestamp 1677580104
transform 1 0 20160 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_4  FILLER_46_38
timestamp 1679577901
transform 1 0 4800 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_94
timestamp 1677579658
transform 1 0 10176 0 1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_116
timestamp 1677579658
transform 1 0 12288 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_138
timestamp 1679581782
transform 1 0 14400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_162
timestamp 1679577901
transform 1 0 16704 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_166
timestamp 1677579658
transform 1 0 17088 0 1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_199
timestamp 1677579658
transform 1 0 20256 0 1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_47_17
timestamp 1679577901
transform 1 0 2784 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_21
timestamp 1677579658
transform 1 0 3168 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_4  FILLER_47_39
timestamp 1679577901
transform 1 0 4896 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_43
timestamp 1677580104
transform 1 0 5280 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_62
timestamp 1677580104
transform 1 0 7104 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_84
timestamp 1677580104
transform 1 0 9216 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_86
timestamp 1677579658
transform 1 0 9408 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_95
timestamp 1677580104
transform 1 0 10272 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_166
timestamp 1677579658
transform 1 0 17088 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_170
timestamp 1679581782
transform 1 0 17472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_177
timestamp 1679581782
transform 1 0 18144 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_184
timestamp 1677579658
transform 1 0 18816 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_188
timestamp 1679581782
transform 1 0 19200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_195
timestamp 1679577901
transform 1 0 19872 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_199
timestamp 1677579658
transform 1 0 20256 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 1152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_7
timestamp 1679577901
transform 1 0 1824 0 1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_48_11
timestamp 1677580104
transform 1 0 2208 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_84
timestamp 1677579658
transform 1 0 9216 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_90
timestamp 1677580104
transform 1 0 9792 0 1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_48_95
timestamp 1677580104
transform 1 0 10272 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_97
timestamp 1677579658
transform 1 0 10464 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_132
timestamp 1679581782
transform 1 0 13824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_139
timestamp 1679581782
transform 1 0 14496 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_170
timestamp 1679581782
transform 1 0 17472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_177
timestamp 1679581782
transform 1 0 18144 0 1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_184
timestamp 1677579658
transform 1 0 18816 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_38
timestamp 1679581782
transform 1 0 4800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_45
timestamp 1679577901
transform 1 0 5472 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_2  FILLER_49_49
timestamp 1677580104
transform 1 0 5856 0 -1 38556
box -48 -56 240 834
use sg13g2_decap_4  FILLER_49_76
timestamp 1679577901
transform 1 0 8448 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_80
timestamp 1677579658
transform 1 0 8832 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_4  FILLER_49_84
timestamp 1679577901
transform 1 0 9216 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_113
timestamp 1677579658
transform 1 0 12000 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_4  FILLER_49_135
timestamp 1679577901
transform 1 0 14112 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_139
timestamp 1677579658
transform 1 0 14496 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_160
timestamp 1679581782
transform 1 0 16512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_170
timestamp 1679581782
transform 1 0 17472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_177
timestamp 1679577901
transform 1 0 18144 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_8  FILLER_50_0
timestamp 1679581782
transform 1 0 1152 0 1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_50_7
timestamp 1679577901
transform 1 0 1824 0 1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_50_11
timestamp 1677579658
transform 1 0 2208 0 1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_50_33
timestamp 1679581782
transform 1 0 4320 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_40
timestamp 1679581782
transform 1 0 4992 0 1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_50_98
timestamp 1679577901
transform 1 0 10560 0 1 38556
box -48 -56 432 834
use sg13g2_decap_8  FILLER_50_160
timestamp 1679581782
transform 1 0 16512 0 1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_50_184
timestamp 1677579658
transform 1 0 18816 0 1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_51_17
timestamp 1679581782
transform 1 0 2784 0 -1 40068
box -48 -56 720 834
use sg13g2_fill_2  FILLER_51_24
timestamp 1677580104
transform 1 0 3456 0 -1 40068
box -48 -56 240 834
use sg13g2_decap_4  FILLER_51_47
timestamp 1679577901
transform 1 0 5664 0 -1 40068
box -48 -56 432 834
use sg13g2_fill_2  FILLER_51_51
timestamp 1677580104
transform 1 0 6048 0 -1 40068
box -48 -56 240 834
use sg13g2_decap_8  FILLER_51_74
timestamp 1679581782
transform 1 0 8256 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_105
timestamp 1679581782
transform 1 0 11232 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_4  FILLER_51_112
timestamp 1679577901
transform 1 0 11904 0 -1 40068
box -48 -56 432 834
use sg13g2_fill_2  FILLER_51_137
timestamp 1677580104
transform 1 0 14304 0 -1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_51_139
timestamp 1677579658
transform 1 0 14496 0 -1 40068
box -48 -56 144 834
use sg13g2_decap_8  FILLER_51_160
timestamp 1679581782
transform 1 0 16512 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_170
timestamp 1679581782
transform 1 0 17472 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_177
timestamp 1679581782
transform 1 0 18144 0 -1 40068
box -48 -56 720 834
use sg13g2_fill_1  FILLER_51_184
timestamp 1677579658
transform 1 0 18816 0 -1 40068
box -48 -56 144 834
use sg13g2_decap_4  FILLER_51_196
timestamp 1679577901
transform 1 0 19968 0 -1 40068
box -48 -56 432 834
use sg13g2_decap_8  FILLER_52_0
timestamp 1679581782
transform 1 0 1152 0 1 40068
box -48 -56 720 834
use sg13g2_fill_2  FILLER_52_78
timestamp 1677580104
transform 1 0 8640 0 1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_52_80
timestamp 1677579658
transform 1 0 8832 0 1 40068
box -48 -56 144 834
use sg13g2_decap_8  FILLER_52_84
timestamp 1679581782
transform 1 0 9216 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_91
timestamp 1679581782
transform 1 0 9888 0 1 40068
box -48 -56 720 834
use sg13g2_fill_1  FILLER_52_98
timestamp 1677579658
transform 1 0 10560 0 1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_52_116
timestamp 1677580104
transform 1 0 12288 0 1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_52_118
timestamp 1677579658
transform 1 0 12480 0 1 40068
box -48 -56 144 834
use sg13g2_decap_8  FILLER_52_160
timestamp 1679581782
transform 1 0 16512 0 1 40068
box -48 -56 720 834
use sg13g2_fill_2  FILLER_52_170
timestamp 1677580104
transform 1 0 17472 0 1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_52_172
timestamp 1677579658
transform 1 0 17664 0 1 40068
box -48 -56 144 834
use sg13g2_decap_8  FILLER_52_177
timestamp 1679581782
transform 1 0 18144 0 1 40068
box -48 -56 720 834
use sg13g2_fill_1  FILLER_52_184
timestamp 1677579658
transform 1 0 18816 0 1 40068
box -48 -56 144 834
use sg13g2_decap_8  FILLER_52_193
timestamp 1679581782
transform 1 0 19680 0 1 40068
box -48 -56 720 834
use sg13g2_decap_4  FILLER_53_0
timestamp 1679577901
transform 1 0 1152 0 -1 41580
box -48 -56 432 834
use sg13g2_fill_2  FILLER_53_4
timestamp 1677580104
transform 1 0 1536 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_2  FILLER_53_23
timestamp 1677580104
transform 1 0 3360 0 -1 41580
box -48 -56 240 834
use sg13g2_decap_8  FILLER_53_46
timestamp 1679581782
transform 1 0 5568 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_4  FILLER_53_53
timestamp 1679577901
transform 1 0 6240 0 -1 41580
box -48 -56 432 834
use sg13g2_fill_1  FILLER_53_57
timestamp 1677579658
transform 1 0 6624 0 -1 41580
box -48 -56 144 834
use sg13g2_decap_8  FILLER_53_96
timestamp 1679581782
transform 1 0 10368 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_4  FILLER_53_103
timestamp 1679577901
transform 1 0 11040 0 -1 41580
box -48 -56 432 834
use sg13g2_fill_2  FILLER_53_107
timestamp 1677580104
transform 1 0 11424 0 -1 41580
box -48 -56 240 834
use sg13g2_decap_8  FILLER_53_129
timestamp 1679581782
transform 1 0 13536 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_160
timestamp 1679581782
transform 1 0 16512 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_170
timestamp 1679581782
transform 1 0 17472 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_177
timestamp 1679581782
transform 1 0 18144 0 -1 41580
box -48 -56 720 834
use sg13g2_fill_1  FILLER_53_184
timestamp 1677579658
transform 1 0 18816 0 -1 41580
box -48 -56 144 834
use sg13g2_decap_4  FILLER_53_196
timestamp 1679577901
transform 1 0 19968 0 -1 41580
box -48 -56 432 834
use sg13g2_decap_8  FILLER_54_0
timestamp 1679581782
transform 1 0 1152 0 1 41580
box -48 -56 720 834
use sg13g2_decap_4  FILLER_54_7
timestamp 1679577901
transform 1 0 1824 0 1 41580
box -48 -56 432 834
use sg13g2_fill_2  FILLER_54_11
timestamp 1677580104
transform 1 0 2208 0 1 41580
box -48 -56 240 834
use sg13g2_decap_8  FILLER_54_51
timestamp 1679581782
transform 1 0 6048 0 1 41580
box -48 -56 720 834
use sg13g2_decap_4  FILLER_54_58
timestamp 1679577901
transform 1 0 6720 0 1 41580
box -48 -56 432 834
use sg13g2_fill_2  FILLER_54_62
timestamp 1677580104
transform 1 0 7104 0 1 41580
box -48 -56 240 834
use sg13g2_fill_2  FILLER_54_84
timestamp 1677580104
transform 1 0 9216 0 1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_54_86
timestamp 1677579658
transform 1 0 9408 0 1 41580
box -48 -56 144 834
use sg13g2_decap_4  FILLER_54_108
timestamp 1679577901
transform 1 0 11520 0 1 41580
box -48 -56 432 834
use sg13g2_fill_2  FILLER_54_112
timestamp 1677580104
transform 1 0 11904 0 1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_54_135
timestamp 1677579658
transform 1 0 14112 0 1 41580
box -48 -56 144 834
use sg13g2_decap_8  FILLER_54_178
timestamp 1679581782
transform 1 0 18240 0 1 41580
box -48 -56 720 834
use sg13g2_decap_4  FILLER_54_196
timestamp 1679577901
transform 1 0 19968 0 1 41580
box -48 -56 432 834
use sg13g2_fill_2  FILLER_55_0
timestamp 1677580104
transform 1 0 1152 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_55_40
timestamp 1677579658
transform 1 0 4992 0 -1 43092
box -48 -56 144 834
use sg13g2_decap_4  FILLER_55_75
timestamp 1679577901
transform 1 0 8352 0 -1 43092
box -48 -56 432 834
use sg13g2_fill_2  FILLER_55_79
timestamp 1677580104
transform 1 0 8736 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_2  FILLER_55_84
timestamp 1677580104
transform 1 0 9216 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_55_86
timestamp 1677579658
transform 1 0 9408 0 -1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_55_90
timestamp 1679581782
transform 1 0 9792 0 -1 43092
box -48 -56 720 834
use sg13g2_fill_2  FILLER_55_97
timestamp 1677580104
transform 1 0 10464 0 -1 43092
box -48 -56 240 834
use sg13g2_decap_4  FILLER_55_116
timestamp 1679577901
transform 1 0 12288 0 -1 43092
box -48 -56 432 834
use sg13g2_fill_2  FILLER_55_137
timestamp 1677580104
transform 1 0 14304 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_55_139
timestamp 1677579658
transform 1 0 14496 0 -1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_55_160
timestamp 1679581782
transform 1 0 16512 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_170
timestamp 1679581782
transform 1 0 17472 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_177
timestamp 1679581782
transform 1 0 18144 0 -1 43092
box -48 -56 720 834
use sg13g2_fill_1  FILLER_55_184
timestamp 1677579658
transform 1 0 18816 0 -1 43092
box -48 -56 144 834
use sg13g2_decap_4  FILLER_55_188
timestamp 1679577901
transform 1 0 19200 0 -1 43092
box -48 -56 432 834
use sg13g2_fill_1  FILLER_55_192
timestamp 1677579658
transform 1 0 19584 0 -1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_56_0
timestamp 1679581782
transform 1 0 1152 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_7
timestamp 1679581782
transform 1 0 1824 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_14
timestamp 1679581782
transform 1 0 2496 0 1 43092
box -48 -56 720 834
use sg13g2_decap_4  FILLER_56_21
timestamp 1679577901
transform 1 0 3168 0 1 43092
box -48 -56 432 834
use sg13g2_fill_2  FILLER_56_76
timestamp 1677580104
transform 1 0 8448 0 1 43092
box -48 -56 240 834
use sg13g2_decap_8  FILLER_56_95
timestamp 1679581782
transform 1 0 10272 0 1 43092
box -48 -56 720 834
use sg13g2_fill_2  FILLER_56_102
timestamp 1677580104
transform 1 0 10944 0 1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_56_104
timestamp 1677579658
transform 1 0 11136 0 1 43092
box -48 -56 144 834
use sg13g2_fill_2  FILLER_56_122
timestamp 1677580104
transform 1 0 12864 0 1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_56_139
timestamp 1677579658
transform 1 0 14496 0 1 43092
box -48 -56 144 834
use sg13g2_fill_1  FILLER_56_165
timestamp 1677579658
transform 1 0 16992 0 1 43092
box -48 -56 144 834
use sg13g2_fill_2  FILLER_56_183
timestamp 1677580104
transform 1 0 18720 0 1 43092
box -48 -56 240 834
use sg13g2_decap_8  FILLER_56_188
timestamp 1679581782
transform 1 0 19200 0 1 43092
box -48 -56 720 834
use sg13g2_decap_4  FILLER_56_195
timestamp 1679577901
transform 1 0 19872 0 1 43092
box -48 -56 432 834
use sg13g2_fill_1  FILLER_56_199
timestamp 1677579658
transform 1 0 20256 0 1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_57_0
timestamp 1679581782
transform 1 0 1152 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_7
timestamp 1679581782
transform 1 0 1824 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_4  FILLER_57_14
timestamp 1679577901
transform 1 0 2496 0 -1 44604
box -48 -56 432 834
use sg13g2_fill_2  FILLER_57_18
timestamp 1677580104
transform 1 0 2880 0 -1 44604
box -48 -56 240 834
use sg13g2_fill_1  FILLER_57_37
timestamp 1677579658
transform 1 0 4704 0 -1 44604
box -48 -56 144 834
use sg13g2_decap_4  FILLER_57_55
timestamp 1679577901
transform 1 0 6432 0 -1 44604
box -48 -56 432 834
use sg13g2_decap_8  FILLER_57_97
timestamp 1679581782
transform 1 0 10464 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_4  FILLER_57_104
timestamp 1679577901
transform 1 0 11136 0 -1 44604
box -48 -56 432 834
use sg13g2_fill_1  FILLER_57_108
timestamp 1677579658
transform 1 0 11520 0 -1 44604
box -48 -56 144 834
use sg13g2_fill_1  FILLER_57_139
timestamp 1677579658
transform 1 0 14496 0 -1 44604
box -48 -56 144 834
use sg13g2_fill_1  FILLER_57_165
timestamp 1677579658
transform 1 0 16992 0 -1 44604
box -48 -56 144 834
use sg13g2_decap_4  FILLER_57_171
timestamp 1679577901
transform 1 0 17568 0 -1 44604
box -48 -56 432 834
use sg13g2_fill_1  FILLER_57_175
timestamp 1677579658
transform 1 0 17952 0 -1 44604
box -48 -56 144 834
use sg13g2_fill_2  FILLER_57_197
timestamp 1677580104
transform 1 0 20064 0 -1 44604
box -48 -56 240 834
use sg13g2_fill_1  FILLER_57_199
timestamp 1677579658
transform 1 0 20256 0 -1 44604
box -48 -56 144 834
use sg13g2_decap_8  FILLER_58_0
timestamp 1679581782
transform 1 0 1152 0 1 44604
box -48 -56 720 834
use sg13g2_fill_1  FILLER_58_7
timestamp 1677579658
transform 1 0 1824 0 1 44604
box -48 -56 144 834
use sg13g2_fill_1  FILLER_58_25
timestamp 1677579658
transform 1 0 3552 0 1 44604
box -48 -56 144 834
use sg13g2_decap_4  FILLER_58_41
timestamp 1679577901
transform 1 0 5088 0 1 44604
box -48 -56 432 834
use sg13g2_fill_2  FILLER_58_75
timestamp 1677580104
transform 1 0 8352 0 1 44604
box -48 -56 240 834
use sg13g2_decap_8  FILLER_58_98
timestamp 1679581782
transform 1 0 10560 0 1 44604
box -48 -56 720 834
use sg13g2_fill_1  FILLER_58_105
timestamp 1677579658
transform 1 0 11232 0 1 44604
box -48 -56 144 834
use sg13g2_fill_2  FILLER_58_123
timestamp 1677580104
transform 1 0 12960 0 1 44604
box -48 -56 240 834
use sg13g2_decap_8  FILLER_58_150
timestamp 1679581782
transform 1 0 15552 0 1 44604
box -48 -56 720 834
use sg13g2_fill_1  FILLER_58_160
timestamp 1677579658
transform 1 0 16512 0 1 44604
box -48 -56 144 834
use sg13g2_fill_1  FILLER_58_199
timestamp 1677579658
transform 1 0 20256 0 1 44604
box -48 -56 144 834
use sg13g2_fill_2  FILLER_59_0
timestamp 1677580104
transform 1 0 1152 0 -1 46116
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_19
timestamp 1677580104
transform 1 0 2976 0 -1 46116
box -48 -56 240 834
use sg13g2_fill_1  FILLER_59_21
timestamp 1677579658
transform 1 0 3168 0 -1 46116
box -48 -56 144 834
use sg13g2_decap_4  FILLER_59_43
timestamp 1679577901
transform 1 0 5280 0 -1 46116
box -48 -56 432 834
use sg13g2_fill_2  FILLER_59_68
timestamp 1677580104
transform 1 0 7680 0 -1 46116
box -48 -56 240 834
use sg13g2_decap_4  FILLER_59_143
timestamp 1679577901
transform 1 0 14880 0 -1 46116
box -48 -56 432 834
use sg13g2_fill_1  FILLER_59_147
timestamp 1677579658
transform 1 0 15264 0 -1 46116
box -48 -56 144 834
use sg13g2_decap_4  FILLER_59_196
timestamp 1679577901
transform 1 0 19968 0 -1 46116
box -48 -56 432 834
use sg13g2_decap_8  FILLER_60_43
timestamp 1679581782
transform 1 0 5280 0 1 46116
box -48 -56 720 834
use sg13g2_fill_1  FILLER_60_50
timestamp 1677579658
transform 1 0 5952 0 1 46116
box -48 -56 144 834
use sg13g2_decap_8  FILLER_60_113
timestamp 1679581782
transform 1 0 12000 0 1 46116
box -48 -56 720 834
use sg13g2_decap_4  FILLER_60_141
timestamp 1679577901
transform 1 0 14688 0 1 46116
box -48 -56 432 834
use sg13g2_fill_2  FILLER_60_145
timestamp 1677580104
transform 1 0 15072 0 1 46116
box -48 -56 240 834
use sg13g2_decap_8  FILLER_60_169
timestamp 1679581782
transform 1 0 17376 0 1 46116
box -48 -56 720 834
use sg13g2_fill_2  FILLER_60_176
timestamp 1677580104
transform 1 0 18048 0 1 46116
box -48 -56 240 834
use sg13g2_fill_1  FILLER_60_178
timestamp 1677579658
transform 1 0 18240 0 1 46116
box -48 -56 144 834
use sg13g2_decap_8  FILLER_61_0
timestamp 1679581782
transform 1 0 1152 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_4  FILLER_61_7
timestamp 1679577901
transform 1 0 1824 0 -1 47628
box -48 -56 432 834
use sg13g2_fill_2  FILLER_61_11
timestamp 1677580104
transform 1 0 2208 0 -1 47628
box -48 -56 240 834
use sg13g2_decap_8  FILLER_61_40
timestamp 1679581782
transform 1 0 4992 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_47
timestamp 1679581782
transform 1 0 5664 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_4  FILLER_61_97
timestamp 1679577901
transform 1 0 10464 0 -1 47628
box -48 -56 432 834
use sg13g2_decap_8  FILLER_61_135
timestamp 1679581782
transform 1 0 14112 0 -1 47628
box -48 -56 720 834
use sg13g2_fill_1  FILLER_61_142
timestamp 1677579658
transform 1 0 14784 0 -1 47628
box -48 -56 144 834
use sg13g2_fill_2  FILLER_61_160
timestamp 1677580104
transform 1 0 16512 0 -1 47628
box -48 -56 240 834
use sg13g2_fill_2  FILLER_61_179
timestamp 1677580104
transform 1 0 18336 0 -1 47628
box -48 -56 240 834
use sg13g2_fill_2  FILLER_61_198
timestamp 1677580104
transform 1 0 20160 0 -1 47628
box -48 -56 240 834
use sg13g2_decap_4  FILLER_62_38
timestamp 1679577901
transform 1 0 4800 0 1 47628
box -48 -56 432 834
use sg13g2_fill_1  FILLER_62_42
timestamp 1677579658
transform 1 0 5184 0 1 47628
box -48 -56 144 834
use sg13g2_decap_8  FILLER_62_70
timestamp 1679581782
transform 1 0 7872 0 1 47628
box -48 -56 720 834
use sg13g2_decap_4  FILLER_62_111
timestamp 1679577901
transform 1 0 11808 0 1 47628
box -48 -56 432 834
use sg13g2_fill_2  FILLER_62_115
timestamp 1677580104
transform 1 0 12192 0 1 47628
box -48 -56 240 834
use sg13g2_fill_2  FILLER_62_138
timestamp 1677580104
transform 1 0 14400 0 1 47628
box -48 -56 240 834
use sg13g2_fill_1  FILLER_62_140
timestamp 1677579658
transform 1 0 14592 0 1 47628
box -48 -56 144 834
use sg13g2_fill_1  FILLER_62_163
timestamp 1677579658
transform 1 0 16800 0 1 47628
box -48 -56 144 834
use sg13g2_fill_2  FILLER_62_198
timestamp 1677580104
transform 1 0 20160 0 1 47628
box -48 -56 240 834
use sg13g2_fill_1  FILLER_63_0
timestamp 1677579658
transform 1 0 1152 0 -1 49140
box -48 -56 144 834
use sg13g2_fill_2  FILLER_63_18
timestamp 1677580104
transform 1 0 2880 0 -1 49140
box -48 -56 240 834
use sg13g2_decap_4  FILLER_63_126
timestamp 1679577901
transform 1 0 13248 0 -1 49140
box -48 -56 432 834
use sg13g2_fill_1  FILLER_63_199
timestamp 1677579658
transform 1 0 20256 0 -1 49140
box -48 -56 144 834
use sg13g2_decap_8  FILLER_64_0
timestamp 1679581782
transform 1 0 1152 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_7
timestamp 1679581782
transform 1 0 1824 0 1 49140
box -48 -56 720 834
use sg13g2_fill_1  FILLER_64_14
timestamp 1677579658
transform 1 0 2496 0 1 49140
box -48 -56 144 834
use sg13g2_decap_4  FILLER_64_41
timestamp 1679577901
transform 1 0 5088 0 1 49140
box -48 -56 432 834
use sg13g2_fill_1  FILLER_64_45
timestamp 1677579658
transform 1 0 5472 0 1 49140
box -48 -56 144 834
use sg13g2_decap_8  FILLER_64_77
timestamp 1679581782
transform 1 0 8544 0 1 49140
box -48 -56 720 834
use sg13g2_fill_2  FILLER_64_84
timestamp 1677580104
transform 1 0 9216 0 1 49140
box -48 -56 240 834
use sg13g2_decap_8  FILLER_64_107
timestamp 1679581782
transform 1 0 11424 0 1 49140
box -48 -56 720 834
use sg13g2_decap_4  FILLER_64_114
timestamp 1679577901
transform 1 0 12096 0 1 49140
box -48 -56 432 834
use sg13g2_fill_2  FILLER_64_118
timestamp 1677580104
transform 1 0 12480 0 1 49140
box -48 -56 240 834
use sg13g2_fill_2  FILLER_64_141
timestamp 1677580104
transform 1 0 14688 0 1 49140
box -48 -56 240 834
use sg13g2_fill_1  FILLER_64_143
timestamp 1677579658
transform 1 0 14880 0 1 49140
box -48 -56 144 834
use sg13g2_fill_1  FILLER_64_163
timestamp 1677579658
transform 1 0 16800 0 1 49140
box -48 -56 144 834
use sg13g2_fill_2  FILLER_64_198
timestamp 1677580104
transform 1 0 20160 0 1 49140
box -48 -56 240 834
use sg13g2_decap_8  FILLER_65_0
timestamp 1679581782
transform 1 0 1152 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_4  FILLER_65_7
timestamp 1679577901
transform 1 0 1824 0 -1 50652
box -48 -56 432 834
use sg13g2_fill_1  FILLER_65_11
timestamp 1677579658
transform 1 0 2208 0 -1 50652
box -48 -56 144 834
use sg13g2_fill_2  FILLER_65_32
timestamp 1677580104
transform 1 0 4224 0 -1 50652
box -48 -56 240 834
use sg13g2_fill_1  FILLER_65_34
timestamp 1677579658
transform 1 0 4416 0 -1 50652
box -48 -56 144 834
use sg13g2_fill_2  FILLER_65_52
timestamp 1677580104
transform 1 0 6144 0 -1 50652
box -48 -56 240 834
use sg13g2_fill_1  FILLER_65_72
timestamp 1677579658
transform 1 0 8064 0 -1 50652
box -48 -56 144 834
use sg13g2_decap_8  FILLER_65_90
timestamp 1679581782
transform 1 0 9792 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_97
timestamp 1679581782
transform 1 0 10464 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_138
timestamp 1679581782
transform 1 0 14400 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_4  FILLER_65_145
timestamp 1679577901
transform 1 0 15072 0 -1 50652
box -48 -56 432 834
use sg13g2_decap_4  FILLER_66_32
timestamp 1679577901
transform 1 0 4224 0 1 50652
box -48 -56 432 834
use sg13g2_decap_8  FILLER_66_91
timestamp 1679581782
transform 1 0 9888 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_98
timestamp 1679581782
transform 1 0 10560 0 1 50652
box -48 -56 720 834
use sg13g2_fill_1  FILLER_66_122
timestamp 1677579658
transform 1 0 12864 0 1 50652
box -48 -56 144 834
use sg13g2_decap_4  FILLER_66_144
timestamp 1679577901
transform 1 0 14976 0 1 50652
box -48 -56 432 834
use sg13g2_fill_1  FILLER_66_148
timestamp 1677579658
transform 1 0 15360 0 1 50652
box -48 -56 144 834
use sg13g2_fill_2  FILLER_66_166
timestamp 1677580104
transform 1 0 17088 0 1 50652
box -48 -56 240 834
use sg13g2_fill_1  FILLER_66_178
timestamp 1677579658
transform 1 0 18240 0 1 50652
box -48 -56 144 834
use sg13g2_fill_2  FILLER_67_0
timestamp 1677580104
transform 1 0 1152 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_2  FILLER_67_40
timestamp 1677580104
transform 1 0 4992 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_67_42
timestamp 1677579658
transform 1 0 5184 0 -1 52164
box -48 -56 144 834
use sg13g2_decap_8  FILLER_67_77
timestamp 1679581782
transform 1 0 8544 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_4  FILLER_67_84
timestamp 1679577901
transform 1 0 9216 0 -1 52164
box -48 -56 432 834
use sg13g2_fill_2  FILLER_67_88
timestamp 1677580104
transform 1 0 9600 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_2  FILLER_67_124
timestamp 1677580104
transform 1 0 13056 0 -1 52164
box -48 -56 240 834
use sg13g2_decap_8  FILLER_67_143
timestamp 1679581782
transform 1 0 14880 0 -1 52164
box -48 -56 720 834
use sg13g2_fill_2  FILLER_67_150
timestamp 1677580104
transform 1 0 15552 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_67_181
timestamp 1677579658
transform 1 0 18528 0 -1 52164
box -48 -56 144 834
use sg13g2_fill_1  FILLER_67_199
timestamp 1677579658
transform 1 0 20256 0 -1 52164
box -48 -56 144 834
use sg13g2_fill_2  FILLER_68_0
timestamp 1677580104
transform 1 0 1152 0 1 52164
box -48 -56 240 834
use sg13g2_fill_2  FILLER_68_29
timestamp 1677580104
transform 1 0 3936 0 1 52164
box -48 -56 240 834
use sg13g2_fill_2  FILLER_68_91
timestamp 1677580104
transform 1 0 9888 0 1 52164
box -48 -56 240 834
use sg13g2_fill_2  FILLER_68_112
timestamp 1677580104
transform 1 0 11904 0 1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_68_114
timestamp 1677579658
transform 1 0 12096 0 1 52164
box -48 -56 144 834
use sg13g2_fill_2  FILLER_68_133
timestamp 1677580104
transform 1 0 13920 0 1 52164
box -48 -56 240 834
use sg13g2_fill_2  FILLER_68_138
timestamp 1677580104
transform 1 0 14400 0 1 52164
box -48 -56 240 834
use sg13g2_fill_2  FILLER_68_157
timestamp 1677580104
transform 1 0 16224 0 1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_68_199
timestamp 1677579658
transform 1 0 20256 0 1 52164
box -48 -56 144 834
use sg13g2_fill_1  FILLER_69_17
timestamp 1677579658
transform 1 0 2784 0 -1 53676
box -48 -56 144 834
use sg13g2_decap_8  FILLER_69_23
timestamp 1679581782
transform 1 0 3360 0 -1 53676
box -48 -56 720 834
use sg13g2_fill_2  FILLER_69_30
timestamp 1677580104
transform 1 0 4032 0 -1 53676
box -48 -56 240 834
use sg13g2_fill_1  FILLER_69_32
timestamp 1677579658
transform 1 0 4224 0 -1 53676
box -48 -56 144 834
use sg13g2_fill_2  FILLER_69_98
timestamp 1677580104
transform 1 0 10560 0 -1 53676
box -48 -56 240 834
use sg13g2_fill_1  FILLER_69_122
timestamp 1677579658
transform 1 0 12864 0 -1 53676
box -48 -56 144 834
use sg13g2_fill_2  FILLER_69_144
timestamp 1677580104
transform 1 0 14976 0 -1 53676
box -48 -56 240 834
use sg13g2_fill_2  FILLER_69_168
timestamp 1677580104
transform 1 0 17280 0 -1 53676
box -48 -56 240 834
use sg13g2_fill_2  FILLER_70_0
timestamp 1677580104
transform 1 0 1152 0 1 53676
box -48 -56 240 834
use sg13g2_fill_1  FILLER_70_62
timestamp 1677579658
transform 1 0 7104 0 1 53676
box -48 -56 144 834
use sg13g2_fill_2  FILLER_70_142
timestamp 1677580104
transform 1 0 14784 0 1 53676
box -48 -56 240 834
use sg13g2_fill_1  FILLER_70_144
timestamp 1677579658
transform 1 0 14976 0 1 53676
box -48 -56 144 834
use sg13g2_fill_2  FILLER_70_175
timestamp 1677580104
transform 1 0 17952 0 1 53676
box -48 -56 240 834
use sg13g2_fill_2  FILLER_70_198
timestamp 1677580104
transform 1 0 20160 0 1 53676
box -48 -56 240 834
use sg13g2_fill_2  FILLER_71_0
timestamp 1677580104
transform 1 0 1152 0 -1 55188
box -48 -56 240 834
use sg13g2_decap_4  FILLER_71_39
timestamp 1679577901
transform 1 0 4896 0 -1 55188
box -48 -56 432 834
use sg13g2_fill_2  FILLER_71_43
timestamp 1677580104
transform 1 0 5280 0 -1 55188
box -48 -56 240 834
use sg13g2_fill_2  FILLER_71_62
timestamp 1677580104
transform 1 0 7104 0 -1 55188
box -48 -56 240 834
use sg13g2_decap_4  FILLER_71_69
timestamp 1679577901
transform 1 0 7776 0 -1 55188
box -48 -56 432 834
use sg13g2_fill_2  FILLER_71_90
timestamp 1677580104
transform 1 0 9792 0 -1 55188
box -48 -56 240 834
use sg13g2_decap_8  FILLER_71_114
timestamp 1679581782
transform 1 0 12096 0 -1 55188
box -48 -56 720 834
use sg13g2_fill_1  FILLER_71_121
timestamp 1677579658
transform 1 0 12768 0 -1 55188
box -48 -56 144 834
use sg13g2_fill_2  FILLER_71_139
timestamp 1677580104
transform 1 0 14496 0 -1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_141
timestamp 1677579658
transform 1 0 14688 0 -1 55188
box -48 -56 144 834
use sg13g2_fill_2  FILLER_71_159
timestamp 1677580104
transform 1 0 16416 0 -1 55188
box -48 -56 240 834
use sg13g2_fill_2  FILLER_71_166
timestamp 1677580104
transform 1 0 17088 0 -1 55188
box -48 -56 240 834
use sg13g2_fill_2  FILLER_71_178
timestamp 1677580104
transform 1 0 18240 0 -1 55188
box -48 -56 240 834
use sg13g2_fill_2  FILLER_71_197
timestamp 1677580104
transform 1 0 20064 0 -1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_199
timestamp 1677579658
transform 1 0 20256 0 -1 55188
box -48 -56 144 834
use sg13g2_fill_1  FILLER_72_0
timestamp 1677579658
transform 1 0 1152 0 1 55188
box -48 -56 144 834
use sg13g2_fill_2  FILLER_72_18
timestamp 1677580104
transform 1 0 2880 0 1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_72_33
timestamp 1677579658
transform 1 0 4320 0 1 55188
box -48 -56 144 834
use sg13g2_decap_8  FILLER_72_115
timestamp 1679581782
transform 1 0 12192 0 1 55188
box -48 -56 720 834
use sg13g2_fill_2  FILLER_72_122
timestamp 1677580104
transform 1 0 12864 0 1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_72_124
timestamp 1677579658
transform 1 0 13056 0 1 55188
box -48 -56 144 834
use sg13g2_decap_8  FILLER_72_142
timestamp 1679581782
transform 1 0 14784 0 1 55188
box -48 -56 720 834
use sg13g2_fill_2  FILLER_72_149
timestamp 1677580104
transform 1 0 15456 0 1 55188
box -48 -56 240 834
use sg13g2_fill_2  FILLER_72_168
timestamp 1677580104
transform 1 0 17280 0 1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_72_170
timestamp 1677579658
transform 1 0 17472 0 1 55188
box -48 -56 144 834
use sg13g2_fill_2  FILLER_72_176
timestamp 1677580104
transform 1 0 18048 0 1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_72_178
timestamp 1677579658
transform 1 0 18240 0 1 55188
box -48 -56 144 834
use sg13g2_decap_4  FILLER_72_196
timestamp 1679577901
transform 1 0 19968 0 1 55188
box -48 -56 432 834
use sg13g2_decap_4  FILLER_73_0
timestamp 1679577901
transform 1 0 1152 0 -1 56700
box -48 -56 432 834
use sg13g2_fill_2  FILLER_73_21
timestamp 1677580104
transform 1 0 3168 0 -1 56700
box -48 -56 240 834
use sg13g2_decap_4  FILLER_73_43
timestamp 1679577901
transform 1 0 5280 0 -1 56700
box -48 -56 432 834
use sg13g2_fill_1  FILLER_73_47
timestamp 1677579658
transform 1 0 5664 0 -1 56700
box -48 -56 144 834
use sg13g2_decap_4  FILLER_73_84
timestamp 1679577901
transform 1 0 9216 0 -1 56700
box -48 -56 432 834
use sg13g2_decap_8  FILLER_73_105
timestamp 1679581782
transform 1 0 11232 0 -1 56700
box -48 -56 720 834
use sg13g2_fill_1  FILLER_73_129
timestamp 1677579658
transform 1 0 13536 0 -1 56700
box -48 -56 144 834
use sg13g2_decap_8  FILLER_73_151
timestamp 1679581782
transform 1 0 15648 0 -1 56700
box -48 -56 720 834
use sg13g2_fill_1  FILLER_73_158
timestamp 1677579658
transform 1 0 16320 0 -1 56700
box -48 -56 144 834
use sg13g2_fill_1  FILLER_73_199
timestamp 1677579658
transform 1 0 20256 0 -1 56700
box -48 -56 144 834
use sg13g2_fill_1  FILLER_74_0
timestamp 1677579658
transform 1 0 1152 0 1 56700
box -48 -56 144 834
use sg13g2_decap_8  FILLER_74_44
timestamp 1679581782
transform 1 0 5376 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_51
timestamp 1679581782
transform 1 0 6048 0 1 56700
box -48 -56 720 834
use sg13g2_fill_2  FILLER_74_58
timestamp 1677580104
transform 1 0 6720 0 1 56700
box -48 -56 240 834
use sg13g2_decap_4  FILLER_74_107
timestamp 1679577901
transform 1 0 11424 0 1 56700
box -48 -56 432 834
use sg13g2_fill_1  FILLER_74_111
timestamp 1677579658
transform 1 0 11808 0 1 56700
box -48 -56 144 834
use sg13g2_decap_8  FILLER_74_150
timestamp 1679581782
transform 1 0 15552 0 1 56700
box -48 -56 720 834
use sg13g2_fill_1  FILLER_75_0
timestamp 1677579658
transform 1 0 1152 0 -1 58212
box -48 -56 144 834
use sg13g2_fill_2  FILLER_75_18
timestamp 1677580104
transform 1 0 2880 0 -1 58212
box -48 -56 240 834
use sg13g2_decap_8  FILLER_75_33
timestamp 1679581782
transform 1 0 4320 0 -1 58212
box -48 -56 720 834
use sg13g2_fill_2  FILLER_75_40
timestamp 1677580104
transform 1 0 4992 0 -1 58212
box -48 -56 240 834
use sg13g2_fill_1  FILLER_75_42
timestamp 1677579658
transform 1 0 5184 0 -1 58212
box -48 -56 144 834
use sg13g2_decap_4  FILLER_75_60
timestamp 1679577901
transform 1 0 6912 0 -1 58212
box -48 -56 432 834
use sg13g2_fill_2  FILLER_75_64
timestamp 1677580104
transform 1 0 7296 0 -1 58212
box -48 -56 240 834
use sg13g2_decap_4  FILLER_75_83
timestamp 1679577901
transform 1 0 9120 0 -1 58212
box -48 -56 432 834
use sg13g2_fill_2  FILLER_75_87
timestamp 1677580104
transform 1 0 9504 0 -1 58212
box -48 -56 240 834
use sg13g2_decap_4  FILLER_75_106
timestamp 1679577901
transform 1 0 11328 0 -1 58212
box -48 -56 432 834
use sg13g2_fill_1  FILLER_75_110
timestamp 1677579658
transform 1 0 11712 0 -1 58212
box -48 -56 144 834
use sg13g2_decap_4  FILLER_75_128
timestamp 1679577901
transform 1 0 13440 0 -1 58212
box -48 -56 432 834
use sg13g2_fill_1  FILLER_75_132
timestamp 1677579658
transform 1 0 13824 0 -1 58212
box -48 -56 144 834
use sg13g2_fill_2  FILLER_75_198
timestamp 1677580104
transform 1 0 20160 0 -1 58212
box -48 -56 240 834
use sg13g2_fill_2  FILLER_76_0
timestamp 1677580104
transform 1 0 1152 0 1 58212
box -48 -56 240 834
use sg13g2_fill_2  FILLER_76_22
timestamp 1677580104
transform 1 0 3264 0 1 58212
box -48 -56 240 834
use sg13g2_fill_2  FILLER_76_62
timestamp 1677580104
transform 1 0 7104 0 1 58212
box -48 -56 240 834
use sg13g2_fill_1  FILLER_76_64
timestamp 1677579658
transform 1 0 7296 0 1 58212
box -48 -56 144 834
use sg13g2_decap_4  FILLER_76_86
timestamp 1679577901
transform 1 0 9408 0 1 58212
box -48 -56 432 834
use sg13g2_fill_1  FILLER_76_90
timestamp 1677579658
transform 1 0 9792 0 1 58212
box -48 -56 144 834
use sg13g2_fill_1  FILLER_76_129
timestamp 1677579658
transform 1 0 13536 0 1 58212
box -48 -56 144 834
use sg13g2_fill_2  FILLER_76_169
timestamp 1677580104
transform 1 0 17376 0 1 58212
box -48 -56 240 834
use sg13g2_fill_1  FILLER_76_188
timestamp 1677579658
transform 1 0 19200 0 1 58212
box -48 -56 144 834
use sg13g2_fill_2  FILLER_76_197
timestamp 1677580104
transform 1 0 20064 0 1 58212
box -48 -56 240 834
use sg13g2_fill_1  FILLER_76_199
timestamp 1677579658
transform 1 0 20256 0 1 58212
box -48 -56 144 834
use sg13g2_decap_8  FILLER_77_0
timestamp 1679581782
transform 1 0 1152 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_7
timestamp 1679581782
transform 1 0 1824 0 -1 59724
box -48 -56 720 834
use sg13g2_fill_2  FILLER_77_14
timestamp 1677580104
transform 1 0 2496 0 -1 59724
box -48 -56 240 834
use sg13g2_decap_8  FILLER_77_40
timestamp 1679581782
transform 1 0 4992 0 -1 59724
box -48 -56 720 834
use sg13g2_fill_2  FILLER_77_47
timestamp 1677580104
transform 1 0 5664 0 -1 59724
box -48 -56 240 834
use sg13g2_fill_1  FILLER_77_49
timestamp 1677579658
transform 1 0 5856 0 -1 59724
box -48 -56 144 834
use sg13g2_fill_2  FILLER_77_67
timestamp 1677580104
transform 1 0 7584 0 -1 59724
box -48 -56 240 834
use sg13g2_decap_8  FILLER_77_107
timestamp 1679581782
transform 1 0 11424 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_114
timestamp 1679581782
transform 1 0 12096 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_121
timestamp 1679581782
transform 1 0 12768 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_4  FILLER_77_128
timestamp 1679577901
transform 1 0 13440 0 -1 59724
box -48 -56 432 834
use sg13g2_fill_1  FILLER_77_132
timestamp 1677579658
transform 1 0 13824 0 -1 59724
box -48 -56 144 834
use sg13g2_fill_2  FILLER_77_158
timestamp 1677580104
transform 1 0 16320 0 -1 59724
box -48 -56 240 834
use sg13g2_fill_1  FILLER_77_160
timestamp 1677579658
transform 1 0 16512 0 -1 59724
box -48 -56 144 834
use sg13g2_fill_2  FILLER_77_197
timestamp 1677580104
transform 1 0 20064 0 -1 59724
box -48 -56 240 834
use sg13g2_fill_1  FILLER_77_199
timestamp 1677579658
transform 1 0 20256 0 -1 59724
box -48 -56 144 834
use sg13g2_fill_2  FILLER_78_17
timestamp 1677580104
transform 1 0 2784 0 1 59724
box -48 -56 240 834
use sg13g2_decap_8  FILLER_78_36
timestamp 1679581782
transform 1 0 4608 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_43
timestamp 1679581782
transform 1 0 5280 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_71
timestamp 1679581782
transform 1 0 7968 0 1 59724
box -48 -56 720 834
use sg13g2_decap_4  FILLER_78_78
timestamp 1679577901
transform 1 0 8640 0 1 59724
box -48 -56 432 834
use sg13g2_fill_1  FILLER_78_82
timestamp 1677579658
transform 1 0 9024 0 1 59724
box -48 -56 144 834
use sg13g2_decap_8  FILLER_78_100
timestamp 1679581782
transform 1 0 10752 0 1 59724
box -48 -56 720 834
use sg13g2_decap_4  FILLER_78_150
timestamp 1679577901
transform 1 0 15552 0 1 59724
box -48 -56 432 834
use sg13g2_decap_4  FILLER_78_171
timestamp 1679577901
transform 1 0 17568 0 1 59724
box -48 -56 432 834
use sg13g2_fill_1  FILLER_78_175
timestamp 1677579658
transform 1 0 17952 0 1 59724
box -48 -56 144 834
use sg13g2_fill_2  FILLER_78_197
timestamp 1677580104
transform 1 0 20064 0 1 59724
box -48 -56 240 834
use sg13g2_fill_1  FILLER_78_199
timestamp 1677579658
transform 1 0 20256 0 1 59724
box -48 -56 144 834
use sg13g2_fill_2  FILLER_79_0
timestamp 1677580104
transform 1 0 1152 0 -1 61236
box -48 -56 240 834
use sg13g2_decap_4  FILLER_79_40
timestamp 1679577901
transform 1 0 4992 0 -1 61236
box -48 -56 432 834
use sg13g2_fill_2  FILLER_79_95
timestamp 1677580104
transform 1 0 10272 0 -1 61236
box -48 -56 240 834
use sg13g2_fill_1  FILLER_79_97
timestamp 1677579658
transform 1 0 10464 0 -1 61236
box -48 -56 144 834
use sg13g2_decap_8  FILLER_79_119
timestamp 1679581782
transform 1 0 12576 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_143
timestamp 1679581782
transform 1 0 14880 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_4  FILLER_79_150
timestamp 1679577901
transform 1 0 15552 0 -1 61236
box -48 -56 432 834
use sg13g2_decap_8  FILLER_80_0
timestamp 1679581782
transform 1 0 1152 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_7
timestamp 1679581782
transform 1 0 1824 0 1 61236
box -48 -56 720 834
use sg13g2_fill_2  FILLER_80_14
timestamp 1677580104
transform 1 0 2496 0 1 61236
box -48 -56 240 834
use sg13g2_decap_4  FILLER_80_37
timestamp 1679577901
transform 1 0 4704 0 1 61236
box -48 -56 432 834
use sg13g2_fill_2  FILLER_80_41
timestamp 1677580104
transform 1 0 5088 0 1 61236
box -48 -56 240 834
use sg13g2_fill_2  FILLER_80_60
timestamp 1677580104
transform 1 0 6912 0 1 61236
box -48 -56 240 834
use sg13g2_decap_4  FILLER_80_134
timestamp 1679577901
transform 1 0 14016 0 1 61236
box -48 -56 432 834
use sg13g2_fill_1  FILLER_80_138
timestamp 1677579658
transform 1 0 14400 0 1 61236
box -48 -56 144 834
use sg13g2_decap_8  FILLER_80_173
timestamp 1679581782
transform 1 0 17760 0 1 61236
box -48 -56 720 834
use sg13g2_fill_1  FILLER_80_180
timestamp 1677579658
transform 1 0 18432 0 1 61236
box -48 -56 144 834
use sg13g2_fill_2  FILLER_80_197
timestamp 1677580104
transform 1 0 20064 0 1 61236
box -48 -56 240 834
use sg13g2_fill_1  FILLER_80_199
timestamp 1677579658
transform 1 0 20256 0 1 61236
box -48 -56 144 834
use sg13g2_fill_1  FILLER_81_17
timestamp 1677579658
transform 1 0 2784 0 -1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_81_52
timestamp 1679581782
transform 1 0 6144 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_4  FILLER_81_59
timestamp 1679577901
transform 1 0 6816 0 -1 62748
box -48 -56 432 834
use sg13g2_fill_2  FILLER_81_63
timestamp 1677580104
transform 1 0 7200 0 -1 62748
box -48 -56 240 834
use sg13g2_decap_8  FILLER_81_86
timestamp 1679581782
transform 1 0 9408 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_93
timestamp 1679581782
transform 1 0 10080 0 -1 62748
box -48 -56 720 834
use sg13g2_fill_1  FILLER_81_100
timestamp 1677579658
transform 1 0 10752 0 -1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_81_118
timestamp 1679581782
transform 1 0 12480 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_4  FILLER_81_125
timestamp 1679577901
transform 1 0 13152 0 -1 62748
box -48 -56 432 834
use sg13g2_fill_2  FILLER_81_129
timestamp 1677580104
transform 1 0 13536 0 -1 62748
box -48 -56 240 834
use sg13g2_decap_8  FILLER_81_152
timestamp 1679581782
transform 1 0 15744 0 -1 62748
box -48 -56 720 834
use sg13g2_fill_1  FILLER_81_159
timestamp 1677579658
transform 1 0 16416 0 -1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_81_164
timestamp 1679581782
transform 1 0 16896 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_4  FILLER_81_171
timestamp 1679577901
transform 1 0 17568 0 -1 62748
box -48 -56 432 834
use sg13g2_decap_8  FILLER_82_0
timestamp 1679581782
transform 1 0 1152 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_7
timestamp 1679581782
transform 1 0 1824 0 1 62748
box -48 -56 720 834
use sg13g2_fill_2  FILLER_82_14
timestamp 1677580104
transform 1 0 2496 0 1 62748
box -48 -56 240 834
use sg13g2_decap_8  FILLER_82_37
timestamp 1679581782
transform 1 0 4704 0 1 62748
box -48 -56 720 834
use sg13g2_fill_2  FILLER_82_44
timestamp 1677580104
transform 1 0 5376 0 1 62748
box -48 -56 240 834
use sg13g2_fill_1  FILLER_82_63
timestamp 1677579658
transform 1 0 7200 0 1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_82_115
timestamp 1679581782
transform 1 0 12192 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_122
timestamp 1679581782
transform 1 0 12864 0 1 62748
box -48 -56 720 834
use sg13g2_fill_2  FILLER_82_129
timestamp 1677580104
transform 1 0 13536 0 1 62748
box -48 -56 240 834
use sg13g2_fill_1  FILLER_82_148
timestamp 1677579658
transform 1 0 15360 0 1 62748
box -48 -56 144 834
use sg13g2_decap_4  FILLER_82_194
timestamp 1679577901
transform 1 0 19776 0 1 62748
box -48 -56 432 834
use sg13g2_fill_2  FILLER_82_198
timestamp 1677580104
transform 1 0 20160 0 1 62748
box -48 -56 240 834
use sg13g2_decap_4  FILLER_83_0
timestamp 1679577901
transform 1 0 1152 0 -1 64260
box -48 -56 432 834
use sg13g2_fill_1  FILLER_83_4
timestamp 1677579658
transform 1 0 1536 0 -1 64260
box -48 -56 144 834
use sg13g2_decap_8  FILLER_83_43
timestamp 1679581782
transform 1 0 5280 0 -1 64260
box -48 -56 720 834
use sg13g2_fill_2  FILLER_83_50
timestamp 1677580104
transform 1 0 5952 0 -1 64260
box -48 -56 240 834
use sg13g2_fill_1  FILLER_83_52
timestamp 1677579658
transform 1 0 6144 0 -1 64260
box -48 -56 144 834
use sg13g2_decap_8  FILLER_83_74
timestamp 1679581782
transform 1 0 8256 0 -1 64260
box -48 -56 720 834
use sg13g2_fill_1  FILLER_83_81
timestamp 1677579658
transform 1 0 8928 0 -1 64260
box -48 -56 144 834
use sg13g2_decap_8  FILLER_83_120
timestamp 1679581782
transform 1 0 12672 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_4  FILLER_83_127
timestamp 1679577901
transform 1 0 13344 0 -1 64260
box -48 -56 432 834
use sg13g2_decap_8  FILLER_83_152
timestamp 1679581782
transform 1 0 15744 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_159
timestamp 1679581782
transform 1 0 16416 0 -1 64260
box -48 -56 720 834
use sg13g2_fill_2  FILLER_83_166
timestamp 1677580104
transform 1 0 17088 0 -1 64260
box -48 -56 240 834
use sg13g2_fill_2  FILLER_83_197
timestamp 1677580104
transform 1 0 20064 0 -1 64260
box -48 -56 240 834
use sg13g2_fill_1  FILLER_83_199
timestamp 1677579658
transform 1 0 20256 0 -1 64260
box -48 -56 144 834
use sg13g2_decap_8  FILLER_84_0
timestamp 1679581782
transform 1 0 1152 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_7
timestamp 1679581782
transform 1 0 1824 0 1 64260
box -48 -56 720 834
use sg13g2_fill_2  FILLER_84_86
timestamp 1677580104
transform 1 0 9408 0 1 64260
box -48 -56 240 834
use sg13g2_decap_8  FILLER_84_109
timestamp 1679581782
transform 1 0 11616 0 1 64260
box -48 -56 720 834
use sg13g2_fill_1  FILLER_84_150
timestamp 1677579658
transform 1 0 15552 0 1 64260
box -48 -56 144 834
use sg13g2_decap_4  FILLER_84_168
timestamp 1679577901
transform 1 0 17280 0 1 64260
box -48 -56 432 834
use sg13g2_fill_2  FILLER_84_197
timestamp 1677580104
transform 1 0 20064 0 1 64260
box -48 -56 240 834
use sg13g2_fill_1  FILLER_84_199
timestamp 1677579658
transform 1 0 20256 0 1 64260
box -48 -56 144 834
use sg13g2_decap_8  FILLER_85_0
timestamp 1679581782
transform 1 0 1152 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_7
timestamp 1679581782
transform 1 0 1824 0 -1 65772
box -48 -56 720 834
use sg13g2_fill_1  FILLER_85_14
timestamp 1677579658
transform 1 0 2496 0 -1 65772
box -48 -56 144 834
use sg13g2_decap_8  FILLER_85_36
timestamp 1679581782
transform 1 0 4608 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_4  FILLER_85_43
timestamp 1679577901
transform 1 0 5280 0 -1 65772
box -48 -56 432 834
use sg13g2_fill_1  FILLER_85_47
timestamp 1677579658
transform 1 0 5664 0 -1 65772
box -48 -56 144 834
use sg13g2_decap_8  FILLER_85_120
timestamp 1679581782
transform 1 0 12672 0 -1 65772
box -48 -56 720 834
use sg13g2_fill_2  FILLER_85_127
timestamp 1677580104
transform 1 0 13344 0 -1 65772
box -48 -56 240 834
use sg13g2_decap_4  FILLER_85_150
timestamp 1679577901
transform 1 0 15552 0 -1 65772
box -48 -56 432 834
use sg13g2_fill_2  FILLER_85_154
timestamp 1677580104
transform 1 0 15936 0 -1 65772
box -48 -56 240 834
use sg13g2_decap_4  FILLER_85_180
timestamp 1679577901
transform 1 0 18432 0 -1 65772
box -48 -56 432 834
use sg13g2_fill_1  FILLER_85_184
timestamp 1677579658
transform 1 0 18816 0 -1 65772
box -48 -56 144 834
use sg13g2_fill_2  FILLER_85_197
timestamp 1677580104
transform 1 0 20064 0 -1 65772
box -48 -56 240 834
use sg13g2_fill_1  FILLER_85_199
timestamp 1677579658
transform 1 0 20256 0 -1 65772
box -48 -56 144 834
use sg13g2_fill_2  FILLER_86_0
timestamp 1677580104
transform 1 0 1152 0 1 65772
box -48 -56 240 834
use sg13g2_decap_4  FILLER_86_19
timestamp 1679577901
transform 1 0 2976 0 1 65772
box -48 -56 432 834
use sg13g2_fill_1  FILLER_86_23
timestamp 1677579658
transform 1 0 3360 0 1 65772
box -48 -56 144 834
use sg13g2_fill_2  FILLER_86_45
timestamp 1677580104
transform 1 0 5472 0 1 65772
box -48 -56 240 834
use sg13g2_decap_8  FILLER_86_68
timestamp 1679581782
transform 1 0 7680 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_75
timestamp 1679581782
transform 1 0 8352 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_150
timestamp 1679581782
transform 1 0 15552 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_157
timestamp 1679581782
transform 1 0 16224 0 1 65772
box -48 -56 720 834
use sg13g2_fill_1  FILLER_86_164
timestamp 1677579658
transform 1 0 16896 0 1 65772
box -48 -56 144 834
use sg13g2_fill_2  FILLER_86_197
timestamp 1677580104
transform 1 0 20064 0 1 65772
box -48 -56 240 834
use sg13g2_fill_1  FILLER_86_199
timestamp 1677579658
transform 1 0 20256 0 1 65772
box -48 -56 144 834
use sg13g2_decap_4  FILLER_87_17
timestamp 1679577901
transform 1 0 2784 0 -1 67284
box -48 -56 432 834
use sg13g2_fill_1  FILLER_87_21
timestamp 1677579658
transform 1 0 3168 0 -1 67284
box -48 -56 144 834
use sg13g2_decap_8  FILLER_87_56
timestamp 1679581782
transform 1 0 6528 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_4  FILLER_87_63
timestamp 1679577901
transform 1 0 7200 0 -1 67284
box -48 -56 432 834
use sg13g2_fill_2  FILLER_87_67
timestamp 1677580104
transform 1 0 7584 0 -1 67284
box -48 -56 240 834
use sg13g2_fill_2  FILLER_87_90
timestamp 1677580104
transform 1 0 9792 0 -1 67284
box -48 -56 240 834
use sg13g2_fill_1  FILLER_87_109
timestamp 1677579658
transform 1 0 11616 0 -1 67284
box -48 -56 144 834
use sg13g2_fill_2  FILLER_87_148
timestamp 1677580104
transform 1 0 15360 0 -1 67284
box -48 -56 240 834
use sg13g2_decap_8  FILLER_87_184
timestamp 1679581782
transform 1 0 18816 0 -1 67284
box -48 -56 720 834
use sg13g2_fill_1  FILLER_87_191
timestamp 1677579658
transform 1 0 19488 0 -1 67284
box -48 -56 144 834
use sg13g2_fill_1  FILLER_88_0
timestamp 1677579658
transform 1 0 1152 0 1 67284
box -48 -56 144 834
use sg13g2_fill_1  FILLER_88_86
timestamp 1677579658
transform 1 0 9408 0 1 67284
box -48 -56 144 834
use sg13g2_fill_2  FILLER_88_125
timestamp 1677580104
transform 1 0 13152 0 1 67284
box -48 -56 240 834
use sg13g2_decap_8  FILLER_88_144
timestamp 1679581782
transform 1 0 14976 0 1 67284
box -48 -56 720 834
use sg13g2_fill_2  FILLER_88_197
timestamp 1677580104
transform 1 0 20064 0 1 67284
box -48 -56 240 834
use sg13g2_fill_1  FILLER_88_199
timestamp 1677579658
transform 1 0 20256 0 1 67284
box -48 -56 144 834
use sg13g2_fill_2  FILLER_89_0
timestamp 1677580104
transform 1 0 1152 0 -1 68796
box -48 -56 240 834
use sg13g2_fill_1  FILLER_89_2
timestamp 1677579658
transform 1 0 1344 0 -1 68796
box -48 -56 144 834
use sg13g2_fill_2  FILLER_89_20
timestamp 1677580104
transform 1 0 3072 0 -1 68796
box -48 -56 240 834
use sg13g2_decap_8  FILLER_89_43
timestamp 1679581782
transform 1 0 5280 0 -1 68796
box -48 -56 720 834
use sg13g2_fill_2  FILLER_89_50
timestamp 1677580104
transform 1 0 5952 0 -1 68796
box -48 -56 240 834
use sg13g2_decap_8  FILLER_89_90
timestamp 1679581782
transform 1 0 9792 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_118
timestamp 1679581782
transform 1 0 12480 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_125
timestamp 1679581782
transform 1 0 13152 0 -1 68796
box -48 -56 720 834
use sg13g2_fill_2  FILLER_89_132
timestamp 1677580104
transform 1 0 13824 0 -1 68796
box -48 -56 240 834
use sg13g2_fill_2  FILLER_89_168
timestamp 1677580104
transform 1 0 17280 0 -1 68796
box -48 -56 240 834
use sg13g2_fill_1  FILLER_89_199
timestamp 1677579658
transform 1 0 20256 0 -1 68796
box -48 -56 144 834
use sg13g2_decap_8  FILLER_90_0
timestamp 1679581782
transform 1 0 1152 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_7
timestamp 1679581782
transform 1 0 1824 0 1 68796
box -48 -56 720 834
use sg13g2_fill_2  FILLER_90_14
timestamp 1677580104
transform 1 0 2496 0 1 68796
box -48 -56 240 834
use sg13g2_fill_2  FILLER_90_54
timestamp 1677580104
transform 1 0 6336 0 1 68796
box -48 -56 240 834
use sg13g2_fill_1  FILLER_90_56
timestamp 1677579658
transform 1 0 6528 0 1 68796
box -48 -56 144 834
use sg13g2_fill_2  FILLER_90_78
timestamp 1677580104
transform 1 0 8640 0 1 68796
box -48 -56 240 834
use sg13g2_fill_1  FILLER_90_97
timestamp 1677579658
transform 1 0 10464 0 1 68796
box -48 -56 144 834
use sg13g2_decap_4  FILLER_90_149
timestamp 1679577901
transform 1 0 15456 0 1 68796
box -48 -56 432 834
use sg13g2_fill_2  FILLER_90_153
timestamp 1677580104
transform 1 0 15840 0 1 68796
box -48 -56 240 834
use sg13g2_fill_2  FILLER_90_197
timestamp 1677580104
transform 1 0 20064 0 1 68796
box -48 -56 240 834
use sg13g2_fill_1  FILLER_90_199
timestamp 1677579658
transform 1 0 20256 0 1 68796
box -48 -56 144 834
use sg13g2_fill_1  FILLER_91_17
timestamp 1677579658
transform 1 0 2784 0 -1 70308
box -48 -56 144 834
use sg13g2_decap_4  FILLER_91_69
timestamp 1679577901
transform 1 0 7776 0 -1 70308
box -48 -56 432 834
use sg13g2_fill_2  FILLER_91_73
timestamp 1677580104
transform 1 0 8160 0 -1 70308
box -48 -56 240 834
use sg13g2_decap_8  FILLER_91_113
timestamp 1679581782
transform 1 0 12000 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_120
timestamp 1679581782
transform 1 0 12672 0 -1 70308
box -48 -56 720 834
use sg13g2_fill_1  FILLER_91_127
timestamp 1677579658
transform 1 0 13344 0 -1 70308
box -48 -56 144 834
use sg13g2_decap_4  FILLER_91_145
timestamp 1679577901
transform 1 0 15072 0 -1 70308
box -48 -56 432 834
use sg13g2_fill_1  FILLER_91_199
timestamp 1677579658
transform 1 0 20256 0 -1 70308
box -48 -56 144 834
use sg13g2_decap_8  FILLER_92_0
timestamp 1679581782
transform 1 0 1152 0 1 70308
box -48 -56 720 834
use sg13g2_decap_4  FILLER_92_7
timestamp 1679577901
transform 1 0 1824 0 1 70308
box -48 -56 432 834
use sg13g2_fill_1  FILLER_92_11
timestamp 1677579658
transform 1 0 2208 0 1 70308
box -48 -56 144 834
use sg13g2_decap_8  FILLER_92_83
timestamp 1679581782
transform 1 0 9120 0 1 70308
box -48 -56 720 834
use sg13g2_decap_4  FILLER_92_90
timestamp 1679577901
transform 1 0 9792 0 1 70308
box -48 -56 432 834
use sg13g2_fill_1  FILLER_92_94
timestamp 1677579658
transform 1 0 10176 0 1 70308
box -48 -56 144 834
use sg13g2_fill_2  FILLER_92_129
timestamp 1677580104
transform 1 0 13536 0 1 70308
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_131
timestamp 1677579658
transform 1 0 13728 0 1 70308
box -48 -56 144 834
use sg13g2_decap_4  FILLER_92_149
timestamp 1679577901
transform 1 0 15456 0 1 70308
box -48 -56 432 834
use sg13g2_fill_2  FILLER_92_153
timestamp 1677580104
transform 1 0 15840 0 1 70308
box -48 -56 240 834
use sg13g2_fill_2  FILLER_92_197
timestamp 1677580104
transform 1 0 20064 0 1 70308
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_199
timestamp 1677579658
transform 1 0 20256 0 1 70308
box -48 -56 144 834
use sg13g2_fill_2  FILLER_93_0
timestamp 1677580104
transform 1 0 1152 0 -1 71820
box -48 -56 240 834
use sg13g2_fill_1  FILLER_93_2
timestamp 1677579658
transform 1 0 1344 0 -1 71820
box -48 -56 144 834
use sg13g2_decap_8  FILLER_93_20
timestamp 1679581782
transform 1 0 3072 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_27
timestamp 1679581782
transform 1 0 3744 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_101
timestamp 1679581782
transform 1 0 10848 0 -1 71820
box -48 -56 720 834
use sg13g2_fill_2  FILLER_93_108
timestamp 1677580104
transform 1 0 11520 0 -1 71820
box -48 -56 240 834
use sg13g2_fill_1  FILLER_93_110
timestamp 1677579658
transform 1 0 11712 0 -1 71820
box -48 -56 144 834
use sg13g2_fill_2  FILLER_93_170
timestamp 1677580104
transform 1 0 17472 0 -1 71820
box -48 -56 240 834
use sg13g2_fill_2  FILLER_93_193
timestamp 1677580104
transform 1 0 19680 0 -1 71820
box -48 -56 240 834
use sg13g2_fill_1  FILLER_93_199
timestamp 1677579658
transform 1 0 20256 0 -1 71820
box -48 -56 144 834
use sg13g2_decap_8  FILLER_94_17
timestamp 1679581782
transform 1 0 2784 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_24
timestamp 1679581782
transform 1 0 3456 0 1 71820
box -48 -56 720 834
use sg13g2_fill_1  FILLER_94_31
timestamp 1677579658
transform 1 0 4128 0 1 71820
box -48 -56 144 834
use sg13g2_decap_8  FILLER_94_83
timestamp 1679581782
transform 1 0 9120 0 1 71820
box -48 -56 720 834
use sg13g2_decap_4  FILLER_94_90
timestamp 1679577901
transform 1 0 9792 0 1 71820
box -48 -56 432 834
use sg13g2_fill_1  FILLER_94_94
timestamp 1677579658
transform 1 0 10176 0 1 71820
box -48 -56 144 834
use sg13g2_fill_2  FILLER_94_129
timestamp 1677580104
transform 1 0 13536 0 1 71820
box -48 -56 240 834
use sg13g2_fill_1  FILLER_94_131
timestamp 1677579658
transform 1 0 13728 0 1 71820
box -48 -56 144 834
use sg13g2_decap_8  FILLER_94_149
timestamp 1679581782
transform 1 0 15456 0 1 71820
box -48 -56 720 834
use sg13g2_decap_4  FILLER_94_156
timestamp 1679577901
transform 1 0 16128 0 1 71820
box -48 -56 432 834
use sg13g2_fill_1  FILLER_94_160
timestamp 1677579658
transform 1 0 16512 0 1 71820
box -48 -56 144 834
use sg13g2_fill_2  FILLER_94_182
timestamp 1677580104
transform 1 0 18624 0 1 71820
box -48 -56 240 834
use sg13g2_fill_1  FILLER_94_184
timestamp 1677579658
transform 1 0 18816 0 1 71820
box -48 -56 144 834
use sg13g2_fill_2  FILLER_94_197
timestamp 1677580104
transform 1 0 20064 0 1 71820
box -48 -56 240 834
use sg13g2_fill_1  FILLER_94_199
timestamp 1677579658
transform 1 0 20256 0 1 71820
box -48 -56 144 834
use sg13g2_decap_8  FILLER_95_0
timestamp 1679581782
transform 1 0 1152 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_7
timestamp 1679581782
transform 1 0 1824 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_14
timestamp 1679581782
transform 1 0 2496 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_21
timestamp 1679581782
transform 1 0 3168 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_45
timestamp 1679581782
transform 1 0 5472 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_52
timestamp 1679581782
transform 1 0 6144 0 -1 73332
box -48 -56 720 834
use sg13g2_fill_2  FILLER_95_59
timestamp 1677580104
transform 1 0 6816 0 -1 73332
box -48 -56 240 834
use sg13g2_decap_8  FILLER_95_133
timestamp 1679581782
transform 1 0 13920 0 -1 73332
box -48 -56 720 834
use sg13g2_fill_2  FILLER_95_140
timestamp 1677580104
transform 1 0 14592 0 -1 73332
box -48 -56 240 834
use sg13g2_fill_1  FILLER_95_142
timestamp 1677579658
transform 1 0 14784 0 -1 73332
box -48 -56 144 834
use sg13g2_fill_2  FILLER_95_197
timestamp 1677580104
transform 1 0 20064 0 -1 73332
box -48 -56 240 834
use sg13g2_fill_1  FILLER_95_199
timestamp 1677579658
transform 1 0 20256 0 -1 73332
box -48 -56 144 834
use sg13g2_decap_8  FILLER_96_0
timestamp 1679581782
transform 1 0 1152 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_7
timestamp 1679581782
transform 1 0 1824 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_14
timestamp 1679581782
transform 1 0 2496 0 1 73332
box -48 -56 720 834
use sg13g2_decap_4  FILLER_96_21
timestamp 1679577901
transform 1 0 3168 0 1 73332
box -48 -56 432 834
use sg13g2_fill_1  FILLER_96_25
timestamp 1677579658
transform 1 0 3552 0 1 73332
box -48 -56 144 834
use sg13g2_decap_8  FILLER_96_64
timestamp 1679581782
transform 1 0 7296 0 1 73332
box -48 -56 720 834
use sg13g2_decap_4  FILLER_96_71
timestamp 1679577901
transform 1 0 7968 0 1 73332
box -48 -56 432 834
use sg13g2_decap_8  FILLER_96_96
timestamp 1679581782
transform 1 0 10368 0 1 73332
box -48 -56 720 834
use sg13g2_fill_2  FILLER_96_103
timestamp 1677580104
transform 1 0 11040 0 1 73332
box -48 -56 240 834
use sg13g2_fill_1  FILLER_96_126
timestamp 1677579658
transform 1 0 13248 0 1 73332
box -48 -56 144 834
use sg13g2_decap_4  FILLER_96_161
timestamp 1679577901
transform 1 0 16608 0 1 73332
box -48 -56 432 834
use sg13g2_fill_1  FILLER_96_165
timestamp 1677579658
transform 1 0 16992 0 1 73332
box -48 -56 144 834
use sg13g2_fill_2  FILLER_96_183
timestamp 1677580104
transform 1 0 18720 0 1 73332
box -48 -56 240 834
use sg13g2_fill_2  FILLER_96_197
timestamp 1677580104
transform 1 0 20064 0 1 73332
box -48 -56 240 834
use sg13g2_fill_1  FILLER_96_199
timestamp 1677579658
transform 1 0 20256 0 1 73332
box -48 -56 144 834
use sg13g2_decap_8  FILLER_97_0
timestamp 1679581782
transform 1 0 1152 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_7
timestamp 1679581782
transform 1 0 1824 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_14
timestamp 1679581782
transform 1 0 2496 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_21
timestamp 1679581782
transform 1 0 3168 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_28
timestamp 1679581782
transform 1 0 3840 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_4  FILLER_97_35
timestamp 1679577901
transform 1 0 4512 0 -1 74844
box -48 -56 432 834
use sg13g2_fill_2  FILLER_97_39
timestamp 1677580104
transform 1 0 4896 0 -1 74844
box -48 -56 240 834
use sg13g2_decap_4  FILLER_97_96
timestamp 1679577901
transform 1 0 10368 0 -1 74844
box -48 -56 432 834
use sg13g2_fill_1  FILLER_97_100
timestamp 1677579658
transform 1 0 10752 0 -1 74844
box -48 -56 144 834
use sg13g2_decap_4  FILLER_97_139
timestamp 1679577901
transform 1 0 14496 0 -1 74844
box -48 -56 432 834
use sg13g2_fill_2  FILLER_97_143
timestamp 1677580104
transform 1 0 14880 0 -1 74844
box -48 -56 240 834
use sg13g2_fill_2  FILLER_97_166
timestamp 1677580104
transform 1 0 17088 0 -1 74844
box -48 -56 240 834
use sg13g2_fill_1  FILLER_97_168
timestamp 1677579658
transform 1 0 17280 0 -1 74844
box -48 -56 144 834
use sg13g2_fill_2  FILLER_97_198
timestamp 1677580104
transform 1 0 20160 0 -1 74844
box -48 -56 240 834
use sg13g2_decap_8  FILLER_98_0
timestamp 1679581782
transform 1 0 1152 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_7
timestamp 1679581782
transform 1 0 1824 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_14
timestamp 1679581782
transform 1 0 2496 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_21
timestamp 1679581782
transform 1 0 3168 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_28
timestamp 1679581782
transform 1 0 3840 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_35
timestamp 1679581782
transform 1 0 4512 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_42
timestamp 1679581782
transform 1 0 5184 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_49
timestamp 1679581782
transform 1 0 5856 0 1 74844
box -48 -56 720 834
use sg13g2_fill_1  FILLER_98_56
timestamp 1677579658
transform 1 0 6528 0 1 74844
box -48 -56 144 834
use sg13g2_decap_4  FILLER_98_77
timestamp 1679577901
transform 1 0 8544 0 1 74844
box -48 -56 432 834
use sg13g2_fill_2  FILLER_98_81
timestamp 1677580104
transform 1 0 8928 0 1 74844
box -48 -56 240 834
use sg13g2_decap_4  FILLER_98_117
timestamp 1679577901
transform 1 0 12384 0 1 74844
box -48 -56 432 834
use sg13g2_fill_2  FILLER_98_121
timestamp 1677580104
transform 1 0 12768 0 1 74844
box -48 -56 240 834
use sg13g2_decap_8  FILLER_98_140
timestamp 1679581782
transform 1 0 14592 0 1 74844
box -48 -56 720 834
use sg13g2_fill_2  FILLER_98_198
timestamp 1677580104
transform 1 0 20160 0 1 74844
box -48 -56 240 834
use sg13g2_decap_8  FILLER_99_0
timestamp 1679581782
transform 1 0 1152 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_7
timestamp 1679581782
transform 1 0 1824 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_14
timestamp 1679581782
transform 1 0 2496 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_21
timestamp 1679581782
transform 1 0 3168 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_28
timestamp 1679581782
transform 1 0 3840 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_35
timestamp 1679581782
transform 1 0 4512 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_42
timestamp 1679581782
transform 1 0 5184 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_49
timestamp 1679581782
transform 1 0 5856 0 -1 76356
box -48 -56 720 834
use sg13g2_fill_1  FILLER_99_56
timestamp 1677579658
transform 1 0 6528 0 -1 76356
box -48 -56 144 834
use sg13g2_fill_1  FILLER_99_77
timestamp 1677579658
transform 1 0 8544 0 -1 76356
box -48 -56 144 834
use sg13g2_decap_8  FILLER_99_98
timestamp 1679581782
transform 1 0 10560 0 -1 76356
box -48 -56 720 834
use sg13g2_fill_2  FILLER_99_105
timestamp 1677580104
transform 1 0 11232 0 -1 76356
box -48 -56 240 834
use sg13g2_fill_2  FILLER_99_124
timestamp 1677580104
transform 1 0 13056 0 -1 76356
box -48 -56 240 834
use sg13g2_fill_2  FILLER_99_143
timestamp 1677580104
transform 1 0 14880 0 -1 76356
box -48 -56 240 834
use sg13g2_fill_1  FILLER_99_145
timestamp 1677579658
transform 1 0 15072 0 -1 76356
box -48 -56 144 834
use sg13g2_fill_1  FILLER_99_199
timestamp 1677579658
transform 1 0 20256 0 -1 76356
box -48 -56 144 834
use sg13g2_decap_8  FILLER_100_0
timestamp 1679581782
transform 1 0 1152 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_7
timestamp 1679581782
transform 1 0 1824 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_14
timestamp 1679581782
transform 1 0 2496 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_21
timestamp 1679581782
transform 1 0 3168 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_28
timestamp 1679581782
transform 1 0 3840 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_35
timestamp 1679581782
transform 1 0 4512 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_42
timestamp 1679581782
transform 1 0 5184 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_49
timestamp 1679581782
transform 1 0 5856 0 1 76356
box -48 -56 720 834
use sg13g2_fill_1  FILLER_100_56
timestamp 1677579658
transform 1 0 6528 0 1 76356
box -48 -56 144 834
use sg13g2_decap_4  FILLER_100_116
timestamp 1679577901
transform 1 0 12288 0 1 76356
box -48 -56 432 834
use sg13g2_fill_2  FILLER_100_120
timestamp 1677580104
transform 1 0 12672 0 1 76356
box -48 -56 240 834
use sg13g2_fill_2  FILLER_100_189
timestamp 1677580104
transform 1 0 19296 0 1 76356
box -48 -56 240 834
use sg13g2_fill_1  FILLER_100_199
timestamp 1677579658
transform 1 0 20256 0 1 76356
box -48 -56 144 834
use sg13g2_decap_8  FILLER_101_0
timestamp 1679581782
transform 1 0 1152 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_7
timestamp 1679581782
transform 1 0 1824 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_14
timestamp 1679581782
transform 1 0 2496 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_21
timestamp 1679581782
transform 1 0 3168 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_28
timestamp 1679581782
transform 1 0 3840 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_35
timestamp 1679581782
transform 1 0 4512 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_42
timestamp 1679581782
transform 1 0 5184 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_49
timestamp 1679581782
transform 1 0 5856 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_56
timestamp 1679581782
transform 1 0 6528 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_63
timestamp 1679581782
transform 1 0 7200 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_4  FILLER_101_70
timestamp 1679577901
transform 1 0 7872 0 -1 77868
box -48 -56 432 834
use sg13g2_fill_2  FILLER_101_77
timestamp 1677580104
transform 1 0 8544 0 -1 77868
box -48 -56 240 834
use sg13g2_fill_2  FILLER_101_96
timestamp 1677580104
transform 1 0 10368 0 -1 77868
box -48 -56 240 834
use sg13g2_decap_8  FILLER_101_115
timestamp 1679581782
transform 1 0 12192 0 -1 77868
box -48 -56 720 834
use sg13g2_fill_1  FILLER_101_122
timestamp 1677579658
transform 1 0 12864 0 -1 77868
box -48 -56 144 834
use sg13g2_decap_4  FILLER_101_140
timestamp 1679577901
transform 1 0 14592 0 -1 77868
box -48 -56 432 834
use sg13g2_fill_2  FILLER_101_169
timestamp 1677580104
transform 1 0 17376 0 -1 77868
box -48 -56 240 834
use sg13g2_fill_1  FILLER_101_171
timestamp 1677579658
transform 1 0 17568 0 -1 77868
box -48 -56 144 834
use sg13g2_fill_2  FILLER_101_197
timestamp 1677580104
transform 1 0 20064 0 -1 77868
box -48 -56 240 834
use sg13g2_fill_1  FILLER_101_199
timestamp 1677579658
transform 1 0 20256 0 -1 77868
box -48 -56 144 834
use sg13g2_decap_8  FILLER_102_0
timestamp 1679581782
transform 1 0 1152 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_7
timestamp 1679581782
transform 1 0 1824 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_14
timestamp 1679581782
transform 1 0 2496 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_21
timestamp 1679581782
transform 1 0 3168 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_28
timestamp 1679581782
transform 1 0 3840 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_35
timestamp 1679581782
transform 1 0 4512 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_42
timestamp 1679581782
transform 1 0 5184 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_49
timestamp 1679581782
transform 1 0 5856 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_56
timestamp 1679581782
transform 1 0 6528 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_63
timestamp 1679581782
transform 1 0 7200 0 1 77868
box -48 -56 720 834
use sg13g2_decap_4  FILLER_102_70
timestamp 1679577901
transform 1 0 7872 0 1 77868
box -48 -56 432 834
use sg13g2_decap_8  FILLER_102_77
timestamp 1679581782
transform 1 0 8544 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_84
timestamp 1679581782
transform 1 0 9216 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_91
timestamp 1679581782
transform 1 0 9888 0 1 77868
box -48 -56 720 834
use sg13g2_fill_1  FILLER_102_98
timestamp 1677579658
transform 1 0 10560 0 1 77868
box -48 -56 144 834
use sg13g2_decap_8  FILLER_102_102
timestamp 1679581782
transform 1 0 10944 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_126
timestamp 1679581782
transform 1 0 13248 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_133
timestamp 1679581782
transform 1 0 13920 0 1 77868
box -48 -56 720 834
use sg13g2_fill_2  FILLER_102_140
timestamp 1677580104
transform 1 0 14592 0 1 77868
box -48 -56 240 834
use sg13g2_decap_8  FILLER_102_163
timestamp 1679581782
transform 1 0 16800 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_170
timestamp 1679581782
transform 1 0 17472 0 1 77868
box -48 -56 720 834
use sg13g2_decap_4  FILLER_102_177
timestamp 1679577901
transform 1 0 18144 0 1 77868
box -48 -56 432 834
use sg13g2_fill_2  FILLER_102_197
timestamp 1677580104
transform 1 0 20064 0 1 77868
box -48 -56 240 834
use sg13g2_fill_1  FILLER_102_199
timestamp 1677579658
transform 1 0 20256 0 1 77868
box -48 -56 144 834
use sg13g2_decap_8  FILLER_103_0
timestamp 1679581782
transform 1 0 1152 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_7
timestamp 1679581782
transform 1 0 1824 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_14
timestamp 1679581782
transform 1 0 2496 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_21
timestamp 1679581782
transform 1 0 3168 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_28
timestamp 1679581782
transform 1 0 3840 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_35
timestamp 1679581782
transform 1 0 4512 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_42
timestamp 1679581782
transform 1 0 5184 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_49
timestamp 1679581782
transform 1 0 5856 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_56
timestamp 1679581782
transform 1 0 6528 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_63
timestamp 1679581782
transform 1 0 7200 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_70
timestamp 1679581782
transform 1 0 7872 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_4  FILLER_103_77
timestamp 1679577901
transform 1 0 8544 0 -1 79380
box -48 -56 432 834
use sg13g2_fill_1  FILLER_103_81
timestamp 1677579658
transform 1 0 8928 0 -1 79380
box -48 -56 144 834
use sg13g2_fill_2  FILLER_103_120
timestamp 1677580104
transform 1 0 12672 0 -1 79380
box -48 -56 240 834
use sg13g2_fill_1  FILLER_103_122
timestamp 1677579658
transform 1 0 12864 0 -1 79380
box -48 -56 144 834
use sg13g2_fill_2  FILLER_103_144
timestamp 1677580104
transform 1 0 14976 0 -1 79380
box -48 -56 240 834
use sg13g2_fill_1  FILLER_103_146
timestamp 1677579658
transform 1 0 15168 0 -1 79380
box -48 -56 144 834
use sg13g2_decap_8  FILLER_103_164
timestamp 1679581782
transform 1 0 16896 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_171
timestamp 1679581782
transform 1 0 17568 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_178
timestamp 1679581782
transform 1 0 18240 0 -1 79380
box -48 -56 720 834
use sg13g2_fill_2  FILLER_103_197
timestamp 1677580104
transform 1 0 20064 0 -1 79380
box -48 -56 240 834
use sg13g2_fill_1  FILLER_103_199
timestamp 1677579658
transform 1 0 20256 0 -1 79380
box -48 -56 144 834
use sg13g2_decap_8  FILLER_104_0
timestamp 1679581782
transform 1 0 1152 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_7
timestamp 1679581782
transform 1 0 1824 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_14
timestamp 1679581782
transform 1 0 2496 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_21
timestamp 1679581782
transform 1 0 3168 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_28
timestamp 1679581782
transform 1 0 3840 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_35
timestamp 1679581782
transform 1 0 4512 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_42
timestamp 1679581782
transform 1 0 5184 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_49
timestamp 1679581782
transform 1 0 5856 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_56
timestamp 1679581782
transform 1 0 6528 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_63
timestamp 1679581782
transform 1 0 7200 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_70
timestamp 1679581782
transform 1 0 7872 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_77
timestamp 1679581782
transform 1 0 8544 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_84
timestamp 1679581782
transform 1 0 9216 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_91
timestamp 1679581782
transform 1 0 9888 0 1 79380
box -48 -56 720 834
use sg13g2_fill_1  FILLER_104_98
timestamp 1677579658
transform 1 0 10560 0 1 79380
box -48 -56 144 834
use sg13g2_decap_8  FILLER_104_119
timestamp 1679581782
transform 1 0 12576 0 1 79380
box -48 -56 720 834
use sg13g2_fill_1  FILLER_104_126
timestamp 1677579658
transform 1 0 13248 0 1 79380
box -48 -56 144 834
use sg13g2_decap_4  FILLER_104_144
timestamp 1679577901
transform 1 0 14976 0 1 79380
box -48 -56 432 834
use sg13g2_fill_1  FILLER_104_148
timestamp 1677579658
transform 1 0 15360 0 1 79380
box -48 -56 144 834
use sg13g2_fill_2  FILLER_104_157
timestamp 1677580104
transform 1 0 16224 0 1 79380
box -48 -56 240 834
use sg13g2_decap_8  FILLER_104_163
timestamp 1679581782
transform 1 0 16800 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_170
timestamp 1679581782
transform 1 0 17472 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_177
timestamp 1679581782
transform 1 0 18144 0 1 79380
box -48 -56 720 834
use sg13g2_fill_1  FILLER_104_184
timestamp 1677579658
transform 1 0 18816 0 1 79380
box -48 -56 144 834
use sg13g2_fill_2  FILLER_104_197
timestamp 1677580104
transform 1 0 20064 0 1 79380
box -48 -56 240 834
use sg13g2_fill_1  FILLER_104_199
timestamp 1677579658
transform 1 0 20256 0 1 79380
box -48 -56 144 834
use sg13g2_decap_8  FILLER_105_0
timestamp 1679581782
transform 1 0 1152 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_7
timestamp 1679581782
transform 1 0 1824 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_14
timestamp 1679581782
transform 1 0 2496 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_21
timestamp 1679581782
transform 1 0 3168 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_28
timestamp 1679581782
transform 1 0 3840 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_35
timestamp 1679581782
transform 1 0 4512 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_42
timestamp 1679581782
transform 1 0 5184 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_49
timestamp 1679581782
transform 1 0 5856 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_56
timestamp 1679581782
transform 1 0 6528 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_63
timestamp 1679581782
transform 1 0 7200 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_70
timestamp 1679581782
transform 1 0 7872 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_77
timestamp 1679581782
transform 1 0 8544 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_84
timestamp 1679581782
transform 1 0 9216 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_91
timestamp 1679581782
transform 1 0 9888 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_98
timestamp 1679581782
transform 1 0 10560 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_105
timestamp 1679581782
transform 1 0 11232 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_112
timestamp 1679581782
transform 1 0 11904 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_4  FILLER_105_119
timestamp 1679577901
transform 1 0 12576 0 -1 80892
box -48 -56 432 834
use sg13g2_fill_2  FILLER_105_123
timestamp 1677580104
transform 1 0 12960 0 -1 80892
box -48 -56 240 834
use sg13g2_decap_8  FILLER_105_142
timestamp 1679581782
transform 1 0 14784 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_149
timestamp 1679581782
transform 1 0 15456 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_156
timestamp 1679581782
transform 1 0 16128 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_163
timestamp 1679581782
transform 1 0 16800 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_170
timestamp 1679581782
transform 1 0 17472 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_4  FILLER_105_177
timestamp 1679577901
transform 1 0 18144 0 -1 80892
box -48 -56 432 834
use sg13g2_fill_1  FILLER_105_181
timestamp 1677579658
transform 1 0 18528 0 -1 80892
box -48 -56 144 834
use sg13g2_fill_2  FILLER_105_186
timestamp 1677580104
transform 1 0 19008 0 -1 80892
box -48 -56 240 834
use sg13g2_fill_1  FILLER_105_188
timestamp 1677579658
transform 1 0 19200 0 -1 80892
box -48 -56 144 834
use sg13g2_fill_2  FILLER_105_197
timestamp 1677580104
transform 1 0 20064 0 -1 80892
box -48 -56 240 834
use sg13g2_fill_1  FILLER_105_199
timestamp 1677579658
transform 1 0 20256 0 -1 80892
box -48 -56 144 834
use sg13g2_decap_8  FILLER_106_0
timestamp 1679581782
transform 1 0 1152 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_7
timestamp 1679581782
transform 1 0 1824 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_14
timestamp 1679581782
transform 1 0 2496 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_21
timestamp 1679581782
transform 1 0 3168 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_28
timestamp 1679581782
transform 1 0 3840 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_35
timestamp 1679581782
transform 1 0 4512 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_42
timestamp 1679581782
transform 1 0 5184 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_49
timestamp 1679581782
transform 1 0 5856 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_56
timestamp 1679581782
transform 1 0 6528 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_63
timestamp 1679581782
transform 1 0 7200 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_70
timestamp 1679581782
transform 1 0 7872 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_77
timestamp 1679581782
transform 1 0 8544 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_84
timestamp 1679581782
transform 1 0 9216 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_91
timestamp 1679581782
transform 1 0 9888 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_98
timestamp 1679581782
transform 1 0 10560 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_105
timestamp 1679581782
transform 1 0 11232 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_112
timestamp 1679581782
transform 1 0 11904 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_119
timestamp 1679581782
transform 1 0 12576 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_126
timestamp 1679581782
transform 1 0 13248 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_133
timestamp 1679581782
transform 1 0 13920 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_140
timestamp 1679581782
transform 1 0 14592 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_147
timestamp 1679581782
transform 1 0 15264 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_154
timestamp 1679581782
transform 1 0 15936 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_161
timestamp 1679581782
transform 1 0 16608 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_168
timestamp 1679581782
transform 1 0 17280 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_175
timestamp 1679581782
transform 1 0 17952 0 1 80892
box -48 -56 720 834
use sg13g2_fill_2  FILLER_106_182
timestamp 1677580104
transform 1 0 18624 0 1 80892
box -48 -56 240 834
use sg13g2_fill_1  FILLER_106_184
timestamp 1677579658
transform 1 0 18816 0 1 80892
box -48 -56 144 834
use sg13g2_decap_8  FILLER_106_193
timestamp 1679581782
transform 1 0 19680 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_0
timestamp 1679581782
transform 1 0 1152 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_7
timestamp 1679581782
transform 1 0 1824 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_14
timestamp 1679581782
transform 1 0 2496 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_21
timestamp 1679581782
transform 1 0 3168 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_28
timestamp 1679581782
transform 1 0 3840 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_35
timestamp 1679581782
transform 1 0 4512 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_42
timestamp 1679581782
transform 1 0 5184 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_49
timestamp 1679581782
transform 1 0 5856 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_56
timestamp 1679581782
transform 1 0 6528 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_63
timestamp 1679581782
transform 1 0 7200 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_70
timestamp 1679581782
transform 1 0 7872 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_77
timestamp 1679581782
transform 1 0 8544 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_84
timestamp 1679581782
transform 1 0 9216 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_91
timestamp 1679581782
transform 1 0 9888 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_98
timestamp 1679581782
transform 1 0 10560 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_105
timestamp 1679581782
transform 1 0 11232 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_112
timestamp 1679581782
transform 1 0 11904 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_119
timestamp 1679581782
transform 1 0 12576 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_126
timestamp 1679581782
transform 1 0 13248 0 -1 82404
box -48 -56 720 834
use sg13g2_fill_1  FILLER_107_133
timestamp 1677579658
transform 1 0 13920 0 -1 82404
box -48 -56 144 834
use sg13g2_decap_8  FILLER_107_138
timestamp 1679581782
transform 1 0 14400 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_4  FILLER_107_145
timestamp 1679577901
transform 1 0 15072 0 -1 82404
box -48 -56 432 834
use sg13g2_decap_8  FILLER_107_153
timestamp 1679581782
transform 1 0 15840 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_160
timestamp 1679581782
transform 1 0 16512 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_167
timestamp 1679581782
transform 1 0 17184 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_174
timestamp 1679581782
transform 1 0 17856 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_181
timestamp 1679581782
transform 1 0 18528 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_188
timestamp 1679581782
transform 1 0 19200 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_4  FILLER_107_195
timestamp 1679577901
transform 1 0 19872 0 -1 82404
box -48 -56 432 834
use sg13g2_fill_1  FILLER_107_199
timestamp 1677579658
transform 1 0 20256 0 -1 82404
box -48 -56 144 834
use sg13g2_decap_8  FILLER_108_0
timestamp 1679581782
transform 1 0 1152 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_7
timestamp 1679581782
transform 1 0 1824 0 1 82404
box -48 -56 720 834
use sg13g2_fill_1  FILLER_108_14
timestamp 1677579658
transform 1 0 2496 0 1 82404
box -48 -56 144 834
use sg13g2_fill_1  FILLER_108_27
timestamp 1677579658
transform 1 0 3744 0 1 82404
box -48 -56 144 834
use sg13g2_fill_2  FILLER_108_32
timestamp 1677580104
transform 1 0 4224 0 1 82404
box -48 -56 240 834
use sg13g2_fill_1  FILLER_108_34
timestamp 1677579658
transform 1 0 4416 0 1 82404
box -48 -56 144 834
use sg13g2_decap_8  FILLER_108_39
timestamp 1679581782
transform 1 0 4896 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_46
timestamp 1679581782
transform 1 0 5568 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_53
timestamp 1679581782
transform 1 0 6240 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_60
timestamp 1679581782
transform 1 0 6912 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_67
timestamp 1679581782
transform 1 0 7584 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_74
timestamp 1679581782
transform 1 0 8256 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_81
timestamp 1679581782
transform 1 0 8928 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_88
timestamp 1679581782
transform 1 0 9600 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_95
timestamp 1679581782
transform 1 0 10272 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_102
timestamp 1679581782
transform 1 0 10944 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_109
timestamp 1679581782
transform 1 0 11616 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_116
timestamp 1679581782
transform 1 0 12288 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_123
timestamp 1679581782
transform 1 0 12960 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_130
timestamp 1679581782
transform 1 0 13632 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_137
timestamp 1679581782
transform 1 0 14304 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_144
timestamp 1679581782
transform 1 0 14976 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_151
timestamp 1679581782
transform 1 0 15648 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_158
timestamp 1679581782
transform 1 0 16320 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_165
timestamp 1679581782
transform 1 0 16992 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_172
timestamp 1679581782
transform 1 0 17664 0 1 82404
box -48 -56 720 834
use sg13g2_decap_4  FILLER_108_179
timestamp 1679577901
transform 1 0 18336 0 1 82404
box -48 -56 432 834
use sg13g2_fill_2  FILLER_108_183
timestamp 1677580104
transform 1 0 18720 0 1 82404
box -48 -56 240 834
use sg13g2_decap_8  FILLER_108_193
timestamp 1679581782
transform 1 0 19680 0 1 82404
box -48 -56 720 834
use sg13g2_fill_2  FILLER_109_0
timestamp 1677580104
transform 1 0 1152 0 -1 83916
box -48 -56 240 834
use sg13g2_fill_1  FILLER_109_2
timestamp 1677579658
transform 1 0 1344 0 -1 83916
box -48 -56 144 834
use sg13g2_fill_2  FILLER_109_47
timestamp 1677580104
transform 1 0 5664 0 -1 83916
box -48 -56 240 834
use sg13g2_fill_2  FILLER_109_53
timestamp 1677580104
transform 1 0 6240 0 -1 83916
box -48 -56 240 834
use sg13g2_fill_1  FILLER_109_59
timestamp 1677579658
transform 1 0 6816 0 -1 83916
box -48 -56 144 834
use sg13g2_decap_8  FILLER_109_80
timestamp 1679581782
transform 1 0 8832 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_109_87
timestamp 1679581782
transform 1 0 9504 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_109_94
timestamp 1679581782
transform 1 0 10176 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_109_101
timestamp 1679581782
transform 1 0 10848 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_109_108
timestamp 1679581782
transform 1 0 11520 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_109_115
timestamp 1679581782
transform 1 0 12192 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_4  FILLER_109_122
timestamp 1679577901
transform 1 0 12864 0 -1 83916
box -48 -56 432 834
use sg13g2_decap_8  FILLER_109_130
timestamp 1679581782
transform 1 0 13632 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_4  FILLER_109_137
timestamp 1679577901
transform 1 0 14304 0 -1 83916
box -48 -56 432 834
use sg13g2_fill_2  FILLER_109_141
timestamp 1677580104
transform 1 0 14688 0 -1 83916
box -48 -56 240 834
use sg13g2_decap_8  FILLER_109_155
timestamp 1679581782
transform 1 0 16032 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_109_162
timestamp 1679581782
transform 1 0 16704 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_109_169
timestamp 1679581782
transform 1 0 17376 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_4  FILLER_109_180
timestamp 1679577901
transform 1 0 18432 0 -1 83916
box -48 -56 432 834
use sg13g2_fill_1  FILLER_109_184
timestamp 1677579658
transform 1 0 18816 0 -1 83916
box -48 -56 144 834
use sg13g2_decap_8  FILLER_109_193
timestamp 1679581782
transform 1 0 19680 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_0
timestamp 1679581782
transform 1 0 1152 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_7
timestamp 1679581782
transform 1 0 1824 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_14
timestamp 1679581782
transform 1 0 2496 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_21
timestamp 1679581782
transform 1 0 3168 0 1 83916
box -48 -56 720 834
use sg13g2_decap_4  FILLER_110_28
timestamp 1679577901
transform 1 0 3840 0 1 83916
box -48 -56 432 834
use sg13g2_decap_8  FILLER_110_36
timestamp 1679581782
transform 1 0 4608 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_43
timestamp 1679581782
transform 1 0 5280 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_50
timestamp 1679581782
transform 1 0 5952 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_57
timestamp 1679581782
transform 1 0 6624 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_64
timestamp 1679581782
transform 1 0 7296 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_71
timestamp 1679581782
transform 1 0 7968 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_78
timestamp 1679581782
transform 1 0 8640 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_85
timestamp 1679581782
transform 1 0 9312 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_92
timestamp 1679581782
transform 1 0 9984 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_99
timestamp 1679581782
transform 1 0 10656 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_106
timestamp 1679581782
transform 1 0 11328 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_113
timestamp 1679581782
transform 1 0 12000 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_120
timestamp 1679581782
transform 1 0 12672 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_127
timestamp 1679581782
transform 1 0 13344 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_134
timestamp 1679581782
transform 1 0 14016 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_141
timestamp 1679581782
transform 1 0 14688 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_148
timestamp 1679581782
transform 1 0 15360 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_155
timestamp 1679581782
transform 1 0 16032 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_162
timestamp 1679581782
transform 1 0 16704 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_169
timestamp 1679581782
transform 1 0 17376 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_176
timestamp 1679581782
transform 1 0 18048 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_183
timestamp 1679581782
transform 1 0 18720 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_190
timestamp 1679581782
transform 1 0 19392 0 1 83916
box -48 -56 720 834
use sg13g2_fill_2  FILLER_110_197
timestamp 1677580104
transform 1 0 20064 0 1 83916
box -48 -56 240 834
use sg13g2_fill_1  FILLER_110_199
timestamp 1677579658
transform 1 0 20256 0 1 83916
box -48 -56 144 834
<< labels >>
flabel metal3 s 0 34820 80 34900 0 FreeSans 320 0 0 0 CLK_TT_PROJECT
port 0 nsew signal output
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 ENA_TT_PROJECT
port 1 nsew signal output
flabel metal3 s 0 35492 80 35572 0 FreeSans 320 0 0 0 RST_N_TT_PROJECT
port 2 nsew signal output
flabel metal3 s 21424 59180 21504 59260 0 FreeSans 320 0 0 0 Tile_X0Y0_E1BEG[0]
port 3 nsew signal output
flabel metal3 s 21424 59516 21504 59596 0 FreeSans 320 0 0 0 Tile_X0Y0_E1BEG[1]
port 4 nsew signal output
flabel metal3 s 21424 59852 21504 59932 0 FreeSans 320 0 0 0 Tile_X0Y0_E1BEG[2]
port 5 nsew signal output
flabel metal3 s 21424 60188 21504 60268 0 FreeSans 320 0 0 0 Tile_X0Y0_E1BEG[3]
port 6 nsew signal output
flabel metal3 s 21424 60524 21504 60604 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEG[0]
port 7 nsew signal output
flabel metal3 s 21424 60860 21504 60940 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEG[1]
port 8 nsew signal output
flabel metal3 s 21424 61196 21504 61276 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEG[2]
port 9 nsew signal output
flabel metal3 s 21424 61532 21504 61612 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEG[3]
port 10 nsew signal output
flabel metal3 s 21424 61868 21504 61948 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEG[4]
port 11 nsew signal output
flabel metal3 s 21424 62204 21504 62284 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEG[5]
port 12 nsew signal output
flabel metal3 s 21424 62540 21504 62620 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEG[6]
port 13 nsew signal output
flabel metal3 s 21424 62876 21504 62956 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEG[7]
port 14 nsew signal output
flabel metal3 s 21424 63212 21504 63292 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEGb[0]
port 15 nsew signal output
flabel metal3 s 21424 63548 21504 63628 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEGb[1]
port 16 nsew signal output
flabel metal3 s 21424 63884 21504 63964 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEGb[2]
port 17 nsew signal output
flabel metal3 s 21424 64220 21504 64300 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEGb[3]
port 18 nsew signal output
flabel metal3 s 21424 64556 21504 64636 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEGb[4]
port 19 nsew signal output
flabel metal3 s 21424 64892 21504 64972 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEGb[5]
port 20 nsew signal output
flabel metal3 s 21424 65228 21504 65308 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEGb[6]
port 21 nsew signal output
flabel metal3 s 21424 65564 21504 65644 0 FreeSans 320 0 0 0 Tile_X0Y0_E2BEGb[7]
port 22 nsew signal output
flabel metal3 s 21424 71276 21504 71356 0 FreeSans 320 0 0 0 Tile_X0Y0_E6BEG[0]
port 23 nsew signal output
flabel metal3 s 21424 74636 21504 74716 0 FreeSans 320 0 0 0 Tile_X0Y0_E6BEG[10]
port 24 nsew signal output
flabel metal3 s 21424 74972 21504 75052 0 FreeSans 320 0 0 0 Tile_X0Y0_E6BEG[11]
port 25 nsew signal output
flabel metal3 s 21424 71612 21504 71692 0 FreeSans 320 0 0 0 Tile_X0Y0_E6BEG[1]
port 26 nsew signal output
flabel metal3 s 21424 71948 21504 72028 0 FreeSans 320 0 0 0 Tile_X0Y0_E6BEG[2]
port 27 nsew signal output
flabel metal3 s 21424 72284 21504 72364 0 FreeSans 320 0 0 0 Tile_X0Y0_E6BEG[3]
port 28 nsew signal output
flabel metal3 s 21424 72620 21504 72700 0 FreeSans 320 0 0 0 Tile_X0Y0_E6BEG[4]
port 29 nsew signal output
flabel metal3 s 21424 72956 21504 73036 0 FreeSans 320 0 0 0 Tile_X0Y0_E6BEG[5]
port 30 nsew signal output
flabel metal3 s 21424 73292 21504 73372 0 FreeSans 320 0 0 0 Tile_X0Y0_E6BEG[6]
port 31 nsew signal output
flabel metal3 s 21424 73628 21504 73708 0 FreeSans 320 0 0 0 Tile_X0Y0_E6BEG[7]
port 32 nsew signal output
flabel metal3 s 21424 73964 21504 74044 0 FreeSans 320 0 0 0 Tile_X0Y0_E6BEG[8]
port 33 nsew signal output
flabel metal3 s 21424 74300 21504 74380 0 FreeSans 320 0 0 0 Tile_X0Y0_E6BEG[9]
port 34 nsew signal output
flabel metal3 s 21424 65900 21504 65980 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[0]
port 35 nsew signal output
flabel metal3 s 21424 69260 21504 69340 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[10]
port 36 nsew signal output
flabel metal3 s 21424 69596 21504 69676 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[11]
port 37 nsew signal output
flabel metal3 s 21424 69932 21504 70012 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[12]
port 38 nsew signal output
flabel metal3 s 21424 70268 21504 70348 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[13]
port 39 nsew signal output
flabel metal3 s 21424 70604 21504 70684 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[14]
port 40 nsew signal output
flabel metal3 s 21424 70940 21504 71020 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[15]
port 41 nsew signal output
flabel metal3 s 21424 66236 21504 66316 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[1]
port 42 nsew signal output
flabel metal3 s 21424 66572 21504 66652 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[2]
port 43 nsew signal output
flabel metal3 s 21424 66908 21504 66988 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[3]
port 44 nsew signal output
flabel metal3 s 21424 67244 21504 67324 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[4]
port 45 nsew signal output
flabel metal3 s 21424 67580 21504 67660 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[5]
port 46 nsew signal output
flabel metal3 s 21424 67916 21504 67996 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[6]
port 47 nsew signal output
flabel metal3 s 21424 68252 21504 68332 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[7]
port 48 nsew signal output
flabel metal3 s 21424 68588 21504 68668 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[8]
port 49 nsew signal output
flabel metal3 s 21424 68924 21504 69004 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4BEG[9]
port 50 nsew signal output
flabel metal3 s 0 36164 80 36244 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[0]
port 51 nsew signal input
flabel metal3 s 0 42884 80 42964 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[10]
port 52 nsew signal input
flabel metal3 s 0 43556 80 43636 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[11]
port 53 nsew signal input
flabel metal3 s 0 44228 80 44308 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[12]
port 54 nsew signal input
flabel metal3 s 0 44900 80 44980 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[13]
port 55 nsew signal input
flabel metal3 s 0 45572 80 45652 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[14]
port 56 nsew signal input
flabel metal3 s 0 46244 80 46324 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[15]
port 57 nsew signal input
flabel metal3 s 0 46916 80 46996 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[16]
port 58 nsew signal input
flabel metal3 s 0 47588 80 47668 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[17]
port 59 nsew signal input
flabel metal3 s 0 48260 80 48340 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[18]
port 60 nsew signal input
flabel metal3 s 0 48932 80 49012 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[19]
port 61 nsew signal input
flabel metal3 s 0 36836 80 36916 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[1]
port 62 nsew signal input
flabel metal3 s 0 49604 80 49684 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[20]
port 63 nsew signal input
flabel metal3 s 0 50276 80 50356 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[21]
port 64 nsew signal input
flabel metal3 s 0 50948 80 51028 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[22]
port 65 nsew signal input
flabel metal3 s 0 51620 80 51700 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[23]
port 66 nsew signal input
flabel metal3 s 0 52292 80 52372 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[24]
port 67 nsew signal input
flabel metal3 s 0 52964 80 53044 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[25]
port 68 nsew signal input
flabel metal3 s 0 53636 80 53716 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[26]
port 69 nsew signal input
flabel metal3 s 0 54308 80 54388 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[27]
port 70 nsew signal input
flabel metal3 s 0 54980 80 55060 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[28]
port 71 nsew signal input
flabel metal3 s 0 55652 80 55732 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[29]
port 72 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[2]
port 73 nsew signal input
flabel metal3 s 0 56324 80 56404 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[30]
port 74 nsew signal input
flabel metal3 s 0 56996 80 57076 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[31]
port 75 nsew signal input
flabel metal3 s 0 38180 80 38260 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[3]
port 76 nsew signal input
flabel metal3 s 0 38852 80 38932 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[4]
port 77 nsew signal input
flabel metal3 s 0 39524 80 39604 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[5]
port 78 nsew signal input
flabel metal3 s 0 40196 80 40276 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[6]
port 79 nsew signal input
flabel metal3 s 0 40868 80 40948 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[7]
port 80 nsew signal input
flabel metal3 s 0 41540 80 41620 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[8]
port 81 nsew signal input
flabel metal3 s 0 42212 80 42292 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[9]
port 82 nsew signal input
flabel metal3 s 21424 75308 21504 75388 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[0]
port 83 nsew signal output
flabel metal3 s 21424 78668 21504 78748 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[10]
port 84 nsew signal output
flabel metal3 s 21424 79004 21504 79084 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[11]
port 85 nsew signal output
flabel metal3 s 21424 79340 21504 79420 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[12]
port 86 nsew signal output
flabel metal3 s 21424 79676 21504 79756 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[13]
port 87 nsew signal output
flabel metal3 s 21424 80012 21504 80092 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[14]
port 88 nsew signal output
flabel metal3 s 21424 80348 21504 80428 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[15]
port 89 nsew signal output
flabel metal3 s 21424 80684 21504 80764 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[16]
port 90 nsew signal output
flabel metal3 s 21424 81020 21504 81100 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[17]
port 91 nsew signal output
flabel metal3 s 21424 81356 21504 81436 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[18]
port 92 nsew signal output
flabel metal3 s 21424 81692 21504 81772 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[19]
port 93 nsew signal output
flabel metal3 s 21424 75644 21504 75724 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[1]
port 94 nsew signal output
flabel metal3 s 21424 82028 21504 82108 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[20]
port 95 nsew signal output
flabel metal3 s 21424 82364 21504 82444 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[21]
port 96 nsew signal output
flabel metal3 s 21424 82700 21504 82780 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[22]
port 97 nsew signal output
flabel metal3 s 21424 83036 21504 83116 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[23]
port 98 nsew signal output
flabel metal3 s 21424 83372 21504 83452 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[24]
port 99 nsew signal output
flabel metal3 s 21424 83708 21504 83788 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[25]
port 100 nsew signal output
flabel metal3 s 21424 84044 21504 84124 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[26]
port 101 nsew signal output
flabel metal3 s 21424 84380 21504 84460 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[27]
port 102 nsew signal output
flabel metal3 s 21424 84716 21504 84796 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[28]
port 103 nsew signal output
flabel metal3 s 21424 85052 21504 85132 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[29]
port 104 nsew signal output
flabel metal3 s 21424 75980 21504 76060 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[2]
port 105 nsew signal output
flabel metal3 s 21424 85388 21504 85468 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[30]
port 106 nsew signal output
flabel metal3 s 21424 85724 21504 85804 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[31]
port 107 nsew signal output
flabel metal3 s 21424 76316 21504 76396 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[3]
port 108 nsew signal output
flabel metal3 s 21424 76652 21504 76732 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[4]
port 109 nsew signal output
flabel metal3 s 21424 76988 21504 77068 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[5]
port 110 nsew signal output
flabel metal3 s 21424 77324 21504 77404 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[6]
port 111 nsew signal output
flabel metal3 s 21424 77660 21504 77740 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[7]
port 112 nsew signal output
flabel metal3 s 21424 77996 21504 78076 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[8]
port 113 nsew signal output
flabel metal3 s 21424 78332 21504 78412 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[9]
port 114 nsew signal output
flabel metal2 s 15800 85936 15880 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[0]
port 115 nsew signal output
flabel metal2 s 17720 85936 17800 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[10]
port 116 nsew signal output
flabel metal2 s 17912 85936 17992 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[11]
port 117 nsew signal output
flabel metal2 s 18104 85936 18184 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[12]
port 118 nsew signal output
flabel metal2 s 18296 85936 18376 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[13]
port 119 nsew signal output
flabel metal2 s 18488 85936 18568 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[14]
port 120 nsew signal output
flabel metal2 s 18680 85936 18760 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[15]
port 121 nsew signal output
flabel metal2 s 18872 85936 18952 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[16]
port 122 nsew signal output
flabel metal2 s 19064 85936 19144 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[17]
port 123 nsew signal output
flabel metal2 s 19256 85936 19336 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[18]
port 124 nsew signal output
flabel metal2 s 19448 85936 19528 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[19]
port 125 nsew signal output
flabel metal2 s 15992 85936 16072 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[1]
port 126 nsew signal output
flabel metal2 s 16184 85936 16264 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[2]
port 127 nsew signal output
flabel metal2 s 16376 85936 16456 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[3]
port 128 nsew signal output
flabel metal2 s 16568 85936 16648 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[4]
port 129 nsew signal output
flabel metal2 s 16760 85936 16840 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[5]
port 130 nsew signal output
flabel metal2 s 16952 85936 17032 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[6]
port 131 nsew signal output
flabel metal2 s 17144 85936 17224 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[7]
port 132 nsew signal output
flabel metal2 s 17336 85936 17416 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[8]
port 133 nsew signal output
flabel metal2 s 17528 85936 17608 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[9]
port 134 nsew signal output
flabel metal2 s 1784 85936 1864 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[0]
port 135 nsew signal output
flabel metal2 s 1976 85936 2056 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[1]
port 136 nsew signal output
flabel metal2 s 2168 85936 2248 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[2]
port 137 nsew signal output
flabel metal2 s 2360 85936 2440 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[3]
port 138 nsew signal output
flabel metal2 s 2552 85936 2632 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[0]
port 139 nsew signal output
flabel metal2 s 2744 85936 2824 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[1]
port 140 nsew signal output
flabel metal2 s 2936 85936 3016 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[2]
port 141 nsew signal output
flabel metal2 s 3128 85936 3208 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[3]
port 142 nsew signal output
flabel metal2 s 3320 85936 3400 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[4]
port 143 nsew signal output
flabel metal2 s 3512 85936 3592 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[5]
port 144 nsew signal output
flabel metal2 s 3704 85936 3784 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[6]
port 145 nsew signal output
flabel metal2 s 3896 85936 3976 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[7]
port 146 nsew signal output
flabel metal2 s 4088 85936 4168 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[0]
port 147 nsew signal output
flabel metal2 s 4280 85936 4360 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[1]
port 148 nsew signal output
flabel metal2 s 4472 85936 4552 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[2]
port 149 nsew signal output
flabel metal2 s 4664 85936 4744 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[3]
port 150 nsew signal output
flabel metal2 s 4856 85936 4936 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[4]
port 151 nsew signal output
flabel metal2 s 5048 85936 5128 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[5]
port 152 nsew signal output
flabel metal2 s 5240 85936 5320 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[6]
port 153 nsew signal output
flabel metal2 s 5432 85936 5512 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[7]
port 154 nsew signal output
flabel metal2 s 5624 85936 5704 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[0]
port 155 nsew signal output
flabel metal2 s 7544 85936 7624 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[10]
port 156 nsew signal output
flabel metal2 s 7736 85936 7816 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[11]
port 157 nsew signal output
flabel metal2 s 7928 85936 8008 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[12]
port 158 nsew signal output
flabel metal2 s 8120 85936 8200 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[13]
port 159 nsew signal output
flabel metal2 s 8312 85936 8392 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[14]
port 160 nsew signal output
flabel metal2 s 8504 85936 8584 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[15]
port 161 nsew signal output
flabel metal2 s 5816 85936 5896 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[1]
port 162 nsew signal output
flabel metal2 s 6008 85936 6088 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[2]
port 163 nsew signal output
flabel metal2 s 6200 85936 6280 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[3]
port 164 nsew signal output
flabel metal2 s 6392 85936 6472 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[4]
port 165 nsew signal output
flabel metal2 s 6584 85936 6664 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[5]
port 166 nsew signal output
flabel metal2 s 6776 85936 6856 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[6]
port 167 nsew signal output
flabel metal2 s 6968 85936 7048 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[7]
port 168 nsew signal output
flabel metal2 s 7160 85936 7240 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[8]
port 169 nsew signal output
flabel metal2 s 7352 85936 7432 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[9]
port 170 nsew signal output
flabel metal2 s 8696 85936 8776 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[0]
port 171 nsew signal input
flabel metal2 s 8888 85936 8968 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[1]
port 172 nsew signal input
flabel metal2 s 9080 85936 9160 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[2]
port 173 nsew signal input
flabel metal2 s 9272 85936 9352 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[3]
port 174 nsew signal input
flabel metal2 s 11000 85936 11080 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[0]
port 175 nsew signal input
flabel metal2 s 11192 85936 11272 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[1]
port 176 nsew signal input
flabel metal2 s 11384 85936 11464 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[2]
port 177 nsew signal input
flabel metal2 s 11576 85936 11656 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[3]
port 178 nsew signal input
flabel metal2 s 11768 85936 11848 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[4]
port 179 nsew signal input
flabel metal2 s 11960 85936 12040 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[5]
port 180 nsew signal input
flabel metal2 s 12152 85936 12232 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[6]
port 181 nsew signal input
flabel metal2 s 12344 85936 12424 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[7]
port 182 nsew signal input
flabel metal2 s 9464 85936 9544 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[0]
port 183 nsew signal input
flabel metal2 s 9656 85936 9736 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[1]
port 184 nsew signal input
flabel metal2 s 9848 85936 9928 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[2]
port 185 nsew signal input
flabel metal2 s 10040 85936 10120 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[3]
port 186 nsew signal input
flabel metal2 s 10232 85936 10312 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[4]
port 187 nsew signal input
flabel metal2 s 10424 85936 10504 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[5]
port 188 nsew signal input
flabel metal2 s 10616 85936 10696 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[6]
port 189 nsew signal input
flabel metal2 s 10808 85936 10888 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[7]
port 190 nsew signal input
flabel metal2 s 12536 85936 12616 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[0]
port 191 nsew signal input
flabel metal2 s 14456 85936 14536 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[10]
port 192 nsew signal input
flabel metal2 s 14648 85936 14728 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[11]
port 193 nsew signal input
flabel metal2 s 14840 85936 14920 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[12]
port 194 nsew signal input
flabel metal2 s 15032 85936 15112 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[13]
port 195 nsew signal input
flabel metal2 s 15224 85936 15304 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[14]
port 196 nsew signal input
flabel metal2 s 15416 85936 15496 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[15]
port 197 nsew signal input
flabel metal2 s 12728 85936 12808 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[1]
port 198 nsew signal input
flabel metal2 s 12920 85936 13000 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[2]
port 199 nsew signal input
flabel metal2 s 13112 85936 13192 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[3]
port 200 nsew signal input
flabel metal2 s 13304 85936 13384 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[4]
port 201 nsew signal input
flabel metal2 s 13496 85936 13576 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[5]
port 202 nsew signal input
flabel metal2 s 13688 85936 13768 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[6]
port 203 nsew signal input
flabel metal2 s 13880 85936 13960 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[7]
port 204 nsew signal input
flabel metal2 s 14072 85936 14152 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[8]
port 205 nsew signal input
flabel metal2 s 14264 85936 14344 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[9]
port 206 nsew signal input
flabel metal2 s 15608 85936 15688 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_UserCLKo
port 207 nsew signal output
flabel metal3 s 21424 43052 21504 43132 0 FreeSans 320 0 0 0 Tile_X0Y0_W1END[0]
port 208 nsew signal input
flabel metal3 s 21424 43388 21504 43468 0 FreeSans 320 0 0 0 Tile_X0Y0_W1END[1]
port 209 nsew signal input
flabel metal3 s 21424 43724 21504 43804 0 FreeSans 320 0 0 0 Tile_X0Y0_W1END[2]
port 210 nsew signal input
flabel metal3 s 21424 44060 21504 44140 0 FreeSans 320 0 0 0 Tile_X0Y0_W1END[3]
port 211 nsew signal input
flabel metal3 s 21424 47084 21504 47164 0 FreeSans 320 0 0 0 Tile_X0Y0_W2END[0]
port 212 nsew signal input
flabel metal3 s 21424 47420 21504 47500 0 FreeSans 320 0 0 0 Tile_X0Y0_W2END[1]
port 213 nsew signal input
flabel metal3 s 21424 47756 21504 47836 0 FreeSans 320 0 0 0 Tile_X0Y0_W2END[2]
port 214 nsew signal input
flabel metal3 s 21424 48092 21504 48172 0 FreeSans 320 0 0 0 Tile_X0Y0_W2END[3]
port 215 nsew signal input
flabel metal3 s 21424 48428 21504 48508 0 FreeSans 320 0 0 0 Tile_X0Y0_W2END[4]
port 216 nsew signal input
flabel metal3 s 21424 48764 21504 48844 0 FreeSans 320 0 0 0 Tile_X0Y0_W2END[5]
port 217 nsew signal input
flabel metal3 s 21424 49100 21504 49180 0 FreeSans 320 0 0 0 Tile_X0Y0_W2END[6]
port 218 nsew signal input
flabel metal3 s 21424 49436 21504 49516 0 FreeSans 320 0 0 0 Tile_X0Y0_W2END[7]
port 219 nsew signal input
flabel metal3 s 21424 44396 21504 44476 0 FreeSans 320 0 0 0 Tile_X0Y0_W2MID[0]
port 220 nsew signal input
flabel metal3 s 21424 44732 21504 44812 0 FreeSans 320 0 0 0 Tile_X0Y0_W2MID[1]
port 221 nsew signal input
flabel metal3 s 21424 45068 21504 45148 0 FreeSans 320 0 0 0 Tile_X0Y0_W2MID[2]
port 222 nsew signal input
flabel metal3 s 21424 45404 21504 45484 0 FreeSans 320 0 0 0 Tile_X0Y0_W2MID[3]
port 223 nsew signal input
flabel metal3 s 21424 45740 21504 45820 0 FreeSans 320 0 0 0 Tile_X0Y0_W2MID[4]
port 224 nsew signal input
flabel metal3 s 21424 46076 21504 46156 0 FreeSans 320 0 0 0 Tile_X0Y0_W2MID[5]
port 225 nsew signal input
flabel metal3 s 21424 46412 21504 46492 0 FreeSans 320 0 0 0 Tile_X0Y0_W2MID[6]
port 226 nsew signal input
flabel metal3 s 21424 46748 21504 46828 0 FreeSans 320 0 0 0 Tile_X0Y0_W2MID[7]
port 227 nsew signal input
flabel metal3 s 21424 55148 21504 55228 0 FreeSans 320 0 0 0 Tile_X0Y0_W6END[0]
port 228 nsew signal input
flabel metal3 s 21424 58508 21504 58588 0 FreeSans 320 0 0 0 Tile_X0Y0_W6END[10]
port 229 nsew signal input
flabel metal3 s 21424 58844 21504 58924 0 FreeSans 320 0 0 0 Tile_X0Y0_W6END[11]
port 230 nsew signal input
flabel metal3 s 21424 55484 21504 55564 0 FreeSans 320 0 0 0 Tile_X0Y0_W6END[1]
port 231 nsew signal input
flabel metal3 s 21424 55820 21504 55900 0 FreeSans 320 0 0 0 Tile_X0Y0_W6END[2]
port 232 nsew signal input
flabel metal3 s 21424 56156 21504 56236 0 FreeSans 320 0 0 0 Tile_X0Y0_W6END[3]
port 233 nsew signal input
flabel metal3 s 21424 56492 21504 56572 0 FreeSans 320 0 0 0 Tile_X0Y0_W6END[4]
port 234 nsew signal input
flabel metal3 s 21424 56828 21504 56908 0 FreeSans 320 0 0 0 Tile_X0Y0_W6END[5]
port 235 nsew signal input
flabel metal3 s 21424 57164 21504 57244 0 FreeSans 320 0 0 0 Tile_X0Y0_W6END[6]
port 236 nsew signal input
flabel metal3 s 21424 57500 21504 57580 0 FreeSans 320 0 0 0 Tile_X0Y0_W6END[7]
port 237 nsew signal input
flabel metal3 s 21424 57836 21504 57916 0 FreeSans 320 0 0 0 Tile_X0Y0_W6END[8]
port 238 nsew signal input
flabel metal3 s 21424 58172 21504 58252 0 FreeSans 320 0 0 0 Tile_X0Y0_W6END[9]
port 239 nsew signal input
flabel metal3 s 21424 49772 21504 49852 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[0]
port 240 nsew signal input
flabel metal3 s 21424 53132 21504 53212 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[10]
port 241 nsew signal input
flabel metal3 s 21424 53468 21504 53548 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[11]
port 242 nsew signal input
flabel metal3 s 21424 53804 21504 53884 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[12]
port 243 nsew signal input
flabel metal3 s 21424 54140 21504 54220 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[13]
port 244 nsew signal input
flabel metal3 s 21424 54476 21504 54556 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[14]
port 245 nsew signal input
flabel metal3 s 21424 54812 21504 54892 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[15]
port 246 nsew signal input
flabel metal3 s 21424 50108 21504 50188 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[1]
port 247 nsew signal input
flabel metal3 s 21424 50444 21504 50524 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[2]
port 248 nsew signal input
flabel metal3 s 21424 50780 21504 50860 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[3]
port 249 nsew signal input
flabel metal3 s 21424 51116 21504 51196 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[4]
port 250 nsew signal input
flabel metal3 s 21424 51452 21504 51532 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[5]
port 251 nsew signal input
flabel metal3 s 21424 51788 21504 51868 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[6]
port 252 nsew signal input
flabel metal3 s 21424 52124 21504 52204 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[7]
port 253 nsew signal input
flabel metal3 s 21424 52460 21504 52540 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[8]
port 254 nsew signal input
flabel metal3 s 21424 52796 21504 52876 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4END[9]
port 255 nsew signal input
flabel metal3 s 21424 16172 21504 16252 0 FreeSans 320 0 0 0 Tile_X0Y1_E1BEG[0]
port 256 nsew signal output
flabel metal3 s 21424 16508 21504 16588 0 FreeSans 320 0 0 0 Tile_X0Y1_E1BEG[1]
port 257 nsew signal output
flabel metal3 s 21424 16844 21504 16924 0 FreeSans 320 0 0 0 Tile_X0Y1_E1BEG[2]
port 258 nsew signal output
flabel metal3 s 21424 17180 21504 17260 0 FreeSans 320 0 0 0 Tile_X0Y1_E1BEG[3]
port 259 nsew signal output
flabel metal3 s 21424 17516 21504 17596 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEG[0]
port 260 nsew signal output
flabel metal3 s 21424 17852 21504 17932 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEG[1]
port 261 nsew signal output
flabel metal3 s 21424 18188 21504 18268 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEG[2]
port 262 nsew signal output
flabel metal3 s 21424 18524 21504 18604 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEG[3]
port 263 nsew signal output
flabel metal3 s 21424 18860 21504 18940 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEG[4]
port 264 nsew signal output
flabel metal3 s 21424 19196 21504 19276 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEG[5]
port 265 nsew signal output
flabel metal3 s 21424 19532 21504 19612 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEG[6]
port 266 nsew signal output
flabel metal3 s 21424 19868 21504 19948 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEG[7]
port 267 nsew signal output
flabel metal3 s 21424 20204 21504 20284 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEGb[0]
port 268 nsew signal output
flabel metal3 s 21424 20540 21504 20620 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEGb[1]
port 269 nsew signal output
flabel metal3 s 21424 20876 21504 20956 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEGb[2]
port 270 nsew signal output
flabel metal3 s 21424 21212 21504 21292 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEGb[3]
port 271 nsew signal output
flabel metal3 s 21424 21548 21504 21628 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEGb[4]
port 272 nsew signal output
flabel metal3 s 21424 21884 21504 21964 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEGb[5]
port 273 nsew signal output
flabel metal3 s 21424 22220 21504 22300 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEGb[6]
port 274 nsew signal output
flabel metal3 s 21424 22556 21504 22636 0 FreeSans 320 0 0 0 Tile_X0Y1_E2BEGb[7]
port 275 nsew signal output
flabel metal3 s 21424 28268 21504 28348 0 FreeSans 320 0 0 0 Tile_X0Y1_E6BEG[0]
port 276 nsew signal output
flabel metal3 s 21424 31628 21504 31708 0 FreeSans 320 0 0 0 Tile_X0Y1_E6BEG[10]
port 277 nsew signal output
flabel metal3 s 21424 31964 21504 32044 0 FreeSans 320 0 0 0 Tile_X0Y1_E6BEG[11]
port 278 nsew signal output
flabel metal3 s 21424 28604 21504 28684 0 FreeSans 320 0 0 0 Tile_X0Y1_E6BEG[1]
port 279 nsew signal output
flabel metal3 s 21424 28940 21504 29020 0 FreeSans 320 0 0 0 Tile_X0Y1_E6BEG[2]
port 280 nsew signal output
flabel metal3 s 21424 29276 21504 29356 0 FreeSans 320 0 0 0 Tile_X0Y1_E6BEG[3]
port 281 nsew signal output
flabel metal3 s 21424 29612 21504 29692 0 FreeSans 320 0 0 0 Tile_X0Y1_E6BEG[4]
port 282 nsew signal output
flabel metal3 s 21424 29948 21504 30028 0 FreeSans 320 0 0 0 Tile_X0Y1_E6BEG[5]
port 283 nsew signal output
flabel metal3 s 21424 30284 21504 30364 0 FreeSans 320 0 0 0 Tile_X0Y1_E6BEG[6]
port 284 nsew signal output
flabel metal3 s 21424 30620 21504 30700 0 FreeSans 320 0 0 0 Tile_X0Y1_E6BEG[7]
port 285 nsew signal output
flabel metal3 s 21424 30956 21504 31036 0 FreeSans 320 0 0 0 Tile_X0Y1_E6BEG[8]
port 286 nsew signal output
flabel metal3 s 21424 31292 21504 31372 0 FreeSans 320 0 0 0 Tile_X0Y1_E6BEG[9]
port 287 nsew signal output
flabel metal3 s 21424 22892 21504 22972 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[0]
port 288 nsew signal output
flabel metal3 s 21424 26252 21504 26332 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[10]
port 289 nsew signal output
flabel metal3 s 21424 26588 21504 26668 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[11]
port 290 nsew signal output
flabel metal3 s 21424 26924 21504 27004 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[12]
port 291 nsew signal output
flabel metal3 s 21424 27260 21504 27340 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[13]
port 292 nsew signal output
flabel metal3 s 21424 27596 21504 27676 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[14]
port 293 nsew signal output
flabel metal3 s 21424 27932 21504 28012 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[15]
port 294 nsew signal output
flabel metal3 s 21424 23228 21504 23308 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[1]
port 295 nsew signal output
flabel metal3 s 21424 23564 21504 23644 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[2]
port 296 nsew signal output
flabel metal3 s 21424 23900 21504 23980 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[3]
port 297 nsew signal output
flabel metal3 s 21424 24236 21504 24316 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[4]
port 298 nsew signal output
flabel metal3 s 21424 24572 21504 24652 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[5]
port 299 nsew signal output
flabel metal3 s 21424 24908 21504 24988 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[6]
port 300 nsew signal output
flabel metal3 s 21424 25244 21504 25324 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[7]
port 301 nsew signal output
flabel metal3 s 21424 25580 21504 25660 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[8]
port 302 nsew signal output
flabel metal3 s 21424 25916 21504 25996 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4BEG[9]
port 303 nsew signal output
flabel metal3 s 0 57668 80 57748 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[0]
port 304 nsew signal input
flabel metal3 s 0 64388 80 64468 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[10]
port 305 nsew signal input
flabel metal3 s 0 65060 80 65140 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[11]
port 306 nsew signal input
flabel metal3 s 0 65732 80 65812 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[12]
port 307 nsew signal input
flabel metal3 s 0 66404 80 66484 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[13]
port 308 nsew signal input
flabel metal3 s 0 67076 80 67156 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[14]
port 309 nsew signal input
flabel metal3 s 0 67748 80 67828 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[15]
port 310 nsew signal input
flabel metal3 s 0 68420 80 68500 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[16]
port 311 nsew signal input
flabel metal3 s 0 69092 80 69172 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[17]
port 312 nsew signal input
flabel metal3 s 0 69764 80 69844 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[18]
port 313 nsew signal input
flabel metal3 s 0 70436 80 70516 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[19]
port 314 nsew signal input
flabel metal3 s 0 58340 80 58420 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[1]
port 315 nsew signal input
flabel metal3 s 0 71108 80 71188 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[20]
port 316 nsew signal input
flabel metal3 s 0 71780 80 71860 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[21]
port 317 nsew signal input
flabel metal3 s 0 72452 80 72532 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[22]
port 318 nsew signal input
flabel metal3 s 0 73124 80 73204 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[23]
port 319 nsew signal input
flabel metal3 s 0 73796 80 73876 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[24]
port 320 nsew signal input
flabel metal3 s 0 74468 80 74548 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[25]
port 321 nsew signal input
flabel metal3 s 0 75140 80 75220 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[26]
port 322 nsew signal input
flabel metal3 s 0 75812 80 75892 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[27]
port 323 nsew signal input
flabel metal3 s 0 76484 80 76564 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[28]
port 324 nsew signal input
flabel metal3 s 0 77156 80 77236 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[29]
port 325 nsew signal input
flabel metal3 s 0 59012 80 59092 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[2]
port 326 nsew signal input
flabel metal3 s 0 77828 80 77908 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[30]
port 327 nsew signal input
flabel metal3 s 0 78500 80 78580 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[31]
port 328 nsew signal input
flabel metal3 s 0 59684 80 59764 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[3]
port 329 nsew signal input
flabel metal3 s 0 60356 80 60436 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[4]
port 330 nsew signal input
flabel metal3 s 0 61028 80 61108 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[5]
port 331 nsew signal input
flabel metal3 s 0 61700 80 61780 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[6]
port 332 nsew signal input
flabel metal3 s 0 62372 80 62452 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[7]
port 333 nsew signal input
flabel metal3 s 0 63044 80 63124 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[8]
port 334 nsew signal input
flabel metal3 s 0 63716 80 63796 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[9]
port 335 nsew signal input
flabel metal3 s 21424 32300 21504 32380 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[0]
port 336 nsew signal output
flabel metal3 s 21424 35660 21504 35740 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[10]
port 337 nsew signal output
flabel metal3 s 21424 35996 21504 36076 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[11]
port 338 nsew signal output
flabel metal3 s 21424 36332 21504 36412 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[12]
port 339 nsew signal output
flabel metal3 s 21424 36668 21504 36748 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[13]
port 340 nsew signal output
flabel metal3 s 21424 37004 21504 37084 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[14]
port 341 nsew signal output
flabel metal3 s 21424 37340 21504 37420 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[15]
port 342 nsew signal output
flabel metal3 s 21424 37676 21504 37756 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[16]
port 343 nsew signal output
flabel metal3 s 21424 38012 21504 38092 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[17]
port 344 nsew signal output
flabel metal3 s 21424 38348 21504 38428 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[18]
port 345 nsew signal output
flabel metal3 s 21424 38684 21504 38764 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[19]
port 346 nsew signal output
flabel metal3 s 21424 32636 21504 32716 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[1]
port 347 nsew signal output
flabel metal3 s 21424 39020 21504 39100 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[20]
port 348 nsew signal output
flabel metal3 s 21424 39356 21504 39436 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[21]
port 349 nsew signal output
flabel metal3 s 21424 39692 21504 39772 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[22]
port 350 nsew signal output
flabel metal3 s 21424 40028 21504 40108 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[23]
port 351 nsew signal output
flabel metal3 s 21424 40364 21504 40444 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[24]
port 352 nsew signal output
flabel metal3 s 21424 40700 21504 40780 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[25]
port 353 nsew signal output
flabel metal3 s 21424 41036 21504 41116 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[26]
port 354 nsew signal output
flabel metal3 s 21424 41372 21504 41452 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[27]
port 355 nsew signal output
flabel metal3 s 21424 41708 21504 41788 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[28]
port 356 nsew signal output
flabel metal3 s 21424 42044 21504 42124 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[29]
port 357 nsew signal output
flabel metal3 s 21424 32972 21504 33052 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[2]
port 358 nsew signal output
flabel metal3 s 21424 42380 21504 42460 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[30]
port 359 nsew signal output
flabel metal3 s 21424 42716 21504 42796 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[31]
port 360 nsew signal output
flabel metal3 s 21424 33308 21504 33388 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[3]
port 361 nsew signal output
flabel metal3 s 21424 33644 21504 33724 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[4]
port 362 nsew signal output
flabel metal3 s 21424 33980 21504 34060 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[5]
port 363 nsew signal output
flabel metal3 s 21424 34316 21504 34396 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[6]
port 364 nsew signal output
flabel metal3 s 21424 34652 21504 34732 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[7]
port 365 nsew signal output
flabel metal3 s 21424 34988 21504 35068 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[8]
port 366 nsew signal output
flabel metal3 s 21424 35324 21504 35404 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[9]
port 367 nsew signal output
flabel metal2 s 15800 0 15880 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[0]
port 368 nsew signal input
flabel metal2 s 17720 0 17800 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[10]
port 369 nsew signal input
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[11]
port 370 nsew signal input
flabel metal2 s 18104 0 18184 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[12]
port 371 nsew signal input
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[13]
port 372 nsew signal input
flabel metal2 s 18488 0 18568 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[14]
port 373 nsew signal input
flabel metal2 s 18680 0 18760 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[15]
port 374 nsew signal input
flabel metal2 s 18872 0 18952 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[16]
port 375 nsew signal input
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[17]
port 376 nsew signal input
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[18]
port 377 nsew signal input
flabel metal2 s 19448 0 19528 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[19]
port 378 nsew signal input
flabel metal2 s 15992 0 16072 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[1]
port 379 nsew signal input
flabel metal2 s 16184 0 16264 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[2]
port 380 nsew signal input
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[3]
port 381 nsew signal input
flabel metal2 s 16568 0 16648 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[4]
port 382 nsew signal input
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[5]
port 383 nsew signal input
flabel metal2 s 16952 0 17032 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[6]
port 384 nsew signal input
flabel metal2 s 17144 0 17224 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[7]
port 385 nsew signal input
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[8]
port 386 nsew signal input
flabel metal2 s 17528 0 17608 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[9]
port 387 nsew signal input
flabel metal2 s 1784 0 1864 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[0]
port 388 nsew signal input
flabel metal2 s 1976 0 2056 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[1]
port 389 nsew signal input
flabel metal2 s 2168 0 2248 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[2]
port 390 nsew signal input
flabel metal2 s 2360 0 2440 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[3]
port 391 nsew signal input
flabel metal2 s 4088 0 4168 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[0]
port 392 nsew signal input
flabel metal2 s 4280 0 4360 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[1]
port 393 nsew signal input
flabel metal2 s 4472 0 4552 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[2]
port 394 nsew signal input
flabel metal2 s 4664 0 4744 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[3]
port 395 nsew signal input
flabel metal2 s 4856 0 4936 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[4]
port 396 nsew signal input
flabel metal2 s 5048 0 5128 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[5]
port 397 nsew signal input
flabel metal2 s 5240 0 5320 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[6]
port 398 nsew signal input
flabel metal2 s 5432 0 5512 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[7]
port 399 nsew signal input
flabel metal2 s 2552 0 2632 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[0]
port 400 nsew signal input
flabel metal2 s 2744 0 2824 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[1]
port 401 nsew signal input
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[2]
port 402 nsew signal input
flabel metal2 s 3128 0 3208 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[3]
port 403 nsew signal input
flabel metal2 s 3320 0 3400 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[4]
port 404 nsew signal input
flabel metal2 s 3512 0 3592 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[5]
port 405 nsew signal input
flabel metal2 s 3704 0 3784 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[6]
port 406 nsew signal input
flabel metal2 s 3896 0 3976 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[7]
port 407 nsew signal input
flabel metal2 s 5624 0 5704 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[0]
port 408 nsew signal input
flabel metal2 s 7544 0 7624 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[10]
port 409 nsew signal input
flabel metal2 s 7736 0 7816 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[11]
port 410 nsew signal input
flabel metal2 s 7928 0 8008 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[12]
port 411 nsew signal input
flabel metal2 s 8120 0 8200 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[13]
port 412 nsew signal input
flabel metal2 s 8312 0 8392 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[14]
port 413 nsew signal input
flabel metal2 s 8504 0 8584 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[15]
port 414 nsew signal input
flabel metal2 s 5816 0 5896 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[1]
port 415 nsew signal input
flabel metal2 s 6008 0 6088 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[2]
port 416 nsew signal input
flabel metal2 s 6200 0 6280 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[3]
port 417 nsew signal input
flabel metal2 s 6392 0 6472 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[4]
port 418 nsew signal input
flabel metal2 s 6584 0 6664 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[5]
port 419 nsew signal input
flabel metal2 s 6776 0 6856 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[6]
port 420 nsew signal input
flabel metal2 s 6968 0 7048 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[7]
port 421 nsew signal input
flabel metal2 s 7160 0 7240 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[8]
port 422 nsew signal input
flabel metal2 s 7352 0 7432 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[9]
port 423 nsew signal input
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[0]
port 424 nsew signal output
flabel metal2 s 8888 0 8968 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[1]
port 425 nsew signal output
flabel metal2 s 9080 0 9160 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[2]
port 426 nsew signal output
flabel metal2 s 9272 0 9352 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[3]
port 427 nsew signal output
flabel metal2 s 9464 0 9544 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[0]
port 428 nsew signal output
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[1]
port 429 nsew signal output
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[2]
port 430 nsew signal output
flabel metal2 s 10040 0 10120 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[3]
port 431 nsew signal output
flabel metal2 s 10232 0 10312 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[4]
port 432 nsew signal output
flabel metal2 s 10424 0 10504 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[5]
port 433 nsew signal output
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[6]
port 434 nsew signal output
flabel metal2 s 10808 0 10888 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[7]
port 435 nsew signal output
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[0]
port 436 nsew signal output
flabel metal2 s 11192 0 11272 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[1]
port 437 nsew signal output
flabel metal2 s 11384 0 11464 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[2]
port 438 nsew signal output
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[3]
port 439 nsew signal output
flabel metal2 s 11768 0 11848 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[4]
port 440 nsew signal output
flabel metal2 s 11960 0 12040 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[5]
port 441 nsew signal output
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[6]
port 442 nsew signal output
flabel metal2 s 12344 0 12424 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[7]
port 443 nsew signal output
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[0]
port 444 nsew signal output
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[10]
port 445 nsew signal output
flabel metal2 s 14648 0 14728 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[11]
port 446 nsew signal output
flabel metal2 s 14840 0 14920 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[12]
port 447 nsew signal output
flabel metal2 s 15032 0 15112 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[13]
port 448 nsew signal output
flabel metal2 s 15224 0 15304 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[14]
port 449 nsew signal output
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[15]
port 450 nsew signal output
flabel metal2 s 12728 0 12808 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[1]
port 451 nsew signal output
flabel metal2 s 12920 0 13000 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[2]
port 452 nsew signal output
flabel metal2 s 13112 0 13192 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[3]
port 453 nsew signal output
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[4]
port 454 nsew signal output
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[5]
port 455 nsew signal output
flabel metal2 s 13688 0 13768 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[6]
port 456 nsew signal output
flabel metal2 s 13880 0 13960 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[7]
port 457 nsew signal output
flabel metal2 s 14072 0 14152 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[8]
port 458 nsew signal output
flabel metal2 s 14264 0 14344 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[9]
port 459 nsew signal output
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 Tile_X0Y1_UserCLK
port 460 nsew signal input
flabel metal3 s 21424 44 21504 124 0 FreeSans 320 0 0 0 Tile_X0Y1_W1END[0]
port 461 nsew signal input
flabel metal3 s 21424 380 21504 460 0 FreeSans 320 0 0 0 Tile_X0Y1_W1END[1]
port 462 nsew signal input
flabel metal3 s 21424 716 21504 796 0 FreeSans 320 0 0 0 Tile_X0Y1_W1END[2]
port 463 nsew signal input
flabel metal3 s 21424 1052 21504 1132 0 FreeSans 320 0 0 0 Tile_X0Y1_W1END[3]
port 464 nsew signal input
flabel metal3 s 21424 4076 21504 4156 0 FreeSans 320 0 0 0 Tile_X0Y1_W2END[0]
port 465 nsew signal input
flabel metal3 s 21424 4412 21504 4492 0 FreeSans 320 0 0 0 Tile_X0Y1_W2END[1]
port 466 nsew signal input
flabel metal3 s 21424 4748 21504 4828 0 FreeSans 320 0 0 0 Tile_X0Y1_W2END[2]
port 467 nsew signal input
flabel metal3 s 21424 5084 21504 5164 0 FreeSans 320 0 0 0 Tile_X0Y1_W2END[3]
port 468 nsew signal input
flabel metal3 s 21424 5420 21504 5500 0 FreeSans 320 0 0 0 Tile_X0Y1_W2END[4]
port 469 nsew signal input
flabel metal3 s 21424 5756 21504 5836 0 FreeSans 320 0 0 0 Tile_X0Y1_W2END[5]
port 470 nsew signal input
flabel metal3 s 21424 6092 21504 6172 0 FreeSans 320 0 0 0 Tile_X0Y1_W2END[6]
port 471 nsew signal input
flabel metal3 s 21424 6428 21504 6508 0 FreeSans 320 0 0 0 Tile_X0Y1_W2END[7]
port 472 nsew signal input
flabel metal3 s 21424 1388 21504 1468 0 FreeSans 320 0 0 0 Tile_X0Y1_W2MID[0]
port 473 nsew signal input
flabel metal3 s 21424 1724 21504 1804 0 FreeSans 320 0 0 0 Tile_X0Y1_W2MID[1]
port 474 nsew signal input
flabel metal3 s 21424 2060 21504 2140 0 FreeSans 320 0 0 0 Tile_X0Y1_W2MID[2]
port 475 nsew signal input
flabel metal3 s 21424 2396 21504 2476 0 FreeSans 320 0 0 0 Tile_X0Y1_W2MID[3]
port 476 nsew signal input
flabel metal3 s 21424 2732 21504 2812 0 FreeSans 320 0 0 0 Tile_X0Y1_W2MID[4]
port 477 nsew signal input
flabel metal3 s 21424 3068 21504 3148 0 FreeSans 320 0 0 0 Tile_X0Y1_W2MID[5]
port 478 nsew signal input
flabel metal3 s 21424 3404 21504 3484 0 FreeSans 320 0 0 0 Tile_X0Y1_W2MID[6]
port 479 nsew signal input
flabel metal3 s 21424 3740 21504 3820 0 FreeSans 320 0 0 0 Tile_X0Y1_W2MID[7]
port 480 nsew signal input
flabel metal3 s 21424 12140 21504 12220 0 FreeSans 320 0 0 0 Tile_X0Y1_W6END[0]
port 481 nsew signal input
flabel metal3 s 21424 15500 21504 15580 0 FreeSans 320 0 0 0 Tile_X0Y1_W6END[10]
port 482 nsew signal input
flabel metal3 s 21424 15836 21504 15916 0 FreeSans 320 0 0 0 Tile_X0Y1_W6END[11]
port 483 nsew signal input
flabel metal3 s 21424 12476 21504 12556 0 FreeSans 320 0 0 0 Tile_X0Y1_W6END[1]
port 484 nsew signal input
flabel metal3 s 21424 12812 21504 12892 0 FreeSans 320 0 0 0 Tile_X0Y1_W6END[2]
port 485 nsew signal input
flabel metal3 s 21424 13148 21504 13228 0 FreeSans 320 0 0 0 Tile_X0Y1_W6END[3]
port 486 nsew signal input
flabel metal3 s 21424 13484 21504 13564 0 FreeSans 320 0 0 0 Tile_X0Y1_W6END[4]
port 487 nsew signal input
flabel metal3 s 21424 13820 21504 13900 0 FreeSans 320 0 0 0 Tile_X0Y1_W6END[5]
port 488 nsew signal input
flabel metal3 s 21424 14156 21504 14236 0 FreeSans 320 0 0 0 Tile_X0Y1_W6END[6]
port 489 nsew signal input
flabel metal3 s 21424 14492 21504 14572 0 FreeSans 320 0 0 0 Tile_X0Y1_W6END[7]
port 490 nsew signal input
flabel metal3 s 21424 14828 21504 14908 0 FreeSans 320 0 0 0 Tile_X0Y1_W6END[8]
port 491 nsew signal input
flabel metal3 s 21424 15164 21504 15244 0 FreeSans 320 0 0 0 Tile_X0Y1_W6END[9]
port 492 nsew signal input
flabel metal3 s 21424 6764 21504 6844 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[0]
port 493 nsew signal input
flabel metal3 s 21424 10124 21504 10204 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[10]
port 494 nsew signal input
flabel metal3 s 21424 10460 21504 10540 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[11]
port 495 nsew signal input
flabel metal3 s 21424 10796 21504 10876 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[12]
port 496 nsew signal input
flabel metal3 s 21424 11132 21504 11212 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[13]
port 497 nsew signal input
flabel metal3 s 21424 11468 21504 11548 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[14]
port 498 nsew signal input
flabel metal3 s 21424 11804 21504 11884 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[15]
port 499 nsew signal input
flabel metal3 s 21424 7100 21504 7180 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[1]
port 500 nsew signal input
flabel metal3 s 21424 7436 21504 7516 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[2]
port 501 nsew signal input
flabel metal3 s 21424 7772 21504 7852 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[3]
port 502 nsew signal input
flabel metal3 s 21424 8108 21504 8188 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[4]
port 503 nsew signal input
flabel metal3 s 21424 8444 21504 8524 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[5]
port 504 nsew signal input
flabel metal3 s 21424 8780 21504 8860 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[6]
port 505 nsew signal input
flabel metal3 s 21424 9116 21504 9196 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[7]
port 506 nsew signal input
flabel metal3 s 21424 9452 21504 9532 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[8]
port 507 nsew signal input
flabel metal3 s 21424 9788 21504 9868 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4END[9]
port 508 nsew signal input
flabel metal3 s 0 28772 80 28852 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT0
port 509 nsew signal output
flabel metal3 s 0 29444 80 29524 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT1
port 510 nsew signal output
flabel metal3 s 0 30116 80 30196 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT2
port 511 nsew signal output
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT3
port 512 nsew signal output
flabel metal3 s 0 31460 80 31540 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT4
port 513 nsew signal output
flabel metal3 s 0 32132 80 32212 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT5
port 514 nsew signal output
flabel metal3 s 0 32804 80 32884 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT6
port 515 nsew signal output
flabel metal3 s 0 33476 80 33556 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT7
port 516 nsew signal output
flabel metal3 s 0 18020 80 18100 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT0
port 517 nsew signal input
flabel metal3 s 0 18692 80 18772 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT1
port 518 nsew signal input
flabel metal3 s 0 19364 80 19444 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT2
port 519 nsew signal input
flabel metal3 s 0 20036 80 20116 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT3
port 520 nsew signal input
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT4
port 521 nsew signal input
flabel metal3 s 0 21380 80 21460 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT5
port 522 nsew signal input
flabel metal3 s 0 22052 80 22132 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT6
port 523 nsew signal input
flabel metal3 s 0 22724 80 22804 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT7
port 524 nsew signal input
flabel metal3 s 0 12644 80 12724 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT0
port 525 nsew signal input
flabel metal3 s 0 13316 80 13396 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT1
port 526 nsew signal input
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT2
port 527 nsew signal input
flabel metal3 s 0 14660 80 14740 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT3
port 528 nsew signal input
flabel metal3 s 0 15332 80 15412 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT4
port 529 nsew signal input
flabel metal3 s 0 16004 80 16084 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT5
port 530 nsew signal input
flabel metal3 s 0 16676 80 16756 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT6
port 531 nsew signal input
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT7
port 532 nsew signal input
flabel metal3 s 0 23396 80 23476 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT0
port 533 nsew signal output
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT1
port 534 nsew signal output
flabel metal3 s 0 24740 80 24820 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT2
port 535 nsew signal output
flabel metal3 s 0 25412 80 25492 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT3
port 536 nsew signal output
flabel metal3 s 0 26084 80 26164 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT4
port 537 nsew signal output
flabel metal3 s 0 26756 80 26836 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT5
port 538 nsew signal output
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT6
port 539 nsew signal output
flabel metal3 s 0 28100 80 28180 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT7
port 540 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT0
port 541 nsew signal input
flabel metal3 s 0 7940 80 8020 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT1
port 542 nsew signal input
flabel metal3 s 0 8612 80 8692 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT2
port 543 nsew signal input
flabel metal3 s 0 9284 80 9364 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT3
port 544 nsew signal input
flabel metal3 s 0 9956 80 10036 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT4
port 545 nsew signal input
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT5
port 546 nsew signal input
flabel metal3 s 0 11300 80 11380 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT6
port 547 nsew signal input
flabel metal3 s 0 11972 80 12052 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT7
port 548 nsew signal input
flabel metal6 s 4892 0 5332 86016 0 FreeSans 2624 90 0 0 VGND
port 549 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 549 nsew ground bidirectional
flabel metal6 s 4892 85688 5332 86016 0 FreeSans 2624 0 0 0 VGND
port 549 nsew ground bidirectional
flabel metal6 s 20012 0 20452 86016 0 FreeSans 2624 90 0 0 VGND
port 549 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 549 nsew ground bidirectional
flabel metal6 s 20012 85688 20452 86016 0 FreeSans 2624 0 0 0 VGND
port 549 nsew ground bidirectional
flabel metal6 s 3652 0 4092 86016 0 FreeSans 2624 90 0 0 VPWR
port 550 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 550 nsew power bidirectional
flabel metal6 s 3652 85688 4092 86016 0 FreeSans 2624 0 0 0 VPWR
port 550 nsew power bidirectional
flabel metal6 s 18772 0 19212 86016 0 FreeSans 2624 90 0 0 VPWR
port 550 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 550 nsew power bidirectional
flabel metal6 s 18772 85688 19212 86016 0 FreeSans 2624 0 0 0 VPWR
port 550 nsew power bidirectional
rlabel metal1 10802 83916 10802 83916 0 VGND
rlabel metal1 10752 84672 10752 84672 0 VPWR
rlabel metal3 990 34860 990 34860 0 CLK_TT_PROJECT
rlabel metal2 2832 33852 2832 33852 0 ENA_TT_PROJECT
rlabel via2 78 35532 78 35532 0 RST_N_TT_PROJECT
rlabel metal2 19968 58968 19968 58968 0 Tile_X0Y0_E1BEG[0]
rlabel metal3 20706 59556 20706 59556 0 Tile_X0Y0_E1BEG[1]
rlabel metal3 20706 59892 20706 59892 0 Tile_X0Y0_E1BEG[2]
rlabel metal3 20850 60228 20850 60228 0 Tile_X0Y0_E1BEG[3]
rlabel metal3 21234 60564 21234 60564 0 Tile_X0Y0_E2BEG[0]
rlabel metal2 19536 58800 19536 58800 0 Tile_X0Y0_E2BEG[1]
rlabel metal3 21378 61236 21378 61236 0 Tile_X0Y0_E2BEG[2]
rlabel metal2 19200 61488 19200 61488 0 Tile_X0Y0_E2BEG[3]
rlabel metal2 19968 61824 19968 61824 0 Tile_X0Y0_E2BEG[4]
rlabel metal2 18768 61740 18768 61740 0 Tile_X0Y0_E2BEG[5]
rlabel metal3 20658 62580 20658 62580 0 Tile_X0Y0_E2BEG[6]
rlabel metal2 20400 62580 20400 62580 0 Tile_X0Y0_E2BEG[7]
rlabel metal3 20562 63252 20562 63252 0 Tile_X0Y0_E2BEGb[0]
rlabel metal2 19584 59388 19584 59388 0 Tile_X0Y0_E2BEGb[1]
rlabel metal2 19584 63840 19584 63840 0 Tile_X0Y0_E2BEGb[2]
rlabel metal3 20256 64344 20256 64344 0 Tile_X0Y0_E2BEGb[3]
rlabel metal2 19584 64512 19584 64512 0 Tile_X0Y0_E2BEGb[4]
rlabel metal2 19296 65058 19296 65058 0 Tile_X0Y0_E2BEGb[5]
rlabel metal2 20016 64848 20016 64848 0 Tile_X0Y0_E2BEGb[6]
rlabel metal2 19968 65436 19968 65436 0 Tile_X0Y0_E2BEGb[7]
rlabel metal2 19680 71736 19680 71736 0 Tile_X0Y0_E6BEG[0]
rlabel metal3 21138 74676 21138 74676 0 Tile_X0Y0_E6BEG[10]
rlabel metal3 20994 75012 20994 75012 0 Tile_X0Y0_E6BEG[11]
rlabel metal4 19968 71946 19968 71946 0 Tile_X0Y0_E6BEG[1]
rlabel metal3 21090 71988 21090 71988 0 Tile_X0Y0_E6BEG[2]
rlabel metal3 20562 72324 20562 72324 0 Tile_X0Y0_E6BEG[3]
rlabel metal3 20466 72660 20466 72660 0 Tile_X0Y0_E6BEG[4]
rlabel metal3 20514 72996 20514 72996 0 Tile_X0Y0_E6BEG[5]
rlabel metal3 20544 73206 20544 73206 0 Tile_X0Y0_E6BEG[6]
rlabel metal2 19200 73584 19200 73584 0 Tile_X0Y0_E6BEG[7]
rlabel metal4 19968 75390 19968 75390 0 Tile_X0Y0_E6BEG[8]
rlabel metal3 21090 74340 21090 74340 0 Tile_X0Y0_E6BEG[9]
rlabel metal3 20514 65940 20514 65940 0 Tile_X0Y0_EE4BEG[0]
rlabel metal3 20994 69300 20994 69300 0 Tile_X0Y0_EE4BEG[10]
rlabel metal2 20064 69846 20064 69846 0 Tile_X0Y0_EE4BEG[11]
rlabel metal2 17952 69636 17952 69636 0 Tile_X0Y0_EE4BEG[12]
rlabel metal3 21378 70308 21378 70308 0 Tile_X0Y0_EE4BEG[13]
rlabel metal2 20064 71106 20064 71106 0 Tile_X0Y0_EE4BEG[14]
rlabel metal3 21042 70980 21042 70980 0 Tile_X0Y0_EE4BEG[15]
rlabel metal3 20706 66276 20706 66276 0 Tile_X0Y0_EE4BEG[1]
rlabel metal2 19584 65352 19584 65352 0 Tile_X0Y0_EE4BEG[2]
rlabel metal2 19968 67200 19968 67200 0 Tile_X0Y0_EE4BEG[3]
rlabel metal3 21378 67284 21378 67284 0 Tile_X0Y0_EE4BEG[4]
rlabel metal2 19680 67914 19680 67914 0 Tile_X0Y0_EE4BEG[5]
rlabel metal3 21042 67956 21042 67956 0 Tile_X0Y0_EE4BEG[6]
rlabel metal2 20064 68418 20064 68418 0 Tile_X0Y0_EE4BEG[7]
rlabel metal3 21138 68628 21138 68628 0 Tile_X0Y0_EE4BEG[8]
rlabel via2 21426 68964 21426 68964 0 Tile_X0Y0_EE4BEG[9]
rlabel metal2 13728 49812 13728 49812 0 Tile_X0Y0_FrameData[0]
rlabel metal2 2208 53592 2208 53592 0 Tile_X0Y0_FrameData[10]
rlabel metal2 18432 55734 18432 55734 0 Tile_X0Y0_FrameData[11]
rlabel metal2 1536 69216 1536 69216 0 Tile_X0Y0_FrameData[12]
rlabel metal2 14880 54600 14880 54600 0 Tile_X0Y0_FrameData[13]
rlabel metal3 1086 45612 1086 45612 0 Tile_X0Y0_FrameData[14]
rlabel metal2 15024 72996 15024 72996 0 Tile_X0Y0_FrameData[15]
rlabel metal2 1536 54012 1536 54012 0 Tile_X0Y0_FrameData[16]
rlabel metal3 1038 47628 1038 47628 0 Tile_X0Y0_FrameData[17]
rlabel metal3 1776 66948 1776 66948 0 Tile_X0Y0_FrameData[18]
rlabel metal2 1344 48888 1344 48888 0 Tile_X0Y0_FrameData[19]
rlabel metal2 2016 44478 2016 44478 0 Tile_X0Y0_FrameData[1]
rlabel metal2 1344 72240 1344 72240 0 Tile_X0Y0_FrameData[20]
rlabel metal3 894 50316 894 50316 0 Tile_X0Y0_FrameData[21]
rlabel metal2 12480 53382 12480 53382 0 Tile_X0Y0_FrameData[22]
rlabel metal3 40 51996 40 51996 0 Tile_X0Y0_FrameData[23]
rlabel metal3 126 52332 126 52332 0 Tile_X0Y0_FrameData[24]
rlabel metal3 16464 82824 16464 82824 0 Tile_X0Y0_FrameData[25]
rlabel metal2 1296 54264 1296 54264 0 Tile_X0Y0_FrameData[26]
rlabel metal3 16608 54852 16608 54852 0 Tile_X0Y0_FrameData[27]
rlabel metal2 1536 72114 1536 72114 0 Tile_X0Y0_FrameData[28]
rlabel metal2 1344 56364 1344 56364 0 Tile_X0Y0_FrameData[29]
rlabel metal2 1296 53340 1296 53340 0 Tile_X0Y0_FrameData[2]
rlabel metal2 19632 83580 19632 83580 0 Tile_X0Y0_FrameData[30]
rlabel metal2 1440 46284 1440 46284 0 Tile_X0Y0_FrameData[31]
rlabel metal3 1728 51828 1728 51828 0 Tile_X0Y0_FrameData[3]
rlabel metal2 1440 52542 1440 52542 0 Tile_X0Y0_FrameData[4]
rlabel metal3 126 39564 126 39564 0 Tile_X0Y0_FrameData[5]
rlabel metal4 11520 49224 11520 49224 0 Tile_X0Y0_FrameData[6]
rlabel metal2 15552 50232 15552 50232 0 Tile_X0Y0_FrameData[7]
rlabel metal3 480 41622 480 41622 0 Tile_X0Y0_FrameData[8]
rlabel metal2 18144 68880 18144 68880 0 Tile_X0Y0_FrameData[9]
rlabel metal3 21042 75348 21042 75348 0 Tile_X0Y0_FrameData_O[0]
rlabel metal2 19680 79128 19680 79128 0 Tile_X0Y0_FrameData_O[10]
rlabel metal2 18768 78456 18768 78456 0 Tile_X0Y0_FrameData_O[11]
rlabel metal3 20544 79422 20544 79422 0 Tile_X0Y0_FrameData_O[12]
rlabel metal2 19968 79632 19968 79632 0 Tile_X0Y0_FrameData_O[13]
rlabel metal2 19584 80178 19584 80178 0 Tile_X0Y0_FrameData_O[14]
rlabel metal2 16704 80178 16704 80178 0 Tile_X0Y0_FrameData_O[15]
rlabel metal2 19248 79968 19248 79968 0 Tile_X0Y0_FrameData_O[16]
rlabel metal2 18912 80724 18912 80724 0 Tile_X0Y0_FrameData_O[17]
rlabel metal2 19968 80892 19968 80892 0 Tile_X0Y0_FrameData_O[18]
rlabel metal2 19584 81606 19584 81606 0 Tile_X0Y0_FrameData_O[19]
rlabel metal2 20064 75894 20064 75894 0 Tile_X0Y0_FrameData_O[1]
rlabel via3 21426 82068 21426 82068 0 Tile_X0Y0_FrameData_O[20]
rlabel metal3 20112 82320 20112 82320 0 Tile_X0Y0_FrameData_O[21]
rlabel via2 21426 82740 21426 82740 0 Tile_X0Y0_FrameData_O[22]
rlabel metal2 15744 82656 15744 82656 0 Tile_X0Y0_FrameData_O[23]
rlabel metal2 19632 82992 19632 82992 0 Tile_X0Y0_FrameData_O[24]
rlabel metal2 19248 82992 19248 82992 0 Tile_X0Y0_FrameData_O[25]
rlabel metal3 21042 84084 21042 84084 0 Tile_X0Y0_FrameData_O[26]
rlabel metal2 20400 67116 20400 67116 0 Tile_X0Y0_FrameData_O[27]
rlabel metal3 20658 84756 20658 84756 0 Tile_X0Y0_FrameData_O[28]
rlabel metal3 20658 85092 20658 85092 0 Tile_X0Y0_FrameData_O[29]
rlabel metal3 20898 76020 20898 76020 0 Tile_X0Y0_FrameData_O[2]
rlabel metal2 19584 84588 19584 84588 0 Tile_X0Y0_FrameData_O[30]
rlabel metal2 19200 84126 19200 84126 0 Tile_X0Y0_FrameData_O[31]
rlabel metal3 20994 76356 20994 76356 0 Tile_X0Y0_FrameData_O[3]
rlabel metal2 18816 76608 18816 76608 0 Tile_X0Y0_FrameData_O[4]
rlabel metal2 20064 77238 20064 77238 0 Tile_X0Y0_FrameData_O[5]
rlabel metal2 15456 76776 15456 76776 0 Tile_X0Y0_FrameData_O[6]
rlabel metal3 20994 77700 20994 77700 0 Tile_X0Y0_FrameData_O[7]
rlabel metal3 21426 78036 21426 78036 0 Tile_X0Y0_FrameData_O[8]
rlabel metal3 20898 78372 20898 78372 0 Tile_X0Y0_FrameData_O[9]
rlabel metal2 15792 79968 15792 79968 0 Tile_X0Y0_FrameStrobe_O[0]
rlabel metal4 20928 28896 20928 28896 0 Tile_X0Y0_FrameStrobe_O[10]
rlabel metal2 17952 85524 17952 85524 0 Tile_X0Y0_FrameStrobe_O[11]
rlabel metal2 18144 85188 18144 85188 0 Tile_X0Y0_FrameStrobe_O[12]
rlabel metal2 18336 85230 18336 85230 0 Tile_X0Y0_FrameStrobe_O[13]
rlabel metal2 18528 85188 18528 85188 0 Tile_X0Y0_FrameStrobe_O[14]
rlabel metal2 18720 85230 18720 85230 0 Tile_X0Y0_FrameStrobe_O[15]
rlabel metal4 20688 28392 20688 28392 0 Tile_X0Y0_FrameStrobe_O[16]
rlabel via2 19104 85944 19104 85944 0 Tile_X0Y0_FrameStrobe_O[17]
rlabel via2 19296 85944 19296 85944 0 Tile_X0Y0_FrameStrobe_O[18]
rlabel metal2 19488 85188 19488 85188 0 Tile_X0Y0_FrameStrobe_O[19]
rlabel metal2 15984 79968 15984 79968 0 Tile_X0Y0_FrameStrobe_O[1]
rlabel metal3 16656 77700 16656 77700 0 Tile_X0Y0_FrameStrobe_O[2]
rlabel metal2 16704 77784 16704 77784 0 Tile_X0Y0_FrameStrobe_O[3]
rlabel metal3 16512 77448 16512 77448 0 Tile_X0Y0_FrameStrobe_O[4]
rlabel metal3 16656 62580 16656 62580 0 Tile_X0Y0_FrameStrobe_O[5]
rlabel metal2 16992 85776 16992 85776 0 Tile_X0Y0_FrameStrobe_O[6]
rlabel metal2 17184 85188 17184 85188 0 Tile_X0Y0_FrameStrobe_O[7]
rlabel metal2 17376 85230 17376 85230 0 Tile_X0Y0_FrameStrobe_O[8]
rlabel metal2 17568 85188 17568 85188 0 Tile_X0Y0_FrameStrobe_O[9]
rlabel metal2 1776 83748 1776 83748 0 Tile_X0Y0_N1BEG[0]
rlabel metal2 1968 83748 1968 83748 0 Tile_X0Y0_N1BEG[1]
rlabel metal2 2688 83286 2688 83286 0 Tile_X0Y0_N1BEG[2]
rlabel metal2 2352 83748 2352 83748 0 Tile_X0Y0_N1BEG[3]
rlabel metal2 2928 82992 2928 82992 0 Tile_X0Y0_N2BEG[0]
rlabel metal2 2736 83748 2736 83748 0 Tile_X0Y0_N2BEG[1]
rlabel metal2 3456 83286 3456 83286 0 Tile_X0Y0_N2BEG[2]
rlabel metal2 3120 83748 3120 83748 0 Tile_X0Y0_N2BEG[3]
rlabel metal2 4032 82992 4032 82992 0 Tile_X0Y0_N2BEG[4]
rlabel metal2 3504 83748 3504 83748 0 Tile_X0Y0_N2BEG[5]
rlabel metal3 3888 84420 3888 84420 0 Tile_X0Y0_N2BEG[6]
rlabel metal2 3840 84126 3840 84126 0 Tile_X0Y0_N2BEG[7]
rlabel metal2 4560 82992 4560 82992 0 Tile_X0Y0_N2BEGb[0]
rlabel metal2 4224 84210 4224 84210 0 Tile_X0Y0_N2BEGb[1]
rlabel metal2 4608 84210 4608 84210 0 Tile_X0Y0_N2BEGb[2]
rlabel metal2 4848 83748 4848 83748 0 Tile_X0Y0_N2BEGb[3]
rlabel metal2 5376 83916 5376 83916 0 Tile_X0Y0_N2BEGb[4]
rlabel metal2 5088 85314 5088 85314 0 Tile_X0Y0_N2BEGb[5]
rlabel metal2 5280 85272 5280 85272 0 Tile_X0Y0_N2BEGb[6]
rlabel metal2 5808 83748 5808 83748 0 Tile_X0Y0_N2BEGb[7]
rlabel metal5 3956 2100 3956 2100 0 Tile_X0Y0_N4BEG[0]
rlabel metal3 7104 83748 7104 83748 0 Tile_X0Y0_N4BEG[10]
rlabel metal2 13296 83748 13296 83748 0 Tile_X0Y0_N4BEG[11]
rlabel metal3 11472 83748 11472 83748 0 Tile_X0Y0_N4BEG[12]
rlabel metal2 7584 83874 7584 83874 0 Tile_X0Y0_N4BEG[13]
rlabel metal2 8352 84852 8352 84852 0 Tile_X0Y0_N4BEG[14]
rlabel metal2 18096 83748 18096 83748 0 Tile_X0Y0_N4BEG[15]
rlabel metal2 5856 85188 5856 85188 0 Tile_X0Y0_N4BEG[1]
rlabel metal2 6144 2142 6144 2142 0 Tile_X0Y0_N4BEG[2]
rlabel metal2 6240 85188 6240 85188 0 Tile_X0Y0_N4BEG[3]
rlabel metal2 6432 85776 6432 85776 0 Tile_X0Y0_N4BEG[4]
rlabel metal2 6624 85230 6624 85230 0 Tile_X0Y0_N4BEG[5]
rlabel metal5 7232 2100 7232 2100 0 Tile_X0Y0_N4BEG[6]
rlabel metal2 7680 2226 7680 2226 0 Tile_X0Y0_N4BEG[7]
rlabel metal2 15744 84798 15744 84798 0 Tile_X0Y0_N4BEG[8]
rlabel metal2 7200 84210 7200 84210 0 Tile_X0Y0_N4BEG[9]
rlabel metal2 8736 84936 8736 84936 0 Tile_X0Y0_S1END[0]
rlabel metal2 3744 61278 3744 61278 0 Tile_X0Y0_S1END[1]
rlabel metal2 3456 69090 3456 69090 0 Tile_X0Y0_S1END[2]
rlabel metal3 9456 83916 9456 83916 0 Tile_X0Y0_S1END[3]
rlabel metal2 11040 84138 11040 84138 0 Tile_X0Y0_S2END[0]
rlabel metal2 11232 84012 11232 84012 0 Tile_X0Y0_S2END[1]
rlabel metal2 11424 84894 11424 84894 0 Tile_X0Y0_S2END[2]
rlabel metal2 11616 83928 11616 83928 0 Tile_X0Y0_S2END[3]
rlabel metal2 11712 79296 11712 79296 0 Tile_X0Y0_S2END[4]
rlabel metal2 12000 84600 12000 84600 0 Tile_X0Y0_S2END[5]
rlabel metal2 12192 85188 12192 85188 0 Tile_X0Y0_S2END[6]
rlabel metal2 12384 84222 12384 84222 0 Tile_X0Y0_S2END[7]
rlabel metal3 10080 16380 10080 16380 0 Tile_X0Y0_S2MID[0]
rlabel metal2 8880 70644 8880 70644 0 Tile_X0Y0_S2MID[1]
rlabel via1 6521 18563 6521 18563 0 Tile_X0Y0_S2MID[2]
rlabel metal3 9264 84420 9264 84420 0 Tile_X0Y0_S2MID[3]
rlabel metal3 10896 41916 10896 41916 0 Tile_X0Y0_S2MID[4]
rlabel metal2 10464 84558 10464 84558 0 Tile_X0Y0_S2MID[5]
rlabel metal2 10656 85188 10656 85188 0 Tile_X0Y0_S2MID[6]
rlabel metal3 11184 38220 11184 38220 0 Tile_X0Y0_S2MID[7]
rlabel metal3 13776 71484 13776 71484 0 Tile_X0Y0_S4END[0]
rlabel metal2 14496 85440 14496 85440 0 Tile_X0Y0_S4END[10]
rlabel metal2 14688 85272 14688 85272 0 Tile_X0Y0_S4END[11]
rlabel metal2 14880 85230 14880 85230 0 Tile_X0Y0_S4END[12]
rlabel metal2 15072 85188 15072 85188 0 Tile_X0Y0_S4END[13]
rlabel metal2 15264 85188 15264 85188 0 Tile_X0Y0_S4END[14]
rlabel metal2 15456 85776 15456 85776 0 Tile_X0Y0_S4END[15]
rlabel metal2 12768 83970 12768 83970 0 Tile_X0Y0_S4END[1]
rlabel metal2 12960 83592 12960 83592 0 Tile_X0Y0_S4END[2]
rlabel metal2 14208 79170 14208 79170 0 Tile_X0Y0_S4END[3]
rlabel metal2 13344 85188 13344 85188 0 Tile_X0Y0_S4END[4]
rlabel metal2 13536 84810 13536 84810 0 Tile_X0Y0_S4END[5]
rlabel metal2 13728 85188 13728 85188 0 Tile_X0Y0_S4END[6]
rlabel metal2 13920 85188 13920 85188 0 Tile_X0Y0_S4END[7]
rlabel metal2 14112 85230 14112 85230 0 Tile_X0Y0_S4END[8]
rlabel metal2 14304 85188 14304 85188 0 Tile_X0Y0_S4END[9]
rlabel metal2 15600 83748 15600 83748 0 Tile_X0Y0_UserCLKo
rlabel metal2 18528 44436 18528 44436 0 Tile_X0Y0_W1END[0]
rlabel metal2 10272 46410 10272 46410 0 Tile_X0Y0_W1END[1]
rlabel metal2 9120 54054 9120 54054 0 Tile_X0Y0_W1END[2]
rlabel metal2 16320 51786 16320 51786 0 Tile_X0Y0_W1END[3]
rlabel metal2 19152 46704 19152 46704 0 Tile_X0Y0_W2END[0]
rlabel metal3 18882 47460 18882 47460 0 Tile_X0Y0_W2END[1]
rlabel metal2 10944 50064 10944 50064 0 Tile_X0Y0_W2END[2]
rlabel metal3 21378 48132 21378 48132 0 Tile_X0Y0_W2END[3]
rlabel metal3 21378 48468 21378 48468 0 Tile_X0Y0_W2END[4]
rlabel metal2 10080 49140 10080 49140 0 Tile_X0Y0_W2END[5]
rlabel metal3 20994 49140 20994 49140 0 Tile_X0Y0_W2END[6]
rlabel metal3 20802 49476 20802 49476 0 Tile_X0Y0_W2END[7]
rlabel metal2 18720 44352 18720 44352 0 Tile_X0Y0_W2MID[0]
rlabel metal3 14976 44856 14976 44856 0 Tile_X0Y0_W2MID[1]
rlabel metal2 10416 53256 10416 53256 0 Tile_X0Y0_W2MID[2]
rlabel metal2 19008 45108 19008 45108 0 Tile_X0Y0_W2MID[3]
rlabel metal2 13248 53298 13248 53298 0 Tile_X0Y0_W2MID[4]
rlabel metal3 15456 45612 15456 45612 0 Tile_X0Y0_W2MID[5]
rlabel metal3 13248 50778 13248 50778 0 Tile_X0Y0_W2MID[6]
rlabel metal2 14400 48132 14400 48132 0 Tile_X0Y0_W2MID[7]
rlabel metal3 20544 55146 20544 55146 0 Tile_X0Y0_W6END[0]
rlabel metal2 5376 51870 5376 51870 0 Tile_X0Y0_W6END[10]
rlabel metal3 20496 53340 20496 53340 0 Tile_X0Y0_W6END[11]
rlabel metal2 4992 49434 4992 49434 0 Tile_X0Y0_W6END[1]
rlabel metal3 15744 56532 15744 56532 0 Tile_X0Y0_W6END[2]
rlabel metal2 20832 51828 20832 51828 0 Tile_X0Y0_W6END[3]
rlabel metal2 13536 53928 13536 53928 0 Tile_X0Y0_W6END[4]
rlabel metal4 19584 53340 19584 53340 0 Tile_X0Y0_W6END[5]
rlabel metal3 20496 52332 20496 52332 0 Tile_X0Y0_W6END[6]
rlabel metal2 15552 52836 15552 52836 0 Tile_X0Y0_W6END[7]
rlabel metal2 20256 50274 20256 50274 0 Tile_X0Y0_W6END[8]
rlabel metal3 21330 58212 21330 58212 0 Tile_X0Y0_W6END[9]
rlabel metal2 20640 49224 20640 49224 0 Tile_X0Y0_WW4END[0]
rlabel metal3 20802 53172 20802 53172 0 Tile_X0Y0_WW4END[10]
rlabel metal2 19488 53760 19488 53760 0 Tile_X0Y0_WW4END[11]
rlabel metal3 20802 53844 20802 53844 0 Tile_X0Y0_WW4END[12]
rlabel via3 21426 54180 21426 54180 0 Tile_X0Y0_WW4END[13]
rlabel metal2 9504 53592 9504 53592 0 Tile_X0Y0_WW4END[14]
rlabel metal3 20802 54852 20802 54852 0 Tile_X0Y0_WW4END[15]
rlabel metal3 21138 50148 21138 50148 0 Tile_X0Y0_WW4END[1]
rlabel metal3 20802 50484 20802 50484 0 Tile_X0Y0_WW4END[2]
rlabel metal3 20256 50862 20256 50862 0 Tile_X0Y0_WW4END[3]
rlabel metal3 18144 51114 18144 51114 0 Tile_X0Y0_WW4END[4]
rlabel metal3 21186 51492 21186 51492 0 Tile_X0Y0_WW4END[5]
rlabel metal3 19554 51828 19554 51828 0 Tile_X0Y0_WW4END[6]
rlabel metal3 20544 52122 20544 52122 0 Tile_X0Y0_WW4END[7]
rlabel metal3 20946 52500 20946 52500 0 Tile_X0Y0_WW4END[8]
rlabel metal4 17952 50568 17952 50568 0 Tile_X0Y0_WW4END[9]
rlabel metal2 11424 74340 11424 74340 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 12960 73801 12960 73801 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit1.Q
rlabel metal3 9312 72996 9312 72996 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 8544 73962 8544 73962 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 7008 73969 7008 73969 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 5472 73626 5472 73626 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 10176 76230 10176 76230 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 8448 76650 8448 76650 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 12048 76755 12048 76755 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 10464 76986 10464 76986 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit17.Q
rlabel metal3 9648 70896 9648 70896 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 9024 71736 9024 71736 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit19.Q
rlabel metal3 2784 61572 2784 61572 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 10176 47541 10176 47541 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 8640 47208 8640 47208 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit21.Q
rlabel via1 12432 79039 12432 79039 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 10848 79086 10848 79086 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 12768 52290 12768 52290 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 12960 52248 12960 52248 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 2880 53340 2880 53340 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 2880 55062 2880 55062 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 3216 57876 3216 57876 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 3360 57582 3360 57582 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit29.Q
rlabel metal3 3648 61068 3648 61068 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 16133 59514 16133 59514 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 15360 59556 15360 59556 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 2784 66360 2784 66360 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 4320 65769 4320 65769 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 12960 76272 12960 76272 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 14592 76993 14592 76993 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 10080 74757 10080 74757 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 8544 74844 8544 74844 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 4992 45024 4992 45024 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 3504 45192 3504 45192 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 2688 60522 2688 60522 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 4704 61317 4704 61317 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 3600 66108 3600 66108 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 5184 66157 5184 66157 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 14976 78876 14976 78876 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 16560 78267 16560 78267 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 12096 72912 12096 72912 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 13632 72863 13632 72863 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit17.Q
rlabel metal3 2832 66696 2832 66696 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 4416 63385 4416 63385 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 3360 51030 3360 51030 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 2880 70560 2880 70560 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 4416 69349 4416 69349 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit21.Q
rlabel metal3 14928 76188 14928 76188 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 16608 76993 16608 76993 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit23.Q
rlabel metal3 12480 74508 12480 74508 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit24.Q
rlabel via1 14256 74503 14256 74503 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit25.Q
rlabel metal3 3312 65100 3312 65100 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 4080 64428 4080 64428 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 3360 68460 3360 68460 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 4992 68541 4992 68541 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 2880 51324 2880 51324 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 13152 78750 13152 78750 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit30.Q
rlabel via1 14736 79039 14736 79039 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 3552 52416 3552 52416 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 17664 53088 17664 53088 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 18192 51828 18192 51828 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 17760 51779 17760 51779 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 12000 71736 12000 71736 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 13488 70896 13488 70896 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 19104 74757 19104 74757 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 17568 75138 17568 75138 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit1.Q
rlabel via1 11760 69967 11760 69967 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 10176 70014 10176 70014 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 8736 61149 8736 61149 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 7200 61110 7200 61110 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 18456 72156 18456 72156 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 16800 72240 16800 72240 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 19584 48510 19584 48510 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 20064 48720 20064 48720 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 18432 50022 18432 50022 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 3168 48678 3168 48678 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 11520 67242 11520 67242 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 2688 47544 2688 47544 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 3408 48804 3408 48804 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 5856 53592 5856 53592 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 5856 52458 5856 52458 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 6240 53379 6240 53379 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 19968 54180 19968 54180 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 16512 52458 16512 52458 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit26.Q
rlabel metal3 19056 55020 19056 55020 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 15552 45654 15552 45654 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 17184 45360 17184 45360 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 9696 67914 9696 67914 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 17088 46029 17088 46029 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 5088 45864 5088 45864 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q
rlabel metal3 6192 71484 6192 71484 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 8160 71733 8160 71733 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 16608 73500 16608 73500 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 18312 72996 18312 72996 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit7.Q
rlabel via1 19248 76015 19248 76015 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 17664 76104 17664 76104 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 16224 67914 16224 67914 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 17760 67963 17760 67963 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 9552 59388 9552 59388 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 11184 57960 11184 57960 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 6816 69426 6816 69426 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 8352 69181 8352 69181 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 15648 70224 15648 70224 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 17184 70263 17184 70263 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 17472 66612 17472 66612 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit16.Q
rlabel via1 19056 66112 19056 66112 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 10656 68712 10656 68712 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 11616 67998 11616 67998 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 7968 67158 7968 67158 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit2.Q
rlabel metal2 6096 60060 6096 60060 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 7680 60361 7680 60361 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 13632 69090 13632 69090 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 15168 69433 15168 69433 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 14016 71736 14016 71736 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit24.Q
rlabel via2 15552 71481 15552 71481 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 5856 66444 5856 66444 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 7392 66787 7392 66787 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit27.Q
rlabel metal3 4992 71484 4992 71484 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 5472 70938 5472 70938 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 9504 67197 9504 67197 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit3.Q
rlabel metal3 15072 73920 15072 73920 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 16800 74757 16800 74757 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 6288 68460 6288 68460 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit4.Q
rlabel metal2 7872 68709 7872 68709 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 17664 70308 17664 70308 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit6.Q
rlabel via1 19248 69967 19248 69967 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 17664 68880 17664 68880 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit8.Q
rlabel via1 19248 68455 19248 68455 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit9.Q
rlabel metal3 17808 60312 17808 60312 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit0.Q
rlabel metal2 19632 60312 19632 60312 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 7584 58884 7584 58884 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 9072 58044 9072 58044 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit11.Q
rlabel metal2 10464 63504 10464 63504 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit12.Q
rlabel metal3 12384 63966 12384 63966 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit13.Q
rlabel metal2 13872 64428 13872 64428 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 15456 64173 15456 64173 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit15.Q
rlabel metal2 17328 64428 17328 64428 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit16.Q
rlabel metal2 19200 64344 19200 64344 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 10848 65688 10848 65688 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit18.Q
rlabel metal2 12384 65685 12384 65685 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit19.Q
rlabel metal2 10560 61665 10560 61665 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit2.Q
rlabel metal2 7584 64554 7584 64554 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit20.Q
rlabel metal2 9120 64897 9120 64897 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit21.Q
rlabel metal2 13728 65688 13728 65688 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit22.Q
rlabel via1 15312 65431 15312 65431 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit23.Q
rlabel metal2 16608 66066 16608 66066 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit24.Q
rlabel via2 18144 65433 18144 65433 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit25.Q
rlabel metal3 8544 64596 8544 64596 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 11328 64897 11328 64897 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit27.Q
rlabel metal2 6480 66780 6480 66780 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit28.Q
rlabel metal3 7632 64428 7632 64428 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 12096 62251 12096 62251 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit3.Q
rlabel metal2 13536 67000 13536 67000 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 15072 67197 15072 67197 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 7584 62706 7584 62706 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 9120 62829 9120 62829 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit5.Q
rlabel metal2 13920 62118 13920 62118 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 15456 62661 15456 62661 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit7.Q
rlabel metal3 17376 63084 17376 63084 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 19488 62622 19488 62622 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 8496 43680 8496 43680 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 10176 43967 10176 43967 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 10176 52458 10176 52458 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q
rlabel metal2 10416 52752 10416 52752 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 10560 53552 10560 53552 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
rlabel metal3 17088 55020 17088 55020 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q
rlabel metal3 16128 53508 16128 53508 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit14.Q
rlabel metal2 16224 53930 16224 53930 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
rlabel metal2 13344 58296 13344 58296 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 11712 58506 11712 58506 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 6816 58298 6816 58298 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit18.Q
rlabel metal2 5280 58506 5280 58506 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit19.Q
rlabel metal2 18192 44268 18192 44268 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 4704 59637 4704 59637 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit20.Q
rlabel metal2 2976 58380 2976 58380 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit21.Q
rlabel metal2 14784 60361 14784 60361 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit22.Q
rlabel metal2 13248 60018 13248 60018 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit23.Q
rlabel metal2 17376 58674 17376 58674 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 19200 58800 19200 58800 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 9600 56994 9600 56994 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit26.Q
rlabel metal2 11136 56786 11136 56786 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 10704 60312 10704 60312 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit28.Q
rlabel via1 12336 60895 12336 60895 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit29.Q
rlabel via1 19824 44263 19824 44263 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit3.Q
rlabel metal2 16080 60900 16080 60900 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit30.Q
rlabel metal2 17664 61149 17664 61149 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit31.Q
rlabel metal3 13200 43260 13200 43260 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q
rlabel metal2 14304 44352 14304 44352 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit5.Q
rlabel metal2 13824 44436 13824 44436 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 5856 45696 5856 45696 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 8256 46032 8256 46032 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit8.Q
rlabel metal2 6240 46515 6240 46515 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
rlabel metal2 15456 49938 15456 49938 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 15648 49896 15648 49896 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit1.Q
rlabel metal2 19488 57414 19488 57414 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 19488 56063 19488 56063 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q
rlabel metal2 14352 45948 14352 45948 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit12.Q
rlabel metal3 12768 45948 12768 45948 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit13.Q
rlabel metal2 2976 46410 2976 46410 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit14.Q
rlabel metal2 4416 46830 4416 46830 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit15.Q
rlabel metal2 3168 53970 3168 53970 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit16.Q
rlabel metal2 4704 54061 4704 54061 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit17.Q
rlabel metal2 13824 56406 13824 56406 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 15360 56991 15360 56991 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit19.Q
rlabel metal2 16992 49011 16992 49011 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q
rlabel metal2 13152 49224 13152 49224 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit20.Q
rlabel via2 12960 49478 12960 49478 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit21.Q
rlabel metal2 8064 50946 8064 50946 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit22.Q
rlabel via1 9648 50992 9648 50992 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit23.Q
rlabel metal2 9792 49434 9792 49434 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit24.Q
rlabel metal2 11376 48967 11376 48967 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit25.Q
rlabel metal3 12912 53340 12912 53340 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit26.Q
rlabel via1 14736 53335 14736 53335 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 19968 45619 19968 45619 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit28.Q
rlabel metal2 18528 43680 18528 43680 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit29.Q
rlabel metal3 5904 50064 5904 50064 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 10176 46410 10176 46410 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit30.Q
rlabel metal2 11712 46034 11712 46034 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit31.Q
rlabel metal3 7488 49728 7488 49728 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit4.Q
rlabel via2 7296 48801 7296 48801 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q
rlabel metal2 8160 55650 8160 55650 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q
rlabel metal2 8352 55608 8352 55608 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit7.Q
rlabel metal3 7248 55020 7248 55020 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 19008 57834 19008 57834 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 4416 50148 4416 50148 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit10.Q
rlabel metal2 2880 49777 2880 49777 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit11.Q
rlabel metal2 3072 57330 3072 57330 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 4848 56532 4848 56532 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit13.Q
rlabel metal2 13728 56994 13728 56994 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 15264 57379 15264 57379 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit15.Q
rlabel metal3 13728 50400 13728 50400 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit16.Q
rlabel metal2 13248 51289 13248 51289 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit17.Q
rlabel metal2 6192 51240 6192 51240 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit18.Q
rlabel via1 6768 51823 6768 51823 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit19.Q
rlabel metal2 9552 48972 9552 48972 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 11664 48216 11664 48216 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit21.Q
rlabel metal3 12864 53508 12864 53508 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 14496 54313 14496 54313 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit23.Q
rlabel metal3 19488 50400 19488 50400 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit24.Q
rlabel metal2 18624 51289 18624 51289 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit25.Q
rlabel metal2 10368 55608 10368 55608 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit26.Q
rlabel metal2 11976 55524 11976 55524 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit27.Q
rlabel metal2 8352 44478 8352 44478 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit28.Q
rlabel metal2 8736 45360 8736 45360 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit29.Q
rlabel metal2 18528 46746 18528 46746 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit30.Q
rlabel via2 20064 46454 20064 46454 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 14064 47460 14064 47460 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit8.Q
rlabel metal2 12480 47460 12480 47460 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit9.Q
rlabel metal3 16608 58632 16608 58632 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E1BEG0
rlabel metal3 15360 59430 15360 59430 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E1BEG1
rlabel metal3 14688 59640 14688 59640 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E1BEG2
rlabel metal3 17520 60816 17520 60816 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E1BEG3
rlabel metal2 19872 58590 19872 58590 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG0
rlabel metal2 11424 57162 11424 57162 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG1
rlabel metal2 12480 61110 12480 61110 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG2
rlabel metal3 18432 61068 18432 61068 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG3
rlabel metal2 19824 61068 19824 61068 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG4
rlabel metal3 15456 61656 15456 61656 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG5
rlabel metal2 19680 62496 19680 62496 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG6
rlabel metal3 17856 62328 17856 62328 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG7
rlabel metal2 19488 63084 19488 63084 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb0
rlabel metal2 13824 59472 13824 59472 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb1
rlabel metal2 19392 63924 19392 63924 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb2
rlabel metal3 17712 63840 17712 63840 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb3
rlabel metal2 19392 64470 19392 64470 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb4
rlabel metal2 19008 65310 19008 65310 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb5
rlabel metal2 19776 64554 19776 64554 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb6
rlabel metal3 17616 65352 17616 65352 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb7
rlabel metal3 17616 71652 17616 71652 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG0
rlabel metal3 11712 72702 11712 72702 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG1
rlabel metal5 16080 75936 16080 75936 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG10
rlabel metal2 18624 71988 18624 71988 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG11
rlabel metal3 7440 71400 7440 71400 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG2
rlabel metal3 18432 74424 18432 74424 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG3
rlabel via1 19470 74430 19470 74430 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG4
rlabel metal3 11856 72996 11856 72996 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG5
rlabel metal2 18624 72744 18624 72744 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG6
rlabel metal3 18720 72996 18720 72996 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG7
rlabel metal3 19536 76104 19536 76104 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG8
rlabel metal2 11904 70854 11904 70854 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG9
rlabel metal3 18864 65520 18864 65520 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG0
rlabel metal3 15648 66192 15648 66192 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG1
rlabel metal2 18912 71484 18912 71484 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG10
rlabel metal2 17376 70182 17376 70182 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG11
rlabel metal3 17904 69216 17904 69216 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG12
rlabel metal2 12384 70014 12384 70014 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG13
rlabel metal5 15504 72240 15504 72240 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG14
rlabel metal3 17328 72240 17328 72240 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG15
rlabel metal2 19440 65352 19440 65352 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG2
rlabel metal3 17520 67116 17520 67116 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG3
rlabel metal2 19968 68166 19968 68166 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG4
rlabel metal2 9696 67284 9696 67284 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG5
rlabel metal2 18912 68838 18912 68838 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG6
rlabel metal2 19776 69258 19776 69258 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG7
rlabel metal2 19536 68628 19536 68628 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG8
rlabel metal3 16608 70728 16608 70728 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG9
rlabel metal2 18720 70602 18720 70602 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG0
rlabel metal2 7344 51828 7344 51828 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG1
rlabel metal2 10656 50778 10656 50778 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG2
rlabel metal2 14208 53676 14208 53676 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG3
rlabel metal3 19200 50988 19200 50988 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG4
rlabel metal3 11808 54012 11808 54012 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG5
rlabel metal3 9072 46872 9072 46872 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG6
rlabel metal3 19536 48048 19536 48048 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG7
rlabel metal2 6720 53592 6720 53592 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG10
rlabel metal3 18912 54054 18912 54054 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG11
rlabel metal2 13056 48090 13056 48090 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG12
rlabel metal2 3840 49602 3840 49602 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG13
rlabel metal3 3600 51828 3600 51828 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG14
rlabel metal2 15072 71526 15072 71526 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG15
rlabel metal2 16080 48720 16080 48720 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG4
rlabel metal3 7008 69132 7008 69132 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG5
rlabel metal3 6624 55020 6624 55020 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG6
rlabel metal2 17184 53970 17184 53970 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG7
rlabel metal2 16512 48720 16512 48720 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG8
rlabel metal2 6912 67410 6912 67410 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG9
rlabel metal5 1844 83496 1844 83496 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1BEG0
rlabel metal4 2112 66444 2112 66444 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1BEG1
rlabel metal3 3840 58296 3840 58296 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1BEG2
rlabel metal2 1968 76860 1968 76860 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1BEG3
rlabel metal3 14640 13104 14640 13104 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END0
rlabel metal4 3264 43596 3264 43596 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END1
rlabel metal2 12816 36036 12816 36036 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END2
rlabel metal2 14832 36792 14832 36792 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END3
rlabel metal2 13056 51240 13056 51240 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG0
rlabel metal3 2592 83496 2592 83496 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG1
rlabel metal3 3600 82824 3600 82824 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG2
rlabel metal2 3312 83496 3312 83496 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG3
rlabel metal3 4128 82782 4128 82782 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG4
rlabel metal3 3168 83328 3168 83328 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG5
rlabel metal3 6720 84336 6720 84336 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG6
rlabel metal3 4032 83538 4032 83538 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG7
rlabel metal3 6240 82824 6240 82824 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb0
rlabel metal2 4416 83412 4416 83412 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb1
rlabel metal3 5184 83160 5184 83160 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb2
rlabel metal2 5184 83370 5184 83370 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb3
rlabel metal2 5568 83580 5568 83580 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb4
rlabel metal3 9024 83496 9024 83496 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb5
rlabel metal3 8112 83160 8112 83160 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb6
rlabel metal3 6222 83496 6222 83496 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb7
rlabel metal3 15264 83496 15264 83496 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N4BEG0
rlabel metal2 8256 49770 8256 49770 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N4BEG1
rlabel metal3 7680 57288 7680 57288 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N4BEG2
rlabel metal2 18096 83496 18096 83496 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N4BEG3
rlabel metal2 13008 47796 13008 47796 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG0
rlabel metal3 10080 1260 10080 1260 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG1
rlabel metal2 11088 1176 11088 1176 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG2
rlabel metal3 13584 50064 13584 50064 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG3
rlabel metal4 11616 21714 11616 21714 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG4
rlabel metal2 11904 43302 11904 43302 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG5
rlabel metal3 10080 39732 10080 39732 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG6
rlabel metal3 12048 1848 12048 1848 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG7
rlabel metal5 14648 17640 14648 17640 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S4BEG0
rlabel metal5 9606 1260 9606 1260 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S4BEG1
rlabel metal4 11712 27468 11712 27468 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S4BEG2
rlabel metal3 16416 35280 16416 35280 0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S4BEG3
rlabel metal3 6768 83160 6768 83160 0 Tile_X0Y0_W_TT_IF2_top.N4BEG_outbuf_10.A
rlabel metal3 13584 83496 13584 83496 0 Tile_X0Y0_W_TT_IF2_top.N4BEG_outbuf_11.A
rlabel metal3 16080 83496 16080 83496 0 Tile_X0Y0_W_TT_IF2_top.N4BEG_outbuf_8.A
rlabel metal3 7104 83496 7104 83496 0 Tile_X0Y0_W_TT_IF2_top.N4BEG_outbuf_9.A
rlabel metal2 19488 16590 19488 16590 0 Tile_X0Y1_E1BEG[0]
rlabel metal3 15120 16632 15120 16632 0 Tile_X0Y1_E1BEG[1]
rlabel metal2 3648 16086 3648 16086 0 Tile_X0Y1_E1BEG[2]
rlabel metal2 16416 17388 16416 17388 0 Tile_X0Y1_E1BEG[3]
rlabel metal2 17856 16968 17856 16968 0 Tile_X0Y1_E2BEG[0]
rlabel metal2 17472 17136 17472 17136 0 Tile_X0Y1_E2BEG[1]
rlabel metal2 16800 18102 16800 18102 0 Tile_X0Y1_E2BEG[2]
rlabel metal3 21234 18564 21234 18564 0 Tile_X0Y1_E2BEG[3]
rlabel metal3 21282 18900 21282 18900 0 Tile_X0Y1_E2BEG[4]
rlabel metal2 17184 17262 17184 17262 0 Tile_X0Y1_E2BEG[5]
rlabel metal2 20400 14196 20400 14196 0 Tile_X0Y1_E2BEG[6]
rlabel metal2 20256 13734 20256 13734 0 Tile_X0Y1_E2BEG[7]
rlabel metal3 17376 16380 17376 16380 0 Tile_X0Y1_E2BEGb[0]
rlabel metal3 21378 20580 21378 20580 0 Tile_X0Y1_E2BEGb[1]
rlabel metal3 21282 20916 21282 20916 0 Tile_X0Y1_E2BEGb[2]
rlabel metal3 21330 21252 21330 21252 0 Tile_X0Y1_E2BEGb[3]
rlabel metal3 21042 21588 21042 21588 0 Tile_X0Y1_E2BEGb[4]
rlabel metal3 21042 21924 21042 21924 0 Tile_X0Y1_E2BEGb[5]
rlabel metal2 15456 22554 15456 22554 0 Tile_X0Y1_E2BEGb[6]
rlabel metal3 21138 22596 21138 22596 0 Tile_X0Y1_E2BEGb[7]
rlabel metal2 19536 30912 19536 30912 0 Tile_X0Y1_E6BEG[0]
rlabel metal2 20256 30366 20256 30366 0 Tile_X0Y1_E6BEG[10]
rlabel metal4 19872 33096 19872 33096 0 Tile_X0Y1_E6BEG[11]
rlabel metal3 20514 28644 20514 28644 0 Tile_X0Y1_E6BEG[1]
rlabel metal3 20802 28980 20802 28980 0 Tile_X0Y1_E6BEG[2]
rlabel via2 21426 29316 21426 29316 0 Tile_X0Y1_E6BEG[3]
rlabel metal2 19968 30030 19968 30030 0 Tile_X0Y1_E6BEG[4]
rlabel metal2 20736 28854 20736 28854 0 Tile_X0Y1_E6BEG[5]
rlabel metal4 20640 29442 20640 29442 0 Tile_X0Y1_E6BEG[6]
rlabel metal2 20640 29988 20640 29988 0 Tile_X0Y1_E6BEG[7]
rlabel metal3 21378 30996 21378 30996 0 Tile_X0Y1_E6BEG[8]
rlabel metal2 17424 30828 17424 30828 0 Tile_X0Y1_E6BEG[9]
rlabel via2 21426 22932 21426 22932 0 Tile_X0Y1_EE4BEG[0]
rlabel metal3 20802 26292 20802 26292 0 Tile_X0Y1_EE4BEG[10]
rlabel metal3 21186 26628 21186 26628 0 Tile_X0Y1_EE4BEG[11]
rlabel metal3 20994 26964 20994 26964 0 Tile_X0Y1_EE4BEG[12]
rlabel metal2 15456 27132 15456 27132 0 Tile_X0Y1_EE4BEG[13]
rlabel metal2 16848 30408 16848 30408 0 Tile_X0Y1_EE4BEG[14]
rlabel metal3 20544 27930 20544 27930 0 Tile_X0Y1_EE4BEG[15]
rlabel metal3 20256 23226 20256 23226 0 Tile_X0Y1_EE4BEG[1]
rlabel metal3 18384 29652 18384 29652 0 Tile_X0Y1_EE4BEG[2]
rlabel metal3 21024 23898 21024 23898 0 Tile_X0Y1_EE4BEG[3]
rlabel metal3 21138 24276 21138 24276 0 Tile_X0Y1_EE4BEG[4]
rlabel metal3 18384 21000 18384 21000 0 Tile_X0Y1_EE4BEG[5]
rlabel metal3 20994 24948 20994 24948 0 Tile_X0Y1_EE4BEG[6]
rlabel metal2 17376 25494 17376 25494 0 Tile_X0Y1_EE4BEG[7]
rlabel metal3 18192 29232 18192 29232 0 Tile_X0Y1_EE4BEG[8]
rlabel metal3 20994 25956 20994 25956 0 Tile_X0Y1_EE4BEG[9]
rlabel metal2 1296 11004 1296 11004 0 Tile_X0Y1_FrameData[0]
rlabel metal2 1248 38052 1248 38052 0 Tile_X0Y1_FrameData[10]
rlabel metal3 1392 40404 1392 40404 0 Tile_X0Y1_FrameData[11]
rlabel metal3 654 65772 654 65772 0 Tile_X0Y1_FrameData[12]
rlabel via2 78 66444 78 66444 0 Tile_X0Y1_FrameData[13]
rlabel metal3 558 67116 558 67116 0 Tile_X0Y1_FrameData[14]
rlabel metal3 1086 67788 1086 67788 0 Tile_X0Y1_FrameData[15]
rlabel metal3 414 68460 414 68460 0 Tile_X0Y1_FrameData[16]
rlabel metal3 318 69132 318 69132 0 Tile_X0Y1_FrameData[17]
rlabel metal2 1296 39732 1296 39732 0 Tile_X0Y1_FrameData[18]
rlabel metal3 462 70476 462 70476 0 Tile_X0Y1_FrameData[19]
rlabel metal2 1824 12222 1824 12222 0 Tile_X0Y1_FrameData[1]
rlabel metal3 222 71148 222 71148 0 Tile_X0Y1_FrameData[20]
rlabel metal3 990 71820 990 71820 0 Tile_X0Y1_FrameData[21]
rlabel metal3 126 72492 126 72492 0 Tile_X0Y1_FrameData[22]
rlabel metal3 990 73164 990 73164 0 Tile_X0Y1_FrameData[23]
rlabel metal3 174 73836 174 73836 0 Tile_X0Y1_FrameData[24]
rlabel metal3 1038 74508 1038 74508 0 Tile_X0Y1_FrameData[25]
rlabel metal3 1920 40320 1920 40320 0 Tile_X0Y1_FrameData[26]
rlabel metal3 174 75852 174 75852 0 Tile_X0Y1_FrameData[27]
rlabel metal3 366 76524 366 76524 0 Tile_X0Y1_FrameData[28]
rlabel metal3 798 77196 798 77196 0 Tile_X0Y1_FrameData[29]
rlabel metal2 1392 42756 1392 42756 0 Tile_X0Y1_FrameData[2]
rlabel via3 78 77868 78 77868 0 Tile_X0Y1_FrameData[30]
rlabel metal3 126 78540 126 78540 0 Tile_X0Y1_FrameData[31]
rlabel metal2 1728 18648 1728 18648 0 Tile_X0Y1_FrameData[3]
rlabel metal2 1920 9030 1920 9030 0 Tile_X0Y1_FrameData[4]
rlabel metal3 1728 17220 1728 17220 0 Tile_X0Y1_FrameData[5]
rlabel metal2 18816 32508 18816 32508 0 Tile_X0Y1_FrameData[6]
rlabel metal2 1440 10164 1440 10164 0 Tile_X0Y1_FrameData[7]
rlabel metal2 17424 13188 17424 13188 0 Tile_X0Y1_FrameData[8]
rlabel metal2 18720 13146 18720 13146 0 Tile_X0Y1_FrameData[9]
rlabel metal4 20736 31206 20736 31206 0 Tile_X0Y1_FrameData_O[0]
rlabel metal2 19728 34608 19728 34608 0 Tile_X0Y1_FrameData_O[10]
rlabel metal2 20016 35028 20016 35028 0 Tile_X0Y1_FrameData_O[11]
rlabel metal4 19680 35700 19680 35700 0 Tile_X0Y1_FrameData_O[12]
rlabel metal3 20802 36708 20802 36708 0 Tile_X0Y1_FrameData_O[13]
rlabel metal3 20544 37002 20544 37002 0 Tile_X0Y1_FrameData_O[14]
rlabel metal3 20850 37380 20850 37380 0 Tile_X0Y1_FrameData_O[15]
rlabel metal3 20082 37716 20082 37716 0 Tile_X0Y1_FrameData_O[16]
rlabel metal3 20850 38052 20850 38052 0 Tile_X0Y1_FrameData_O[17]
rlabel metal3 20466 38388 20466 38388 0 Tile_X0Y1_FrameData_O[18]
rlabel metal3 20466 38724 20466 38724 0 Tile_X0Y1_FrameData_O[19]
rlabel metal3 21408 32634 21408 32634 0 Tile_X0Y1_FrameData_O[1]
rlabel metal3 20658 39060 20658 39060 0 Tile_X0Y1_FrameData_O[20]
rlabel metal3 19824 39480 19824 39480 0 Tile_X0Y1_FrameData_O[21]
rlabel metal2 19872 39648 19872 39648 0 Tile_X0Y1_FrameData_O[22]
rlabel metal2 19200 40110 19200 40110 0 Tile_X0Y1_FrameData_O[23]
rlabel metal2 18048 40488 18048 40488 0 Tile_X0Y1_FrameData_O[24]
rlabel metal2 19584 40698 19584 40698 0 Tile_X0Y1_FrameData_O[25]
rlabel metal3 20466 41076 20466 41076 0 Tile_X0Y1_FrameData_O[26]
rlabel metal3 20658 41412 20658 41412 0 Tile_X0Y1_FrameData_O[27]
rlabel metal3 20466 41748 20466 41748 0 Tile_X0Y1_FrameData_O[28]
rlabel metal3 20658 42084 20658 42084 0 Tile_X0Y1_FrameData_O[29]
rlabel metal2 19968 32256 19968 32256 0 Tile_X0Y1_FrameData_O[2]
rlabel metal2 18144 42294 18144 42294 0 Tile_X0Y1_FrameData_O[30]
rlabel metal3 20850 42756 20850 42756 0 Tile_X0Y1_FrameData_O[31]
rlabel metal2 18768 33096 18768 33096 0 Tile_X0Y1_FrameData_O[3]
rlabel via3 21426 33684 21426 33684 0 Tile_X0Y1_FrameData_O[4]
rlabel metal3 20544 34062 20544 34062 0 Tile_X0Y1_FrameData_O[5]
rlabel metal3 20802 34356 20802 34356 0 Tile_X0Y1_FrameData_O[6]
rlabel metal3 20802 34692 20802 34692 0 Tile_X0Y1_FrameData_O[7]
rlabel metal4 19968 34440 19968 34440 0 Tile_X0Y1_FrameData_O[8]
rlabel metal4 20736 34650 20736 34650 0 Tile_X0Y1_FrameData_O[9]
rlabel metal2 2496 70014 2496 70014 0 Tile_X0Y1_FrameStrobe[0]
rlabel metal2 17760 282 17760 282 0 Tile_X0Y1_FrameStrobe[10]
rlabel metal2 17952 198 17952 198 0 Tile_X0Y1_FrameStrobe[11]
rlabel metal2 18144 618 18144 618 0 Tile_X0Y1_FrameStrobe[12]
rlabel metal2 18336 114 18336 114 0 Tile_X0Y1_FrameStrobe[13]
rlabel metal2 18528 618 18528 618 0 Tile_X0Y1_FrameStrobe[14]
rlabel metal2 18720 576 18720 576 0 Tile_X0Y1_FrameStrobe[15]
rlabel metal2 18912 618 18912 618 0 Tile_X0Y1_FrameStrobe[16]
rlabel metal2 19104 702 19104 702 0 Tile_X0Y1_FrameStrobe[17]
rlabel metal2 19296 618 19296 618 0 Tile_X0Y1_FrameStrobe[18]
rlabel metal2 19488 72 19488 72 0 Tile_X0Y1_FrameStrobe[19]
rlabel metal2 2448 38220 2448 38220 0 Tile_X0Y1_FrameStrobe[1]
rlabel metal2 2496 19656 2496 19656 0 Tile_X0Y1_FrameStrobe[2]
rlabel metal2 16416 576 16416 576 0 Tile_X0Y1_FrameStrobe[3]
rlabel metal2 16608 660 16608 660 0 Tile_X0Y1_FrameStrobe[4]
rlabel metal2 2496 14910 2496 14910 0 Tile_X0Y1_FrameStrobe[5]
rlabel metal2 2400 47166 2400 47166 0 Tile_X0Y1_FrameStrobe[6]
rlabel metal2 2496 51156 2496 51156 0 Tile_X0Y1_FrameStrobe[7]
rlabel metal2 17376 954 17376 954 0 Tile_X0Y1_FrameStrobe[8]
rlabel metal2 17568 954 17568 954 0 Tile_X0Y1_FrameStrobe[9]
rlabel metal2 1824 4902 1824 4902 0 Tile_X0Y1_N1END[0]
rlabel metal2 1968 10752 1968 10752 0 Tile_X0Y1_N1END[1]
rlabel metal2 2496 17682 2496 17682 0 Tile_X0Y1_N1END[2]
rlabel metal2 2400 3180 2400 3180 0 Tile_X0Y1_N1END[3]
rlabel metal2 4128 996 4128 996 0 Tile_X0Y1_N2END[0]
rlabel metal2 4320 282 4320 282 0 Tile_X0Y1_N2END[1]
rlabel metal3 4272 13188 4272 13188 0 Tile_X0Y1_N2END[2]
rlabel metal2 5328 13188 5328 13188 0 Tile_X0Y1_N2END[3]
rlabel metal2 4896 114 4896 114 0 Tile_X0Y1_N2END[4]
rlabel metal2 5088 156 5088 156 0 Tile_X0Y1_N2END[5]
rlabel metal2 5280 282 5280 282 0 Tile_X0Y1_N2END[6]
rlabel metal2 5472 324 5472 324 0 Tile_X0Y1_N2END[7]
rlabel metal2 2592 492 2592 492 0 Tile_X0Y1_N2MID[0]
rlabel metal2 2784 324 2784 324 0 Tile_X0Y1_N2MID[1]
rlabel metal2 2976 660 2976 660 0 Tile_X0Y1_N2MID[2]
rlabel metal2 10464 10206 10464 10206 0 Tile_X0Y1_N2MID[3]
rlabel via2 3360 72 3360 72 0 Tile_X0Y1_N2MID[4]
rlabel metal2 3552 450 3552 450 0 Tile_X0Y1_N2MID[5]
rlabel metal2 3744 618 3744 618 0 Tile_X0Y1_N2MID[6]
rlabel metal2 3936 198 3936 198 0 Tile_X0Y1_N2MID[7]
rlabel metal2 5664 408 5664 408 0 Tile_X0Y1_N4END[0]
rlabel metal2 7584 744 7584 744 0 Tile_X0Y1_N4END[10]
rlabel metal2 7776 1038 7776 1038 0 Tile_X0Y1_N4END[11]
rlabel metal2 7968 954 7968 954 0 Tile_X0Y1_N4END[12]
rlabel metal2 8160 702 8160 702 0 Tile_X0Y1_N4END[13]
rlabel metal2 8352 660 8352 660 0 Tile_X0Y1_N4END[14]
rlabel metal2 8544 492 8544 492 0 Tile_X0Y1_N4END[15]
rlabel metal2 2352 16380 2352 16380 0 Tile_X0Y1_N4END[1]
rlabel metal2 6048 660 6048 660 0 Tile_X0Y1_N4END[2]
rlabel metal2 6240 114 6240 114 0 Tile_X0Y1_N4END[3]
rlabel metal2 6432 240 6432 240 0 Tile_X0Y1_N4END[4]
rlabel metal2 6624 576 6624 576 0 Tile_X0Y1_N4END[5]
rlabel metal2 6816 660 6816 660 0 Tile_X0Y1_N4END[6]
rlabel via2 7008 72 7008 72 0 Tile_X0Y1_N4END[7]
rlabel metal2 5952 1680 5952 1680 0 Tile_X0Y1_N4END[8]
rlabel metal2 7392 618 7392 618 0 Tile_X0Y1_N4END[9]
rlabel metal2 8736 492 8736 492 0 Tile_X0Y1_S1BEG[0]
rlabel metal2 8928 870 8928 870 0 Tile_X0Y1_S1BEG[1]
rlabel metal2 9120 282 9120 282 0 Tile_X0Y1_S1BEG[2]
rlabel metal2 9312 870 9312 870 0 Tile_X0Y1_S1BEG[3]
rlabel metal2 9504 366 9504 366 0 Tile_X0Y1_S2BEG[0]
rlabel metal2 9696 450 9696 450 0 Tile_X0Y1_S2BEG[1]
rlabel metal2 9888 408 9888 408 0 Tile_X0Y1_S2BEG[2]
rlabel metal2 10080 870 10080 870 0 Tile_X0Y1_S2BEG[3]
rlabel metal2 10272 324 10272 324 0 Tile_X0Y1_S2BEG[4]
rlabel metal2 10464 1290 10464 1290 0 Tile_X0Y1_S2BEG[5]
rlabel metal2 10656 450 10656 450 0 Tile_X0Y1_S2BEG[6]
rlabel metal2 10848 744 10848 744 0 Tile_X0Y1_S2BEG[7]
rlabel metal2 11040 408 11040 408 0 Tile_X0Y1_S2BEGb[0]
rlabel metal2 11232 492 11232 492 0 Tile_X0Y1_S2BEGb[1]
rlabel metal2 11424 492 11424 492 0 Tile_X0Y1_S2BEGb[2]
rlabel metal2 11616 1890 11616 1890 0 Tile_X0Y1_S2BEGb[3]
rlabel metal2 11808 492 11808 492 0 Tile_X0Y1_S2BEGb[4]
rlabel metal2 11232 1386 11232 1386 0 Tile_X0Y1_S2BEGb[5]
rlabel metal3 10752 1302 10752 1302 0 Tile_X0Y1_S2BEGb[6]
rlabel metal2 12384 870 12384 870 0 Tile_X0Y1_S2BEGb[7]
rlabel metal2 12576 534 12576 534 0 Tile_X0Y1_S4BEG[0]
rlabel metal2 14496 702 14496 702 0 Tile_X0Y1_S4BEG[10]
rlabel metal2 14688 492 14688 492 0 Tile_X0Y1_S4BEG[11]
rlabel metal2 14880 870 14880 870 0 Tile_X0Y1_S4BEG[12]
rlabel metal2 15072 450 15072 450 0 Tile_X0Y1_S4BEG[13]
rlabel metal3 14880 2436 14880 2436 0 Tile_X0Y1_S4BEG[14]
rlabel metal2 15456 744 15456 744 0 Tile_X0Y1_S4BEG[15]
rlabel metal2 12768 870 12768 870 0 Tile_X0Y1_S4BEG[1]
rlabel metal2 12960 282 12960 282 0 Tile_X0Y1_S4BEG[2]
rlabel metal2 13152 198 13152 198 0 Tile_X0Y1_S4BEG[3]
rlabel metal2 13344 240 13344 240 0 Tile_X0Y1_S4BEG[4]
rlabel metal2 13536 492 13536 492 0 Tile_X0Y1_S4BEG[5]
rlabel metal2 13728 660 13728 660 0 Tile_X0Y1_S4BEG[6]
rlabel metal2 13920 786 13920 786 0 Tile_X0Y1_S4BEG[7]
rlabel metal2 14016 1596 14016 1596 0 Tile_X0Y1_S4BEG[8]
rlabel metal2 14304 492 14304 492 0 Tile_X0Y1_S4BEG[9]
rlabel metal2 15648 660 15648 660 0 Tile_X0Y1_UserCLK
rlabel metal2 17712 1764 17712 1764 0 Tile_X0Y1_W1END[0]
rlabel metal3 9894 1512 9894 1512 0 Tile_X0Y1_W1END[1]
rlabel metal3 21426 756 21426 756 0 Tile_X0Y1_W1END[2]
rlabel metal3 21378 1092 21378 1092 0 Tile_X0Y1_W1END[3]
rlabel metal2 15936 5628 15936 5628 0 Tile_X0Y1_W2END[0]
rlabel metal2 9216 7812 9216 7812 0 Tile_X0Y1_W2END[1]
rlabel via2 6144 11508 6144 11508 0 Tile_X0Y1_W2END[2]
rlabel metal2 1248 13524 1248 13524 0 Tile_X0Y1_W2END[3]
rlabel metal2 11808 10878 11808 10878 0 Tile_X0Y1_W2END[4]
rlabel metal2 4032 13986 4032 13986 0 Tile_X0Y1_W2END[5]
rlabel metal3 18144 14406 18144 14406 0 Tile_X0Y1_W2END[6]
rlabel metal3 21378 6468 21378 6468 0 Tile_X0Y1_W2END[7]
rlabel metal3 15840 1806 15840 1806 0 Tile_X0Y1_W2MID[0]
rlabel metal3 21426 1764 21426 1764 0 Tile_X0Y1_W2MID[1]
rlabel metal3 20802 2100 20802 2100 0 Tile_X0Y1_W2MID[2]
rlabel metal3 20802 2436 20802 2436 0 Tile_X0Y1_W2MID[3]
rlabel metal2 11616 10836 11616 10836 0 Tile_X0Y1_W2MID[4]
rlabel metal3 12816 11256 12816 11256 0 Tile_X0Y1_W2MID[5]
rlabel metal3 13842 3444 13842 3444 0 Tile_X0Y1_W2MID[6]
rlabel metal2 13584 14028 13584 14028 0 Tile_X0Y1_W2MID[7]
rlabel metal2 19248 12432 19248 12432 0 Tile_X0Y1_W6END[0]
rlabel metal4 16416 15456 16416 15456 0 Tile_X0Y1_W6END[10]
rlabel metal3 12432 16044 12432 16044 0 Tile_X0Y1_W6END[11]
rlabel metal2 5664 30534 5664 30534 0 Tile_X0Y1_W6END[1]
rlabel metal2 7872 12684 7872 12684 0 Tile_X0Y1_W6END[2]
rlabel metal3 11424 14658 11424 14658 0 Tile_X0Y1_W6END[3]
rlabel metal3 12816 13188 12816 13188 0 Tile_X0Y1_W6END[4]
rlabel metal4 18048 14910 18048 14910 0 Tile_X0Y1_W6END[5]
rlabel metal2 7728 17724 7728 17724 0 Tile_X0Y1_W6END[6]
rlabel metal2 14064 14700 14064 14700 0 Tile_X0Y1_W6END[7]
rlabel metal2 16608 11928 16608 11928 0 Tile_X0Y1_W6END[8]
rlabel metal2 8160 16884 8160 16884 0 Tile_X0Y1_W6END[9]
rlabel metal2 18624 12558 18624 12558 0 Tile_X0Y1_WW4END[0]
rlabel metal3 14544 19488 14544 19488 0 Tile_X0Y1_WW4END[10]
rlabel metal3 13968 25452 13968 25452 0 Tile_X0Y1_WW4END[11]
rlabel metal2 15984 12684 15984 12684 0 Tile_X0Y1_WW4END[12]
rlabel metal5 15832 11214 15832 11214 0 Tile_X0Y1_WW4END[13]
rlabel metal3 17616 11424 17616 11424 0 Tile_X0Y1_WW4END[14]
rlabel metal3 17760 24612 17760 24612 0 Tile_X0Y1_WW4END[15]
rlabel metal4 14784 14910 14784 14910 0 Tile_X0Y1_WW4END[1]
rlabel metal3 5616 7476 5616 7476 0 Tile_X0Y1_WW4END[2]
rlabel metal2 13440 26628 13440 26628 0 Tile_X0Y1_WW4END[3]
rlabel metal2 19296 10332 19296 10332 0 Tile_X0Y1_WW4END[4]
rlabel metal3 15744 8064 15744 8064 0 Tile_X0Y1_WW4END[5]
rlabel metal3 3168 22260 3168 22260 0 Tile_X0Y1_WW4END[6]
rlabel metal3 20016 24528 20016 24528 0 Tile_X0Y1_WW4END[7]
rlabel metal2 19152 12264 19152 12264 0 Tile_X0Y1_WW4END[8]
rlabel metal4 5568 20286 5568 20286 0 Tile_X0Y1_WW4END[9]
rlabel metal2 12192 37632 12192 37632 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 13776 37632 13776 37632 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit1.Q
rlabel metal3 9360 36540 9360 36540 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 12192 35952 12192 35952 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 5184 17766 5184 17766 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 2160 17808 2160 17808 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 9408 11046 9408 11046 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 9792 10206 9792 10206 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 9696 41874 9696 41874 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit16.Q
rlabel metal3 9744 40656 9744 40656 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 8544 41874 8544 41874 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 10080 41283 10080 41283 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit19.Q
rlabel metal3 3312 41244 3312 41244 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 9408 40026 9408 40026 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit20.Q
rlabel metal3 9888 37632 9888 37632 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 10176 38640 10176 38640 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 11712 38469 11712 38469 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit23.Q
rlabel via1 14861 9492 14861 9492 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 13920 8820 13920 8820 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 3394 32679 3394 32679 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q
rlabel metal3 4032 32172 4032 32172 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 4224 16296 4224 16296 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 4704 17640 4704 17640 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit29.Q
rlabel via1 5328 41239 5328 41239 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit3.Q
rlabel via1 15045 21588 15045 21588 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 14784 21294 14784 21294 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 2496 38640 2496 38640 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit4.Q
rlabel metal3 3120 36876 3120 36876 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit5.Q
rlabel metal3 12336 39732 12336 39732 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit6.Q
rlabel metal3 13248 39060 13248 39060 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 8544 15120 8544 15120 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q
rlabel metal3 8832 14196 8832 14196 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit9.Q
rlabel metal3 3552 12474 3552 12474 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 6432 13440 6432 13440 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 2688 39060 2688 39060 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 5376 40149 5376 40149 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 2736 33096 2736 33096 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 4560 35931 4560 35931 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 14400 42210 14400 42210 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 15984 41979 15984 41979 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 13248 36750 13248 36750 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 14688 35280 14688 35280 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 2736 39900 2736 39900 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit18.Q
rlabel metal3 4320 42168 4320 42168 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 6048 14196 6048 14196 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 2640 32340 2640 32340 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit20.Q
rlabel metal3 3408 33432 3408 33432 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 14112 40950 14112 40950 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit22.Q
rlabel via1 15984 41239 15984 41239 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 14400 38850 14400 38850 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 16080 38388 16080 38388 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 3264 41664 3264 41664 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 5760 42217 5760 42217 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 2736 34608 2736 34608 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 4032 37632 4032 37632 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 3120 13440 3120 13440 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 12240 41916 12240 41916 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit30.Q
rlabel metal3 13632 41412 13632 41412 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit31.Q
rlabel metal3 3888 8652 3888 8652 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
rlabel metal3 1728 12516 1728 12516 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 1536 12180 1536 12180 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 2880 10290 2880 10290 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit7.Q
rlabel metal3 14784 36120 14784 36120 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 16416 35238 16416 35238 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 15984 33852 15984 33852 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 14496 34314 14496 34314 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 19824 13188 19824 13188 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit10.Q
rlabel metal3 4752 30660 4752 30660 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit11.Q
rlabel metal3 6240 29820 6240 29820 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 6048 30030 6048 30030 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 1344 23898 1344 23898 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q
rlabel via2 3936 24609 3936 24609 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 2688 22554 2688 22554 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 13536 25326 13536 25326 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q
rlabel metal3 12528 24780 12528 24780 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 11616 25704 11616 25704 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 9072 32907 9072 32907 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 16992 9324 16992 9324 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 17184 10542 17184 10542 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit21.Q
rlabel metal3 18624 9660 18624 9660 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit22.Q
rlabel metal3 4560 29148 4560 29148 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 3072 28014 3072 28014 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit24.Q
rlabel metal3 3932 29064 3932 29064 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit25.Q
rlabel metal3 3168 21588 3168 21588 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q
rlabel via1 3072 22272 3072 22272 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 4512 21462 4512 21462 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 20256 21378 20256 21378 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 7488 32802 7488 32802 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit3.Q
rlabel metal3 19008 23100 19008 23100 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 20016 23100 20016 23100 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 11616 32594 11616 32594 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit4.Q
rlabel metal3 9984 32340 9984 32340 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 20400 32340 20400 32340 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit6.Q
rlabel metal3 18192 33852 18192 33852 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 18529 10072 18529 10072 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 20064 12597 20064 12597 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit9.Q
rlabel metal3 18816 26292 18816 26292 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 18096 23940 18096 23940 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 8304 27804 8304 27804 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 6816 28266 6816 28266 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 10656 31290 10656 31290 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 12240 31395 12240 31395 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 18720 30408 18720 30408 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit14.Q
rlabel metal3 16032 30828 16032 30828 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 15168 36750 15168 36750 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit16.Q
rlabel metal2 17568 36120 17568 36120 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 6384 39732 6384 39732 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit18.Q
rlabel metal3 7584 39060 7584 39060 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit19.Q
rlabel metal3 8928 26292 8928 26292 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit2.Q
rlabel metal3 5904 37632 5904 37632 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit20.Q
rlabel metal3 7488 37632 7488 37632 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 14688 39942 14688 39942 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 17232 39060 17232 39060 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 18240 33145 18240 33145 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 16944 31500 16944 31500 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 8736 29397 8736 29397 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit26.Q
rlabel metal3 7104 29148 7104 29148 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 9216 30909 9216 30909 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 7680 30912 7680 30912 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 7776 26754 7776 26754 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 16416 30954 16416 30954 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit30.Q
rlabel metal3 15024 31500 15024 31500 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 10176 26964 10176 26964 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit4.Q
rlabel metal2 11520 27090 11520 27090 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit5.Q
rlabel metal3 19584 29316 19584 29316 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 17664 29400 17664 29400 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 13248 32256 13248 32256 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit8.Q
rlabel via1 14832 32167 14832 32167 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit9.Q
rlabel via2 19200 17472 19200 17472 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q
rlabel metal2 19488 18144 19488 18144 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 9600 22554 9600 22554 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 9888 22470 9888 22470 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit11.Q
rlabel metal2 11616 23688 11616 23688 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q
rlabel metal2 9696 23478 9696 23478 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit13.Q
rlabel metal3 19056 19740 19056 19740 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q
rlabel metal3 17856 19908 17856 19908 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit15.Q
rlabel metal2 17184 32550 17184 32550 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit16.Q
rlabel metal2 19296 32130 19296 32130 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 9408 24311 9408 24311 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit18.Q
rlabel metal3 7680 23940 7680 23940 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit19.Q
rlabel metal3 10752 18564 10752 18564 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q
rlabel metal2 9888 28098 9888 28098 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit20.Q
rlabel metal2 11760 28560 11760 28560 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit21.Q
rlabel metal2 18864 23268 18864 23268 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit22.Q
rlabel metal3 17184 26292 17184 26292 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit23.Q
rlabel metal2 14256 29316 14256 29316 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit24.Q
rlabel metal3 15648 29484 15648 29484 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit25.Q
rlabel metal3 8064 24780 8064 24780 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 6960 25284 6960 25284 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit27.Q
rlabel metal2 10608 30072 10608 30072 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit28.Q
rlabel metal2 12480 30324 12480 30324 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 10656 19320 10656 19320 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit3.Q
rlabel metal3 19104 25578 19104 25578 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit30.Q
rlabel metal3 16224 29148 16224 29148 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit31.Q
rlabel metal3 13056 20076 13056 20076 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 13056 19488 13056 19488 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit5.Q
rlabel metal2 17280 21546 17280 21546 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q
rlabel metal3 16800 21588 16800 21588 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit7.Q
rlabel metal2 19104 21840 19104 21840 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 19872 21630 19872 21630 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 11808 34064 11808 34064 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 12672 35778 12672 35778 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 4128 30828 4128 30828 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit10.Q
rlabel metal3 2256 31332 2256 31332 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 3072 16632 3072 16632 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 2400 17556 2400 17556 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit13.Q
rlabel metal2 16560 17220 16560 17220 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit14.Q
rlabel metal2 14976 18648 14976 18648 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit15.Q
rlabel metal2 19392 15582 19392 15582 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 19104 15960 19104 15960 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 9408 17094 9408 17094 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q
rlabel metal2 9504 17808 9504 17808 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit19.Q
rlabel metal2 6528 23142 6528 23142 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 13200 16968 13200 16968 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q
rlabel metal2 13632 17556 13632 17556 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit21.Q
rlabel metal2 19200 7014 19200 7014 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q
rlabel via1 19298 7140 19298 7140 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit23.Q
rlabel metal3 19248 7728 19248 7728 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 19776 9198 19776 9198 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 8064 19866 8064 19866 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q
rlabel metal2 8208 20076 8208 20076 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 11616 20832 11616 20832 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q
rlabel metal2 11328 20118 11328 20118 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit29.Q
rlabel metal2 7968 22344 7968 22344 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q
rlabel metal2 19104 18606 19104 18606 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q
rlabel metal2 19680 19320 19680 19320 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit31.Q
rlabel metal2 6864 21000 6864 21000 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit4.Q
rlabel metal2 15984 24612 15984 24612 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q
rlabel metal2 17568 24903 17568 24903 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 17376 24192 17376 24192 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 14880 16716 14880 16716 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit8.Q
rlabel metal2 13056 17094 13056 17094 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit9.Q
rlabel metal3 4272 27468 4272 27468 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit0.Q
rlabel metal3 14304 25116 14304 25116 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q
rlabel metal2 12672 22302 12672 22302 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 14112 21672 14112 21672 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit11.Q
rlabel metal2 13200 14028 13200 14028 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit12.Q
rlabel metal2 14976 14319 14976 14319 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit13.Q
rlabel metal2 7584 17094 7584 17094 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit14.Q
rlabel metal2 9120 16751 9120 16751 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit15.Q
rlabel metal2 6912 15792 6912 15792 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit16.Q
rlabel metal3 8304 14952 8304 14952 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit17.Q
rlabel metal2 10848 12768 10848 12768 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 12336 11928 12336 11928 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit19.Q
rlabel metal2 13536 27006 13536 27006 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q
rlabel via1 12624 7975 12624 7975 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit20.Q
rlabel metal2 11040 8148 11040 8148 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit21.Q
rlabel metal2 9888 6888 9888 6888 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit22.Q
rlabel metal2 8256 7098 8256 7098 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit23.Q
rlabel metal2 10368 8400 10368 8400 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit24.Q
rlabel metal2 8688 8148 8688 8148 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit25.Q
rlabel metal2 14208 6890 14208 6890 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit26.Q
rlabel metal2 12672 7224 12672 7224 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 15792 14028 15792 14028 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q
rlabel metal2 17088 15372 17088 15372 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q
rlabel metal3 14256 28140 14256 28140 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit3.Q
rlabel metal3 17616 15708 17616 15708 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit30.Q
rlabel metal2 10272 34398 10272 34398 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q
rlabel metal2 13152 10332 13152 10332 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit4.Q
rlabel metal2 14832 10416 14832 10416 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit5.Q
rlabel metal2 5664 33096 5664 33096 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit6.Q
rlabel via1 7440 33679 7440 33679 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit7.Q
rlabel metal2 4560 19488 4560 19488 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit8.Q
rlabel metal3 6144 19488 6144 19488 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 14496 12938 14496 12938 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit0.Q
rlabel metal2 12960 13146 12960 13146 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit1.Q
rlabel metal3 7008 17724 7008 17724 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit10.Q
rlabel metal2 8640 18193 8640 18193 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit11.Q
rlabel metal3 3648 14196 3648 14196 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 5472 15239 5472 15239 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit13.Q
rlabel metal2 11328 11046 11328 11046 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 12864 10703 12864 10703 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit15.Q
rlabel metal2 10368 14994 10368 14994 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit16.Q
rlabel metal2 11424 14238 11424 14238 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit17.Q
rlabel metal3 6864 11928 6864 11928 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 9024 11970 9024 11970 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit19.Q
rlabel metal2 3456 33723 3456 33723 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit2.Q
rlabel metal2 6384 8904 6384 8904 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 8448 8904 8448 8904 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 14880 6510 14880 6510 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 16512 6678 16512 6678 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit23.Q
rlabel metal2 15696 11508 15696 11508 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q
rlabel metal2 17376 11634 17376 11634 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q
rlabel metal3 16896 11508 16896 11508 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit26.Q
rlabel metal2 5472 35112 5472 35112 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q
rlabel metal2 5952 34146 5952 34146 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q
rlabel metal3 5952 36540 5952 36540 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit29.Q
rlabel metal2 4368 32340 4368 32340 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit3.Q
rlabel metal2 1536 25998 1536 25998 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q
rlabel metal2 3312 23940 3312 23940 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q
rlabel metal3 4416 19908 4416 19908 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit4.Q
rlabel metal2 2736 18732 2736 18732 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit5.Q
rlabel metal2 14688 23349 14688 23349 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit6.Q
rlabel metal2 13152 23142 13152 23142 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit7.Q
rlabel metal2 13056 14448 13056 14448 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit8.Q
rlabel via1 15024 14704 15024 14704 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 19296 17052 19296 17052 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E1BEG0
rlabel metal2 4320 31332 4320 31332 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E1BEG1
rlabel metal2 3456 16170 3456 16170 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E1BEG2
rlabel metal2 16224 18228 16224 18228 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E1BEG3
rlabel metal3 18432 16296 18432 16296 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG0
rlabel metal2 11136 16926 11136 16926 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG1
rlabel metal3 14880 17808 14880 17808 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG2
rlabel metal2 20064 7476 20064 7476 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG3
rlabel metal2 20016 8736 20016 8736 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG4
rlabel metal2 16992 17220 16992 17220 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG5
rlabel metal3 12288 15036 12288 15036 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG6
rlabel metal3 20016 13272 20016 13272 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG7
rlabel metal2 15264 17010 15264 17010 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb0
rlabel metal3 12672 19614 12672 19614 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb1
rlabel metal3 16752 14784 16752 14784 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb2
rlabel metal3 17904 15456 17904 15456 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb3
rlabel metal4 19680 19908 19680 19908 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb4
rlabel metal2 20064 16716 20064 16716 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb5
rlabel metal2 11712 23310 11712 23310 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb6
rlabel metal3 19008 17640 19008 17640 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb7
rlabel metal2 19680 37380 19680 37380 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG0
rlabel metal2 19584 38976 19584 38976 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG1
rlabel metal3 18768 29904 18768 29904 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG10
rlabel metal2 19728 34440 19728 34440 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG11
rlabel metal3 13632 37464 13632 37464 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG2
rlabel metal2 20064 39438 20064 39438 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG3
rlabel metal2 19872 31668 19872 31668 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG4
rlabel metal2 19872 28014 19872 28014 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG5
rlabel metal2 19584 28602 19584 28602 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG6
rlabel metal2 17184 30408 17184 30408 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG7
rlabel metal2 19392 31458 19392 31458 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG8
rlabel metal2 17184 30996 17184 30996 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG9
rlabel metal2 20064 33348 20064 33348 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG0
rlabel metal2 16992 18144 16992 18144 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG1
rlabel metal2 15264 24612 15264 24612 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG10
rlabel metal2 19296 28392 19296 28392 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG11
rlabel metal2 20064 29106 20064 29106 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG12
rlabel metal2 8544 27510 8544 27510 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG13
rlabel metal2 16800 30870 16800 30870 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG14
rlabel metal3 19248 30408 19248 30408 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG15
rlabel metal2 12000 29694 12000 29694 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG2
rlabel metal2 19392 26334 19392 26334 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG3
rlabel metal2 16128 29652 16128 29652 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG4
rlabel metal2 16800 23562 16800 23562 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG5
rlabel metal2 12480 30744 12480 30744 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG6
rlabel metal3 17664 27552 17664 27552 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG7
rlabel metal2 16848 29904 16848 29904 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG8
rlabel metal3 16176 18816 16176 18816 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG9
rlabel metal2 16656 17976 16656 17976 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG12
rlabel metal2 10944 29316 10944 29316 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG13
rlabel metal5 3696 26292 3696 26292 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG14
rlabel metal2 18144 33432 18144 33432 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG15
rlabel metal3 9648 1176 9648 1176 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S1BEG0
rlabel metal3 7872 33768 7872 33768 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S1BEG1
rlabel metal2 7056 1176 7056 1176 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S1BEG2
rlabel metal3 12822 2436 12822 2436 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S1BEG3
rlabel metal3 15504 12684 15504 12684 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG0
rlabel metal2 9072 1848 9072 1848 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG1
rlabel metal2 8640 2184 8640 2184 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG2
rlabel metal2 12624 12600 12624 12600 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG3
rlabel metal2 11712 7224 11712 7224 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG4
rlabel metal2 10176 6678 10176 6678 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG5
rlabel metal3 10128 4116 10128 4116 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG6
rlabel metal3 13872 6972 13872 6972 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG7
rlabel metal3 16992 15288 16992 15288 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S4BEG0
rlabel metal3 12576 5040 12576 5040 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S4BEG1
rlabel metal4 14400 12096 14400 12096 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S4BEG2
rlabel metal3 16704 1848 16704 1848 0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S4BEG3
rlabel metal3 16224 48552 16224 48552 0 UIO_IN_TT_PROJECT0
rlabel metal3 1182 29484 1182 29484 0 UIO_IN_TT_PROJECT1
rlabel metal3 2766 30156 2766 30156 0 UIO_IN_TT_PROJECT2
rlabel metal3 606 30828 606 30828 0 UIO_IN_TT_PROJECT3
rlabel metal3 366 31500 366 31500 0 UIO_IN_TT_PROJECT4
rlabel metal3 1134 32172 1134 32172 0 UIO_IN_TT_PROJECT5
rlabel metal3 1326 32844 1326 32844 0 UIO_IN_TT_PROJECT6
rlabel metal3 654 33516 654 33516 0 UIO_IN_TT_PROJECT7
rlabel metal3 654 18060 654 18060 0 UIO_OE_TT_PROJECT0
rlabel metal3 654 18732 654 18732 0 UIO_OE_TT_PROJECT1
rlabel metal4 6816 68208 6816 68208 0 UIO_OE_TT_PROJECT2
rlabel metal3 174 20076 174 20076 0 UIO_OE_TT_PROJECT3
rlabel metal3 17520 65436 17520 65436 0 UIO_OE_TT_PROJECT4
rlabel metal3 654 21420 654 21420 0 UIO_OE_TT_PROJECT5
rlabel metal3 7488 64344 7488 64344 0 UIO_OE_TT_PROJECT6
rlabel metal2 11568 33348 11568 33348 0 UIO_OE_TT_PROJECT7
rlabel metal2 17088 59136 17088 59136 0 UIO_OUT_TT_PROJECT0
rlabel metal2 13728 59976 13728 59976 0 UIO_OUT_TT_PROJECT1
rlabel metal3 78 14028 78 14028 0 UIO_OUT_TT_PROJECT2
rlabel metal3 654 14700 654 14700 0 UIO_OUT_TT_PROJECT3
rlabel metal3 126 15372 126 15372 0 UIO_OUT_TT_PROJECT4
rlabel metal3 2094 16044 2094 16044 0 UIO_OUT_TT_PROJECT5
rlabel metal3 510 16716 510 16716 0 UIO_OUT_TT_PROJECT6
rlabel metal3 126 17388 126 17388 0 UIO_OUT_TT_PROJECT7
rlabel metal3 126 23436 126 23436 0 UI_IN_TT_PROJECT0
rlabel metal3 78 24108 78 24108 0 UI_IN_TT_PROJECT1
rlabel metal2 3072 24402 3072 24402 0 UI_IN_TT_PROJECT2
rlabel metal2 12480 25662 12480 25662 0 UI_IN_TT_PROJECT3
rlabel metal3 960 10752 960 10752 0 UI_IN_TT_PROJECT4
rlabel metal3 654 26796 654 26796 0 UI_IN_TT_PROJECT5
rlabel metal2 3936 22092 3936 22092 0 UI_IN_TT_PROJECT6
rlabel metal3 654 28140 654 28140 0 UI_IN_TT_PROJECT7
rlabel via3 78 7308 78 7308 0 UO_OUT_TT_PROJECT0
rlabel metal3 1278 7980 1278 7980 0 UO_OUT_TT_PROJECT1
rlabel metal3 222 8652 222 8652 0 UO_OUT_TT_PROJECT2
rlabel metal3 17568 35868 17568 35868 0 UO_OUT_TT_PROJECT3
rlabel metal3 78 9996 78 9996 0 UO_OUT_TT_PROJECT4
rlabel metal3 798 10668 798 10668 0 UO_OUT_TT_PROJECT5
rlabel metal3 270 11340 270 11340 0 UO_OUT_TT_PROJECT6
rlabel metal3 654 12012 654 12012 0 UO_OUT_TT_PROJECT7
rlabel metal2 16608 13734 16608 13734 0 _0000_
rlabel metal2 8352 12138 8352 12138 0 _0001_
rlabel metal2 12096 20916 12096 20916 0 _0002_
rlabel metal2 17184 18480 17184 18480 0 _0003_
rlabel metal3 12816 52332 12816 52332 0 _0004_
rlabel metal2 13248 52710 13248 52710 0 _0005_
rlabel metal2 13632 49602 13632 49602 0 _0006_
rlabel metal2 13632 16842 13632 16842 0 _0007_
rlabel metal2 14400 9744 14400 9744 0 _0008_
rlabel metal3 14016 9492 14016 9492 0 _0009_
rlabel metal2 14400 11109 14400 11109 0 _0010_
rlabel metal2 17568 54810 17568 54810 0 _0011_
rlabel metal3 7392 54180 7392 54180 0 _0012_
rlabel metal3 7680 53592 7680 53592 0 _0013_
rlabel metal2 16272 54180 16272 54180 0 _0014_
rlabel metal2 17472 48552 17472 48552 0 _0015_
rlabel metal2 17376 49056 17376 49056 0 _0016_
rlabel metal2 15744 49980 15744 49980 0 _0017_
rlabel metal3 17184 50988 17184 50988 0 _0018_
rlabel metal2 15072 49518 15072 49518 0 _0019_
rlabel metal2 17232 48972 17232 48972 0 _0020_
rlabel metal3 16224 49476 16224 49476 0 _0021_
rlabel metal2 7296 47880 7296 47880 0 _0022_
rlabel metal2 7776 49140 7776 49140 0 _0023_
rlabel metal3 7248 50400 7248 50400 0 _0024_
rlabel metal3 6672 51828 6672 51828 0 _0025_
rlabel metal3 7392 49476 7392 49476 0 _0026_
rlabel metal2 7680 48846 7680 48846 0 _0027_
rlabel metal3 7968 48636 7968 48636 0 _0028_
rlabel metal2 7632 56532 7632 56532 0 _0029_
rlabel metal2 8256 55776 8256 55776 0 _0030_
rlabel metal2 8496 55524 8496 55524 0 _0031_
rlabel metal2 8736 56448 8736 56448 0 _0032_
rlabel metal3 8400 56196 8400 56196 0 _0033_
rlabel metal2 7968 55776 7968 55776 0 _0034_
rlabel metal2 8880 56196 8880 56196 0 _0035_
rlabel metal2 17760 57792 17760 57792 0 _0036_
rlabel metal3 18480 57876 18480 57876 0 _0037_
rlabel metal3 19632 57036 19632 57036 0 _0038_
rlabel metal2 18768 57624 18768 57624 0 _0039_
rlabel metal2 17952 57120 17952 57120 0 _0040_
rlabel metal2 19680 56826 19680 56826 0 _0041_
rlabel metal2 18144 57162 18144 57162 0 _0042_
rlabel metal3 13920 43428 13920 43428 0 _0043_
rlabel metal2 13440 43512 13440 43512 0 _0044_
rlabel metal3 13104 44268 13104 44268 0 _0045_
rlabel metal2 16800 43302 16800 43302 0 _0046_
rlabel metal2 13632 43932 13632 43932 0 _0047_
rlabel metal2 14304 43344 14304 43344 0 _0048_
rlabel metal3 15648 43260 15648 43260 0 _0049_
rlabel metal2 15456 44604 15456 44604 0 _0050_
rlabel metal3 15984 43428 15984 43428 0 _0051_
rlabel metal2 6432 47040 6432 47040 0 _0052_
rlabel metal3 6816 46452 6816 46452 0 _0053_
rlabel metal2 8160 45024 8160 45024 0 _0054_
rlabel metal3 8016 44940 8016 44940 0 _0055_
rlabel metal2 6720 46578 6720 46578 0 _0056_
rlabel metal2 7392 44856 7392 44856 0 _0057_
rlabel metal2 7584 44940 7584 44940 0 _0058_
rlabel metal2 7584 45822 7584 45822 0 _0059_
rlabel metal2 8016 44940 8016 44940 0 _0060_
rlabel metal3 9744 52500 9744 52500 0 _0061_
rlabel metal3 10464 52332 10464 52332 0 _0062_
rlabel metal2 10464 52290 10464 52290 0 _0063_
rlabel metal2 10944 53592 10944 53592 0 _0064_
rlabel metal2 8064 53172 8064 53172 0 _0065_
rlabel metal2 11424 53802 11424 53802 0 _0066_
rlabel metal3 10512 53340 10512 53340 0 _0067_
rlabel metal2 11616 53172 11616 53172 0 _0068_
rlabel metal2 11712 52962 11712 52962 0 _0069_
rlabel metal2 17568 56070 17568 56070 0 _0070_
rlabel metal3 16464 53340 16464 53340 0 _0071_
rlabel metal2 15936 51870 15936 51870 0 _0072_
rlabel metal2 15840 52458 15840 52458 0 _0073_
rlabel metal2 17952 55104 17952 55104 0 _0074_
rlabel metal2 17472 54894 17472 54894 0 _0075_
rlabel metal2 17184 54852 17184 54852 0 _0076_
rlabel metal2 15360 53970 15360 53970 0 _0077_
rlabel metal3 15984 54180 15984 54180 0 _0078_
rlabel metal2 19872 50211 19872 50211 0 _0079_
rlabel metal2 20160 48888 20160 48888 0 _0080_
rlabel metal2 17904 48972 17904 48972 0 _0081_
rlabel metal2 19872 48888 19872 48888 0 _0082_
rlabel metal3 3456 48888 3456 48888 0 _0083_
rlabel metal2 2784 47796 2784 47796 0 _0084_
rlabel metal2 3072 48468 3072 48468 0 _0085_
rlabel metal2 2496 47544 2496 47544 0 _0086_
rlabel metal2 6336 53130 6336 53130 0 _0087_
rlabel metal2 5664 51996 5664 51996 0 _0088_
rlabel metal2 6048 52968 6048 52968 0 _0089_
rlabel metal2 5952 52080 5952 52080 0 _0090_
rlabel metal3 19776 52878 19776 52878 0 _0091_
rlabel metal2 19968 53130 19968 53130 0 _0092_
rlabel metal2 16704 52710 16704 52710 0 _0093_
rlabel metal2 16608 52542 16608 52542 0 _0094_
rlabel metal2 18048 45654 18048 45654 0 _0095_
rlabel metal2 17952 46032 17952 46032 0 _0096_
rlabel metal2 17424 44268 17424 44268 0 _0097_
rlabel metal3 17040 44268 17040 44268 0 _0098_
rlabel metal2 16752 44100 16752 44100 0 _0099_
rlabel metal2 4512 45864 4512 45864 0 _0100_
rlabel metal3 4416 44940 4416 44940 0 _0101_
rlabel metal2 4704 45402 4704 45402 0 _0102_
rlabel metal2 4416 44852 4416 44852 0 _0103_
rlabel metal2 4224 45108 4224 45108 0 _0104_
rlabel metal2 3552 51534 3552 51534 0 _0105_
rlabel metal2 3840 51114 3840 51114 0 _0106_
rlabel metal2 3072 52248 3072 52248 0 _0107_
rlabel metal2 3120 50988 3120 50988 0 _0108_
rlabel metal2 3072 51450 3072 51450 0 _0109_
rlabel metal2 17568 52584 17568 52584 0 _0110_
rlabel metal2 17664 52626 17664 52626 0 _0111_
rlabel metal2 18433 51919 18433 51919 0 _0112_
rlabel metal2 18096 50988 18096 50988 0 _0113_
rlabel metal3 17760 51156 17760 51156 0 _0114_
rlabel metal3 19680 16044 19680 16044 0 _0115_
rlabel metal2 19008 16086 19008 16086 0 _0116_
rlabel metal3 10464 17724 10464 17724 0 _0117_
rlabel metal2 10656 17682 10656 17682 0 _0118_
rlabel metal2 13152 16212 13152 16212 0 _0119_
rlabel metal2 13632 17808 13632 17808 0 _0120_
rlabel metal3 19536 8652 19536 8652 0 _0121_
rlabel metal2 19296 7980 19296 7980 0 _0122_
rlabel metal4 19584 8232 19584 8232 0 _0123_
rlabel metal2 19968 8358 19968 8358 0 _0124_
rlabel metal2 9408 20076 9408 20076 0 _0125_
rlabel metal2 8352 20034 8352 20034 0 _0126_
rlabel metal2 11904 20580 11904 20580 0 _0127_
rlabel metal2 11520 20286 11520 20286 0 _0128_
rlabel metal2 19392 19425 19392 19425 0 _0129_
rlabel metal2 19776 19740 19776 19740 0 _0130_
rlabel metal3 19680 17724 19680 17724 0 _0131_
rlabel metal2 19584 18060 19584 18060 0 _0132_
rlabel metal2 10848 18984 10848 18984 0 _0133_
rlabel metal2 10464 18564 10464 18564 0 _0134_
rlabel metal3 14016 19068 14016 19068 0 _0135_
rlabel metal3 13152 20916 13152 20916 0 _0136_
rlabel metal3 15696 20580 15696 20580 0 _0137_
rlabel metal2 17136 21420 17136 21420 0 _0138_
rlabel metal2 19344 21756 19344 21756 0 _0139_
rlabel metal2 19824 21420 19824 21420 0 _0140_
rlabel metal2 10080 22008 10080 22008 0 _0141_
rlabel metal2 9792 22386 9792 22386 0 _0142_
rlabel metal2 11520 23604 11520 23604 0 _0143_
rlabel metal3 10272 23268 10272 23268 0 _0144_
rlabel metal3 17616 19992 17616 19992 0 _0145_
rlabel metal3 19296 20076 19296 20076 0 _0146_
rlabel metal2 15936 37548 15936 37548 0 _0147_
rlabel metal2 7392 31920 7392 31920 0 _0148_
rlabel metal3 7680 35280 7680 35280 0 _0149_
rlabel metal2 15648 14448 15648 14448 0 _0150_
rlabel metal2 18624 27594 18624 27594 0 _0151_
rlabel metal2 7968 32802 7968 32802 0 _0152_
rlabel metal2 4464 35364 4464 35364 0 _0153_
rlabel metal2 15552 13650 15552 13650 0 _0154_
rlabel metal3 15360 26124 15360 26124 0 _0155_
rlabel metal2 1632 24948 1632 24948 0 _0156_
rlabel metal2 10656 33558 10656 33558 0 _0157_
rlabel metal2 16896 14868 16896 14868 0 _0158_
rlabel metal2 17760 11928 17760 11928 0 _0159_
rlabel metal3 16464 12516 16464 12516 0 _0160_
rlabel metal2 17088 11130 17088 11130 0 _0161_
rlabel metal3 17472 11172 17472 11172 0 _0162_
rlabel metal3 16416 11928 16416 11928 0 _0163_
rlabel metal2 15408 12600 15408 12600 0 _0164_
rlabel metal2 15216 12516 15216 12516 0 _0165_
rlabel metal2 7872 33558 7872 33558 0 _0166_
rlabel metal3 7584 32340 7584 32340 0 _0167_
rlabel metal2 5328 33852 5328 33852 0 _0168_
rlabel metal2 5136 35196 5136 35196 0 _0169_
rlabel metal2 6864 35532 6864 35532 0 _0170_
rlabel metal3 7872 38220 7872 38220 0 _0171_
rlabel metal2 7248 35868 7248 35868 0 _0172_
rlabel metal2 5952 25788 5952 25788 0 _0173_
rlabel metal2 6144 25158 6144 25158 0 _0174_
rlabel metal2 2112 24444 2112 24444 0 _0175_
rlabel metal3 5136 23940 5136 23940 0 _0176_
rlabel metal3 6000 27048 6000 27048 0 _0177_
rlabel metal3 3840 27636 3840 27636 0 _0178_
rlabel metal2 6624 27510 6624 27510 0 _0179_
rlabel metal3 15024 26796 15024 26796 0 _0180_
rlabel metal3 14448 29064 14448 29064 0 _0181_
rlabel metal2 13824 25074 13824 25074 0 _0182_
rlabel metal2 16608 28014 16608 28014 0 _0183_
rlabel metal3 12960 29820 12960 29820 0 _0184_
rlabel metal2 15936 27552 15936 27552 0 _0185_
rlabel metal2 15984 29400 15984 29400 0 _0186_
rlabel metal2 17856 13944 17856 13944 0 _0187_
rlabel metal2 18000 14196 18000 14196 0 _0188_
rlabel metal2 16992 14070 16992 14070 0 _0189_
rlabel metal2 17232 14952 17232 14952 0 _0190_
rlabel metal2 17568 14280 17568 14280 0 _0191_
rlabel metal3 17808 15540 17808 15540 0 _0192_
rlabel metal3 12192 33978 12192 33978 0 _0193_
rlabel metal2 12288 34188 12288 34188 0 _0194_
rlabel metal2 11520 35994 11520 35994 0 _0195_
rlabel metal2 12192 34650 12192 34650 0 _0196_
rlabel metal2 12480 35784 12480 35784 0 _0197_
rlabel metal2 12528 34356 12528 34356 0 _0198_
rlabel metal3 7536 22260 7536 22260 0 _0199_
rlabel metal2 7680 22596 7680 22596 0 _0200_
rlabel metal2 8256 22260 8256 22260 0 _0201_
rlabel metal2 7776 23016 7776 23016 0 _0202_
rlabel metal2 5472 22218 5472 22218 0 _0203_
rlabel metal3 6384 22428 6384 22428 0 _0204_
rlabel metal2 19008 26292 19008 26292 0 _0205_
rlabel metal2 16080 23100 16080 23100 0 _0206_
rlabel metal2 18240 23772 18240 23772 0 _0207_
rlabel metal2 15936 23310 15936 23310 0 _0208_
rlabel metal2 17760 24234 17760 24234 0 _0209_
rlabel metal3 16944 23100 16944 23100 0 _0210_
rlabel metal2 19728 13356 19728 13356 0 _0211_
rlabel metal2 18336 10374 18336 10374 0 _0212_
rlabel metal3 19488 12684 19488 12684 0 _0213_
rlabel metal2 19392 13860 19392 13860 0 _0214_
rlabel metal2 5952 30660 5952 30660 0 _0215_
rlabel metal2 6240 30114 6240 30114 0 _0216_
rlabel metal2 6528 30282 6528 30282 0 _0217_
rlabel metal3 6768 30072 6768 30072 0 _0218_
rlabel metal2 1440 25116 1440 25116 0 _0219_
rlabel metal2 1488 24780 1488 24780 0 _0220_
rlabel metal3 3792 23772 3792 23772 0 _0221_
rlabel metal2 1920 24402 1920 24402 0 _0222_
rlabel metal2 13440 24864 13440 24864 0 _0223_
rlabel metal3 14016 24612 14016 24612 0 _0224_
rlabel metal3 12336 26124 12336 26124 0 _0225_
rlabel metal2 12768 25914 12768 25914 0 _0226_
rlabel metal3 19584 8022 19584 8022 0 _0227_
rlabel metal2 17376 10584 17376 10584 0 _0228_
rlabel metal2 17760 11004 17760 11004 0 _0229_
rlabel metal2 17184 8652 17184 8652 0 _0230_
rlabel metal2 17760 10332 17760 10332 0 _0231_
rlabel metal2 4656 29148 4656 29148 0 _0232_
rlabel metal2 1344 26880 1344 26880 0 _0233_
rlabel metal3 1776 27888 1776 27888 0 _0234_
rlabel metal3 4368 29316 4368 29316 0 _0235_
rlabel metal2 1440 28224 1440 28224 0 _0236_
rlabel metal3 4464 21756 4464 21756 0 _0237_
rlabel metal2 3552 22764 3552 22764 0 _0238_
rlabel metal2 4128 21798 4128 21798 0 _0239_
rlabel metal2 5328 23772 5328 23772 0 _0240_
rlabel metal2 5376 23058 5376 23058 0 _0241_
rlabel metal2 20256 24318 20256 24318 0 _0242_
rlabel metal2 19872 25788 19872 25788 0 _0243_
rlabel metal2 20064 25746 20064 25746 0 _0244_
rlabel metal3 19776 25116 19776 25116 0 _0245_
rlabel metal2 19584 25452 19584 25452 0 _0246_
rlabel metal2 6000 12516 6000 12516 0 _0247_
rlabel metal2 6864 11928 6864 11928 0 _0248_
rlabel metal3 5712 12348 5712 12348 0 _0249_
rlabel metal2 3600 11676 3600 11676 0 _0250_
rlabel metal3 4272 11844 4272 11844 0 _0251_
rlabel metal2 7104 13140 7104 13140 0 _0252_
rlabel metal2 7200 13818 7200 13818 0 _0253_
rlabel metal3 4800 12516 4800 12516 0 _0254_
rlabel metal3 4800 14028 4800 14028 0 _0255_
rlabel metal2 3456 12432 3456 12432 0 _0256_
rlabel metal2 3648 12894 3648 12894 0 _0257_
rlabel metal2 4128 13902 4128 13902 0 _0258_
rlabel metal2 4224 12768 4224 12768 0 _0259_
rlabel metal3 3696 11676 3696 11676 0 _0260_
rlabel metal2 4320 11970 4320 11970 0 _0261_
rlabel metal2 3648 14154 3648 14154 0 _0262_
rlabel metal2 3936 12558 3936 12558 0 _0263_
rlabel metal5 3648 12516 3648 12516 0 _0264_
rlabel metal2 5568 9996 5568 9996 0 _0265_
rlabel metal3 5376 10164 5376 10164 0 _0266_
rlabel metal2 4512 8862 4512 8862 0 _0267_
rlabel metal2 4224 9156 4224 9156 0 _0268_
rlabel metal3 4464 8904 4464 8904 0 _0269_
rlabel metal2 7008 9954 7008 9954 0 _0270_
rlabel metal2 5664 10248 5664 10248 0 _0271_
rlabel metal2 6048 9618 6048 9618 0 _0272_
rlabel metal2 6000 9324 6000 9324 0 _0273_
rlabel metal2 5616 11004 5616 11004 0 _0274_
rlabel metal2 5376 10290 5376 10290 0 _0275_
rlabel metal2 5088 9576 5088 9576 0 _0276_
rlabel metal3 5184 9534 5184 9534 0 _0277_
rlabel metal3 5088 8148 5088 8148 0 _0278_
rlabel metal2 4656 7812 4656 7812 0 _0279_
rlabel metal2 4224 8232 4224 8232 0 _0280_
rlabel metal3 3744 8148 3744 8148 0 _0281_
rlabel metal2 1440 12012 1440 12012 0 _0282_
rlabel metal3 3264 7980 3264 7980 0 _0283_
rlabel metal2 1536 11550 1536 11550 0 _0284_
rlabel metal3 2352 11508 2352 11508 0 _0285_
rlabel metal2 3696 8148 3696 8148 0 _0286_
rlabel metal2 3312 55776 3312 55776 0 _0287_
rlabel metal2 5232 56532 5232 56532 0 _0288_
rlabel metal2 15648 58002 15648 58002 0 _0289_
rlabel metal3 13920 52500 13920 52500 0 _0290_
rlabel metal3 19776 50316 19776 50316 0 _0291_
rlabel metal2 3264 49434 3264 49434 0 _0292_
rlabel metal3 5952 51996 5952 51996 0 _0293_
rlabel metal2 20064 53508 20064 53508 0 _0294_
rlabel metal2 3264 8148 3264 8148 0 _0295_
rlabel metal2 4800 10458 4800 10458 0 _0296_
rlabel metal3 15072 21588 15072 21588 0 _0297_
rlabel metal2 3360 17010 3360 17010 0 _0298_
rlabel metal2 4896 32340 4896 32340 0 _0299_
rlabel metal3 15024 8820 15024 8820 0 _0300_
rlabel metal2 17376 14700 17376 14700 0 _0301_
rlabel metal3 11232 35196 11232 35196 0 _0302_
rlabel metal2 7296 20790 7296 20790 0 _0303_
rlabel metal2 17952 24570 17952 24570 0 _0304_
rlabel metal3 5328 13944 5328 13944 0 _0305_
rlabel metal3 3456 11802 3456 11802 0 _0306_
rlabel metal2 3792 8064 3792 8064 0 _0307_
rlabel metal3 3744 55608 3744 55608 0 _0308_
rlabel metal2 3216 55020 3216 55020 0 _0309_
rlabel metal2 3408 49476 3408 49476 0 _0310_
rlabel metal2 4272 35448 4272 35448 0 _0311_
rlabel metal3 3360 32844 3360 32844 0 _0312_
rlabel metal2 4464 32004 4464 32004 0 _0313_
rlabel metal3 5424 33684 5424 33684 0 _0314_
rlabel metal3 4512 57876 4512 57876 0 _0315_
rlabel metal2 3648 57750 3648 57750 0 _0316_
rlabel metal2 4176 54012 4176 54012 0 _0317_
rlabel metal3 2880 17808 2880 17808 0 _0318_
rlabel metal2 3936 16212 3936 16212 0 _0319_
rlabel metal3 4128 17052 4128 17052 0 _0320_
rlabel metal3 3792 19824 3792 19824 0 _0321_
rlabel metal2 15744 59254 15744 59254 0 _0322_
rlabel metal2 15648 59556 15648 59556 0 _0323_
rlabel metal2 14784 57624 14784 57624 0 _0324_
rlabel metal2 14016 29484 14016 29484 0 _0325_
rlabel metal2 14592 21714 14592 21714 0 _0326_
rlabel metal2 14496 21840 14496 21840 0 _0327_
rlabel metal2 13728 22092 13728 22092 0 _0328_
rlabel metal3 9408 14700 9408 14700 0 _0329_
rlabel metal2 10080 13608 10080 13608 0 _0330_
rlabel metal3 7680 13020 7680 13020 0 _0331_
rlabel metal3 9264 13188 9264 13188 0 _0332_
rlabel metal2 8160 12978 8160 12978 0 _0333_
rlabel metal3 14880 12012 14880 12012 0 _0334_
rlabel metal2 14448 14700 14448 14700 0 _0335_
rlabel metal3 11040 35868 11040 35868 0 _0336_
rlabel metal2 12096 35406 12096 35406 0 _0337_
rlabel metal2 9600 37128 9600 37128 0 _0338_
rlabel metal2 9696 37590 9696 37590 0 _0339_
rlabel metal2 9600 34398 9600 34398 0 _0340_
rlabel metal2 9792 33936 9792 33936 0 _0341_
rlabel metal2 11712 30576 11712 30576 0 _0342_
rlabel metal2 5232 18564 5232 18564 0 _0343_
rlabel metal2 5664 18606 5664 18606 0 _0344_
rlabel metal3 2112 17745 2112 17745 0 _0345_
rlabel metal2 1824 18018 1824 18018 0 _0346_
rlabel metal2 2112 18228 2112 18228 0 _0347_
rlabel metal2 6144 19320 6144 19320 0 _0348_
rlabel metal3 6672 18396 6672 18396 0 _0349_
rlabel metal2 11040 10248 11040 10248 0 _0350_
rlabel metal2 10704 11676 10704 11676 0 _0351_
rlabel metal2 9888 11424 9888 11424 0 _0352_
rlabel metal2 9504 10458 9504 10458 0 _0353_
rlabel metal3 9792 10038 9792 10038 0 _0354_
rlabel metal2 19837 8701 19837 8701 0 _0355_
rlabel metal2 11952 12516 11952 12516 0 _0356_
rlabel metal3 8304 51660 8304 51660 0 clknet_0_Tile_X0Y1_UserCLK
rlabel metal2 2112 36414 2112 36414 0 clknet_1_0__leaf_Tile_X0Y1_UserCLK
rlabel metal2 15360 82698 15360 82698 0 clknet_1_1__leaf_Tile_X0Y1_UserCLK
<< properties >>
string FIXED_BBOX 0 0 21504 86016
<< end >>
