module S_IO (A_I_top,
    A_O_top,
    A_T_top,
    A_config_C_bit0,
    A_config_C_bit1,
    A_config_C_bit2,
    A_config_C_bit3,
    B_I_top,
    B_O_top,
    B_T_top,
    B_config_C_bit0,
    B_config_C_bit1,
    B_config_C_bit2,
    B_config_C_bit3,
    Co,
    UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 output A_I_top;
 input A_O_top;
 output A_T_top;
 output A_config_C_bit0;
 output A_config_C_bit1;
 output A_config_C_bit2;
 output A_config_C_bit3;
 output B_I_top;
 input B_O_top;
 output B_T_top;
 output B_config_C_bit0;
 output B_config_C_bit1;
 output B_config_C_bit2;
 output B_config_C_bit3;
 output Co;
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire \Inst_A_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_S_IO_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_S_IO_switch_matrix.N1BEG0 ;
 wire \Inst_S_IO_switch_matrix.N1BEG1 ;
 wire \Inst_S_IO_switch_matrix.N1BEG2 ;
 wire \Inst_S_IO_switch_matrix.N1BEG3 ;
 wire \Inst_S_IO_switch_matrix.N2BEG0 ;
 wire \Inst_S_IO_switch_matrix.N2BEG1 ;
 wire \Inst_S_IO_switch_matrix.N2BEG2 ;
 wire \Inst_S_IO_switch_matrix.N2BEG3 ;
 wire \Inst_S_IO_switch_matrix.N2BEG4 ;
 wire \Inst_S_IO_switch_matrix.N2BEG5 ;
 wire \Inst_S_IO_switch_matrix.N2BEG6 ;
 wire \Inst_S_IO_switch_matrix.N2BEG7 ;
 wire \Inst_S_IO_switch_matrix.N2BEGb0 ;
 wire \Inst_S_IO_switch_matrix.N2BEGb1 ;
 wire \Inst_S_IO_switch_matrix.N2BEGb2 ;
 wire \Inst_S_IO_switch_matrix.N2BEGb3 ;
 wire \Inst_S_IO_switch_matrix.N2BEGb4 ;
 wire \Inst_S_IO_switch_matrix.N2BEGb5 ;
 wire \Inst_S_IO_switch_matrix.N2BEGb6 ;
 wire \Inst_S_IO_switch_matrix.N2BEGb7 ;
 wire \Inst_S_IO_switch_matrix.N4BEG0 ;
 wire \Inst_S_IO_switch_matrix.N4BEG1 ;
 wire \Inst_S_IO_switch_matrix.N4BEG10 ;
 wire \Inst_S_IO_switch_matrix.N4BEG11 ;
 wire \Inst_S_IO_switch_matrix.N4BEG12 ;
 wire \Inst_S_IO_switch_matrix.N4BEG13 ;
 wire \Inst_S_IO_switch_matrix.N4BEG14 ;
 wire \Inst_S_IO_switch_matrix.N4BEG15 ;
 wire \Inst_S_IO_switch_matrix.N4BEG2 ;
 wire \Inst_S_IO_switch_matrix.N4BEG3 ;
 wire \Inst_S_IO_switch_matrix.N4BEG4 ;
 wire \Inst_S_IO_switch_matrix.N4BEG5 ;
 wire \Inst_S_IO_switch_matrix.N4BEG6 ;
 wire \Inst_S_IO_switch_matrix.N4BEG7 ;
 wire \Inst_S_IO_switch_matrix.N4BEG8 ;
 wire \Inst_S_IO_switch_matrix.N4BEG9 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG0 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG1 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG10 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG11 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG12 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG13 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG14 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG15 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG2 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG3 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG4 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG5 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG6 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG7 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG8 ;
 wire \Inst_S_IO_switch_matrix.NN4BEG9 ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_1_0__leaf_UserCLK_regs;
 wire clknet_1_1__leaf_UserCLK_regs;
 wire [0:0] \Inst_S_IO_switch_matrix.DEBUG_select_N1BEG0 ;
 wire [0:0] \Inst_S_IO_switch_matrix.DEBUG_select_N1BEG1 ;
 wire [0:0] \Inst_S_IO_switch_matrix.DEBUG_select_N1BEG2 ;
 wire [0:0] \Inst_S_IO_switch_matrix.DEBUG_select_N1BEG3 ;

 sg13g2_mux4_1 _047_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(S1END[2]),
    .A1(S4END[15]),
    .A2(SS4END[15]),
    .A3(A_O_top),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit19.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG0 ));
 sg13g2_mux4_1 _048_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit16.Q ),
    .A0(S2END[0]),
    .A1(S4END[0]),
    .A2(SS4END[0]),
    .A3(SS4END[8]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit17.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEGb7 ));
 sg13g2_mux4_1 _049_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(S2END[1]),
    .A1(S4END[1]),
    .A2(SS4END[1]),
    .A3(SS4END[9]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit15.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEGb6 ));
 sg13g2_mux4_1 _050_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(S2END[2]),
    .A1(S4END[2]),
    .A2(SS4END[2]),
    .A3(SS4END[10]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit13.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEGb5 ));
 sg13g2_mux4_1 _051_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit10.Q ),
    .A0(S2END[3]),
    .A1(S4END[3]),
    .A2(SS4END[3]),
    .A3(SS4END[11]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit11.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEGb4 ));
 sg13g2_mux4_1 _052_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(S2END[4]),
    .A1(S4END[4]),
    .A2(SS4END[4]),
    .A3(SS4END[12]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit9.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEGb3 ));
 sg13g2_mux4_1 _053_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(S2END[5]),
    .A1(S4END[5]),
    .A2(SS4END[5]),
    .A3(SS4END[13]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit7.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEGb2 ));
 sg13g2_mux4_1 _054_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(S2END[6]),
    .A1(S4END[6]),
    .A2(SS4END[6]),
    .A3(SS4END[14]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit5.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEGb1 ));
 sg13g2_mux4_1 _055_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(S2END[7]),
    .A1(S4END[7]),
    .A2(SS4END[7]),
    .A3(SS4END[15]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit3.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEGb0 ));
 sg13g2_mux4_1 _056_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(S2MID[0]),
    .A1(S4END[0]),
    .A2(SS4END[0]),
    .A3(SS4END[8]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit1.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEG7 ));
 sg13g2_mux4_1 _057_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame3_bit30.Q ),
    .A0(S2MID[1]),
    .A1(S4END[1]),
    .A2(SS4END[1]),
    .A3(SS4END[9]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame3_bit31.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEG6 ));
 sg13g2_mux4_1 _058_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(S2MID[2]),
    .A1(S4END[2]),
    .A2(SS4END[2]),
    .A3(SS4END[10]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame3_bit29.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEG5 ));
 sg13g2_mux4_1 _059_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame3_bit26.Q ),
    .A0(S2MID[3]),
    .A1(S4END[3]),
    .A2(SS4END[3]),
    .A3(SS4END[11]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame3_bit27.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEG4 ));
 sg13g2_mux4_1 _060_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame3_bit24.Q ),
    .A0(S2MID[4]),
    .A1(S4END[4]),
    .A2(SS4END[4]),
    .A3(SS4END[12]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame3_bit25.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEG3 ));
 sg13g2_mux4_1 _061_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(S2MID[5]),
    .A1(S4END[5]),
    .A2(SS4END[5]),
    .A3(SS4END[13]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame3_bit23.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEG2 ));
 sg13g2_mux4_1 _062_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(S2MID[6]),
    .A1(S4END[6]),
    .A2(SS4END[6]),
    .A3(SS4END[14]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame3_bit21.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEG1 ));
 sg13g2_mux4_1 _063_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(S2MID[7]),
    .A1(S4END[7]),
    .A2(SS4END[7]),
    .A3(SS4END[15]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame3_bit19.Q ),
    .X(\Inst_S_IO_switch_matrix.N2BEG0 ));
 sg13g2_mux2_1 _064_ (.A0(S1END[0]),
    .A1(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_S_IO_switch_matrix.DEBUG_select_N1BEG3 [0]),
    .X(\Inst_S_IO_switch_matrix.N1BEG3 ));
 sg13g2_mux2_1 _065_ (.A0(S1END[1]),
    .A1(B_O_top),
    .S(\Inst_S_IO_switch_matrix.DEBUG_select_N1BEG2 [0]),
    .X(\Inst_S_IO_switch_matrix.N1BEG2 ));
 sg13g2_mux2_1 _066_ (.A0(S1END[2]),
    .A1(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_S_IO_switch_matrix.DEBUG_select_N1BEG1 [0]),
    .X(\Inst_S_IO_switch_matrix.N1BEG1 ));
 sg13g2_mux2_1 _067_ (.A0(S1END[3]),
    .A1(A_O_top),
    .S(\Inst_S_IO_switch_matrix.DEBUG_select_N1BEG0 [0]),
    .X(\Inst_S_IO_switch_matrix.N1BEG0 ));
 sg13g2_nand2b_1 _068_ (.Y(_032_),
    .B(\Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .A_N(S2END[3]));
 sg13g2_o21ai_1 _069_ (.B1(_032_),
    .Y(_033_),
    .A1(S2MID[7]),
    .A2(\Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nand3_1 _070_ (.B(\Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .C(_001_),
    .A(S2END[1]),
    .Y(_034_));
 sg13g2_o21ai_1 _071_ (.B1(_034_),
    .Y(_035_),
    .A1(\Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(_033_));
 sg13g2_nand3b_1 _072_ (.B(_001_),
    .C(S2END[0]),
    .Y(_036_),
    .A_N(\Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_o21ai_1 _073_ (.B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .Y(_037_),
    .A1(S2END[2]),
    .A2(\Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nand2_1 _074_ (.Y(_038_),
    .A(S2END[4]),
    .B(\Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nand4_1 _075_ (.B(_036_),
    .C(_037_),
    .A(\Inst_S_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .Y(_039_),
    .D(_038_));
 sg13g2_o21ai_1 _076_ (.B1(_039_),
    .Y(A_T_top),
    .A1(\Inst_S_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .A2(_035_));
 sg13g2_nand2b_1 _077_ (.Y(_040_),
    .B(S2END[5]),
    .A_N(\Inst_S_IO_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_mux4_1 _078_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .A0(S2MID[6]),
    .A1(S2MID[7]),
    .A2(S2END[0]),
    .A3(S2END[4]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_041_));
 sg13g2_o21ai_1 _079_ (.B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_042_),
    .A1(S2END[6]),
    .A2(\Inst_S_IO_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_o21ai_1 _080_ (.B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_043_),
    .A1(\Inst_S_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_040_));
 sg13g2_nand2b_1 _081_ (.Y(_044_),
    .B(_042_),
    .A_N(_043_));
 sg13g2_o21ai_1 _082_ (.B1(_044_),
    .Y(B_T_top),
    .A1(\Inst_S_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_041_));
 sg13g2_inv_1 _083_ (.Y(_000_),
    .A(S2END[1]));
 sg13g2_inv_1 _084_ (.Y(_001_),
    .A(\Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_mux2_1 _085_ (.A0(S2END[2]),
    .A1(S2END[3]),
    .S(\Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_002_));
 sg13g2_or2_1 _086_ (.X(_003_),
    .B(S2END[0]),
    .A(\Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_a21oi_1 _087_ (.A1(\Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_000_),
    .Y(_004_),
    .B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_a221oi_1 _088_ (.B2(_004_),
    .C1(\Inst_S_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .B1(_003_),
    .A1(\Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_005_),
    .A2(_002_));
 sg13g2_nand2_1 _089_ (.Y(_006_),
    .A(\Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .B(S2END[5]));
 sg13g2_nand2b_1 _090_ (.Y(_007_),
    .B(S2END[4]),
    .A_N(\Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_a21oi_1 _091_ (.A1(_006_),
    .A2(_007_),
    .Y(_008_),
    .B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_nor2b_1 _092_ (.A(S2END[7]),
    .B_N(\Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_009_));
 sg13g2_o21ai_1 _093_ (.B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_010_),
    .A1(\Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(S2END[6]));
 sg13g2_o21ai_1 _094_ (.B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_011_),
    .A1(_009_),
    .A2(_010_));
 sg13g2_o21ai_1 _095_ (.B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .Y(_012_),
    .A1(_008_),
    .A2(_011_));
 sg13g2_mux4_1 _096_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .A0(S2MID[4]),
    .A1(S2MID[5]),
    .A2(S2MID[6]),
    .A3(S2MID[7]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_013_));
 sg13g2_mux4_1 _097_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .A0(S2MID[0]),
    .A1(S2MID[1]),
    .A2(S2MID[2]),
    .A3(S2MID[3]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_014_));
 sg13g2_mux2_1 _098_ (.A0(_014_),
    .A1(_013_),
    .S(\Inst_S_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_015_));
 sg13g2_nand2b_1 _099_ (.Y(_016_),
    .B(_015_),
    .A_N(\Inst_S_IO_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_o21ai_1 _100_ (.B1(_016_),
    .Y(B_I_top),
    .A1(_005_),
    .A2(_012_));
 sg13g2_mux2_1 _101_ (.A0(S2END[2]),
    .A1(S2END[3]),
    .S(\Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_017_));
 sg13g2_or2_1 _102_ (.X(_018_),
    .B(\Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .A(S2END[0]));
 sg13g2_a21oi_1 _103_ (.A1(_000_),
    .A2(\Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .Y(_019_),
    .B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_a221oi_1 _104_ (.B2(_019_),
    .C1(\Inst_S_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .B1(_018_),
    .A1(\Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .Y(_020_),
    .A2(_017_));
 sg13g2_nand2_1 _105_ (.Y(_021_),
    .A(S2END[5]),
    .B(\Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_nand2b_1 _106_ (.Y(_022_),
    .B(S2END[4]),
    .A_N(\Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_a21oi_1 _107_ (.A1(_021_),
    .A2(_022_),
    .Y(_023_),
    .B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_nor2b_1 _108_ (.A(S2END[7]),
    .B_N(\Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .Y(_024_));
 sg13g2_o21ai_1 _109_ (.B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .Y(_025_),
    .A1(S2END[6]),
    .A2(\Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_o21ai_1 _110_ (.B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .Y(_026_),
    .A1(_024_),
    .A2(_025_));
 sg13g2_o21ai_1 _111_ (.B1(\Inst_S_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .Y(_027_),
    .A1(_023_),
    .A2(_026_));
 sg13g2_mux4_1 _112_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(S2MID[0]),
    .A1(S2MID[1]),
    .A2(S2MID[2]),
    .A3(S2MID[3]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_028_));
 sg13g2_mux4_1 _113_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(S2MID[4]),
    .A1(S2MID[5]),
    .A2(S2MID[6]),
    .A3(S2MID[7]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_029_));
 sg13g2_mux2_1 _114_ (.A0(_028_),
    .A1(_029_),
    .S(\Inst_S_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_030_));
 sg13g2_nand2b_1 _115_ (.Y(_031_),
    .B(_030_),
    .A_N(\Inst_S_IO_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_o21ai_1 _116_ (.B1(_031_),
    .Y(A_I_top),
    .A1(_020_),
    .A2(_027_));
 sg13g2_mux4_1 _117_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit17.Q ),
    .A0(S2MID[1]),
    .A1(S2MID[5]),
    .A2(S2MID[3]),
    .A3(S2MID[7]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit16.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG15 ));
 sg13g2_mux4_1 _118_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit15.Q ),
    .A0(S2MID[0]),
    .A1(S2MID[4]),
    .A2(S2MID[2]),
    .A3(S2MID[6]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit14.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG14 ));
 sg13g2_mux4_1 _119_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit12.Q ),
    .A0(S4END[7]),
    .A1(S4END[9]),
    .A2(S4END[11]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit13.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG13 ));
 sg13g2_mux4_1 _120_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(S4END[1]),
    .A1(S4END[3]),
    .A2(S4END[5]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit11.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG12 ));
 sg13g2_mux4_1 _121_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit8.Q ),
    .A0(S4END[6]),
    .A1(S4END[8]),
    .A2(S4END[10]),
    .A3(B_O_top),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit9.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG11 ));
 sg13g2_mux4_1 _122_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(S4END[0]),
    .A1(S4END[2]),
    .A2(S4END[4]),
    .A3(A_O_top),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG10 ));
 sg13g2_mux4_1 _123_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(S4END[1]),
    .A1(S4END[3]),
    .A2(S4END[5]),
    .A3(S4END[7]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG9 ));
 sg13g2_mux4_1 _124_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit3.Q ),
    .A0(S4END[4]),
    .A1(S4END[8]),
    .A2(S4END[6]),
    .A3(S4END[10]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit2.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG8 ));
 sg13g2_mux4_1 _125_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame0_bit1.Q ),
    .A0(S2MID[1]),
    .A1(S2MID[5]),
    .A2(S2MID[3]),
    .A3(S2MID[7]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame0_bit0.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG7 ));
 sg13g2_mux4_1 _126_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit31.Q ),
    .A0(S2MID[0]),
    .A1(S2MID[4]),
    .A2(S2MID[2]),
    .A3(S2MID[6]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit30.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG6 ));
 sg13g2_mux4_1 _127_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(S2END[1]),
    .A1(S2END[3]),
    .A2(S2END[5]),
    .A3(S2END[7]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG5 ));
 sg13g2_mux4_1 _128_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(S2END[0]),
    .A1(S2END[2]),
    .A2(S2END[4]),
    .A3(S2END[6]),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG4 ));
 sg13g2_mux4_1 _129_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(S4END[7]),
    .A1(S4END[9]),
    .A2(S4END[11]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG3 ));
 sg13g2_mux4_1 _130_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(S4END[1]),
    .A1(S4END[3]),
    .A2(S4END[5]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG2 ));
 sg13g2_mux4_1 _131_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(S4END[6]),
    .A1(S4END[8]),
    .A2(S4END[10]),
    .A3(B_O_top),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG1 ));
 sg13g2_mux4_1 _132_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(S4END[0]),
    .A1(S4END[2]),
    .A2(S4END[4]),
    .A3(A_O_top),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Inst_S_IO_switch_matrix.NN4BEG0 ));
 sg13g2_mux4_1 _133_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(S4END[0]),
    .A1(SS4END[0]),
    .A2(SS4END[12]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG15 ));
 sg13g2_mux4_1 _134_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(S4END[1]),
    .A1(SS4END[1]),
    .A2(SS4END[13]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit15.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG14 ));
 sg13g2_mux4_1 _135_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit13.Q ),
    .A0(S1END[0]),
    .A1(SS4END[4]),
    .A2(S4END[4]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit12.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG13 ));
 sg13g2_mux4_1 _136_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit11.Q ),
    .A0(S1END[1]),
    .A1(SS4END[5]),
    .A2(S4END[5]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit10.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG12 ));
 sg13g2_mux4_1 _137_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit9.Q ),
    .A0(S4END[8]),
    .A1(SS4END[12]),
    .A2(SS4END[8]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit8.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG11 ));
 sg13g2_mux4_1 _138_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit7.Q ),
    .A0(S4END[9]),
    .A1(SS4END[13]),
    .A2(SS4END[9]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit6.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG10 ));
 sg13g2_mux4_1 _139_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit4.Q ),
    .A0(S1END[0]),
    .A1(S4END[12]),
    .A2(SS4END[12]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit5.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG9 ));
 sg13g2_mux4_1 _140_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit2.Q ),
    .A0(S1END[1]),
    .A1(S4END[13]),
    .A2(SS4END[13]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit3.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG8 ));
 sg13g2_mux4_1 _141_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame1_bit0.Q ),
    .A0(S4END[2]),
    .A1(SS4END[2]),
    .A2(SS4END[14]),
    .A3(B_O_top),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame1_bit1.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG7 ));
 sg13g2_mux4_1 _142_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit30.Q ),
    .A0(S4END[3]),
    .A1(SS4END[3]),
    .A2(SS4END[15]),
    .A3(A_O_top),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit31.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG6 ));
 sg13g2_mux4_1 _143_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit29.Q ),
    .A0(S1END[3]),
    .A1(SS4END[6]),
    .A2(S4END[6]),
    .A3(B_O_top),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit28.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG5 ));
 sg13g2_mux4_1 _144_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit27.Q ),
    .A0(S1END[2]),
    .A1(SS4END[7]),
    .A2(S4END[7]),
    .A3(A_O_top),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit26.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG4 ));
 sg13g2_mux4_1 _145_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit25.Q ),
    .A0(S4END[10]),
    .A1(SS4END[14]),
    .A2(SS4END[10]),
    .A3(B_O_top),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit24.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG3 ));
 sg13g2_mux4_1 _146_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit23.Q ),
    .A0(S4END[11]),
    .A1(SS4END[15]),
    .A2(SS4END[11]),
    .A3(A_O_top),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit22.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG2 ));
 sg13g2_mux4_1 _147_ (.S0(\Inst_S_IO_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(S1END[3]),
    .A1(S4END[14]),
    .A2(SS4END[14]),
    .A3(B_O_top),
    .S1(\Inst_S_IO_ConfigMem.Inst_frame2_bit21.Q ),
    .X(\Inst_S_IO_switch_matrix.N4BEG1 ));
 sg13g2_dlhq_1 _148_ (.D(FrameData[6]),
    .GATE(FrameStrobe[3]),
    .Q(A_config_C_bit0));
 sg13g2_dlhq_1 _149_ (.D(FrameData[7]),
    .GATE(FrameStrobe[3]),
    .Q(A_config_C_bit1));
 sg13g2_dlhq_1 _150_ (.D(FrameData[8]),
    .GATE(FrameStrobe[3]),
    .Q(A_config_C_bit2));
 sg13g2_dlhq_1 _151_ (.D(FrameData[9]),
    .GATE(FrameStrobe[3]),
    .Q(A_config_C_bit3));
 sg13g2_dlhq_1 _152_ (.D(FrameData[10]),
    .GATE(FrameStrobe[3]),
    .Q(B_config_C_bit0));
 sg13g2_dlhq_1 _153_ (.D(FrameData[11]),
    .GATE(FrameStrobe[3]),
    .Q(B_config_C_bit1));
 sg13g2_dlhq_1 _154_ (.D(FrameData[12]),
    .GATE(FrameStrobe[3]),
    .Q(B_config_C_bit2));
 sg13g2_dlhq_1 _155_ (.D(FrameData[13]),
    .GATE(FrameStrobe[3]),
    .Q(B_config_C_bit3));
 sg13g2_dlhq_1 _156_ (.D(FrameData[14]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_switch_matrix.DEBUG_select_N1BEG0 [0]));
 sg13g2_dlhq_1 _157_ (.D(FrameData[15]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_switch_matrix.DEBUG_select_N1BEG1 [0]));
 sg13g2_dlhq_1 _158_ (.D(FrameData[16]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_switch_matrix.DEBUG_select_N1BEG2 [0]));
 sg13g2_dlhq_1 _159_ (.D(FrameData[17]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_switch_matrix.DEBUG_select_N1BEG3 [0]));
 sg13g2_dlhq_1 _160_ (.D(FrameData[18]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_dlhq_1 _161_ (.D(FrameData[19]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_dlhq_1 _162_ (.D(FrameData[20]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_dlhq_1 _163_ (.D(FrameData[21]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_dlhq_1 _164_ (.D(FrameData[22]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _165_ (.D(FrameData[23]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _166_ (.D(FrameData[24]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _167_ (.D(FrameData[25]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _168_ (.D(FrameData[26]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _169_ (.D(FrameData[27]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _170_ (.D(FrameData[28]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _171_ (.D(FrameData[29]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _172_ (.D(FrameData[30]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _173_ (.D(FrameData[31]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _174_ (.D(FrameData[0]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _175_ (.D(FrameData[1]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _176_ (.D(FrameData[2]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _177_ (.D(FrameData[3]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _178_ (.D(FrameData[4]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _179_ (.D(FrameData[5]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _180_ (.D(FrameData[6]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _181_ (.D(FrameData[7]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _182_ (.D(FrameData[8]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _183_ (.D(FrameData[9]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _184_ (.D(FrameData[10]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _185_ (.D(FrameData[11]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _186_ (.D(FrameData[12]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _187_ (.D(FrameData[13]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _188_ (.D(FrameData[14]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _189_ (.D(FrameData[15]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _190_ (.D(FrameData[16]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _191_ (.D(FrameData[17]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _192_ (.D(FrameData[18]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _193_ (.D(FrameData[19]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _194_ (.D(FrameData[20]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _195_ (.D(FrameData[21]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _196_ (.D(FrameData[22]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _197_ (.D(FrameData[23]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _198_ (.D(FrameData[24]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _199_ (.D(FrameData[25]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _200_ (.D(FrameData[26]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _201_ (.D(FrameData[27]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _202_ (.D(FrameData[28]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _203_ (.D(FrameData[29]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _204_ (.D(FrameData[30]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _205_ (.D(FrameData[31]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _206_ (.D(FrameData[0]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _207_ (.D(FrameData[1]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _208_ (.D(FrameData[2]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _209_ (.D(FrameData[3]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _210_ (.D(FrameData[4]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _211_ (.D(FrameData[5]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _212_ (.D(FrameData[6]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _213_ (.D(FrameData[7]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _214_ (.D(FrameData[8]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _215_ (.D(FrameData[9]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _216_ (.D(FrameData[10]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _217_ (.D(FrameData[11]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _218_ (.D(FrameData[12]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _219_ (.D(FrameData[13]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _220_ (.D(FrameData[14]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _221_ (.D(FrameData[15]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _222_ (.D(FrameData[16]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _223_ (.D(FrameData[17]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _224_ (.D(FrameData[18]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _225_ (.D(FrameData[19]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _226_ (.D(FrameData[20]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _227_ (.D(FrameData[21]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _228_ (.D(FrameData[22]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _229_ (.D(FrameData[23]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _230_ (.D(FrameData[24]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _231_ (.D(FrameData[25]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _232_ (.D(FrameData[26]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _233_ (.D(FrameData[27]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _234_ (.D(FrameData[28]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _235_ (.D(FrameData[29]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _236_ (.D(FrameData[30]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _237_ (.D(FrameData[31]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _238_ (.D(FrameData[0]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _239_ (.D(FrameData[1]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _240_ (.D(FrameData[2]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _241_ (.D(FrameData[3]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _242_ (.D(FrameData[4]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _243_ (.D(FrameData[5]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _244_ (.D(FrameData[6]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _245_ (.D(FrameData[7]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _246_ (.D(FrameData[8]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _247_ (.D(FrameData[9]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _248_ (.D(FrameData[10]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _249_ (.D(FrameData[11]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _250_ (.D(FrameData[12]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _251_ (.D(FrameData[13]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _252_ (.D(FrameData[14]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _253_ (.D(FrameData[15]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _254_ (.D(FrameData[16]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _255_ (.D(FrameData[17]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _256_ (.D(FrameData[18]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _257_ (.D(FrameData[19]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _258_ (.D(FrameData[20]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _259_ (.D(FrameData[21]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _260_ (.D(FrameData[22]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _261_ (.D(FrameData[23]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _262_ (.D(FrameData[24]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _263_ (.D(FrameData[25]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _264_ (.D(FrameData[26]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _265_ (.D(FrameData[27]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _266_ (.D(FrameData[28]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _267_ (.D(FrameData[29]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _268_ (.D(FrameData[30]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _269_ (.D(FrameData[31]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_S_IO_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_dfrbpq_1 _270_ (.RESET_B(_045_),
    .D(A_O_top),
    .Q(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .CLK(clknet_1_1__leaf_UserCLK_regs));
 sg13g2_dfrbpq_1 _271_ (.RESET_B(_046_),
    .D(B_O_top),
    .Q(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .CLK(clknet_1_0__leaf_UserCLK_regs));
 sg13g2_tiehi _272_ (.L_HI(_045_));
 sg13g2_tiehi _273_ (.L_HI(_046_));
 sg13g2_tielo _274_ (.L_LO(Co));
 sg13g2_buf_1 _275_ (.A(FrameData[0]),
    .X(FrameData_O[0]));
 sg13g2_buf_1 _276_ (.A(FrameData[1]),
    .X(FrameData_O[1]));
 sg13g2_buf_1 _277_ (.A(FrameData[2]),
    .X(FrameData_O[2]));
 sg13g2_buf_1 _278_ (.A(FrameData[3]),
    .X(FrameData_O[3]));
 sg13g2_buf_1 _279_ (.A(FrameData[4]),
    .X(FrameData_O[4]));
 sg13g2_buf_1 _280_ (.A(FrameData[5]),
    .X(FrameData_O[5]));
 sg13g2_buf_1 _281_ (.A(FrameData[6]),
    .X(FrameData_O[6]));
 sg13g2_buf_1 _282_ (.A(FrameData[7]),
    .X(FrameData_O[7]));
 sg13g2_buf_1 _283_ (.A(FrameData[8]),
    .X(FrameData_O[8]));
 sg13g2_buf_1 _284_ (.A(FrameData[9]),
    .X(FrameData_O[9]));
 sg13g2_buf_1 _285_ (.A(FrameData[10]),
    .X(FrameData_O[10]));
 sg13g2_buf_1 _286_ (.A(FrameData[11]),
    .X(FrameData_O[11]));
 sg13g2_buf_1 _287_ (.A(FrameData[12]),
    .X(FrameData_O[12]));
 sg13g2_buf_1 _288_ (.A(FrameData[13]),
    .X(FrameData_O[13]));
 sg13g2_buf_1 _289_ (.A(FrameData[14]),
    .X(FrameData_O[14]));
 sg13g2_buf_1 _290_ (.A(FrameData[15]),
    .X(FrameData_O[15]));
 sg13g2_buf_1 _291_ (.A(FrameData[16]),
    .X(FrameData_O[16]));
 sg13g2_buf_1 _292_ (.A(FrameData[17]),
    .X(FrameData_O[17]));
 sg13g2_buf_1 _293_ (.A(FrameData[18]),
    .X(FrameData_O[18]));
 sg13g2_buf_1 _294_ (.A(FrameData[19]),
    .X(FrameData_O[19]));
 sg13g2_buf_1 _295_ (.A(FrameData[20]),
    .X(FrameData_O[20]));
 sg13g2_buf_1 _296_ (.A(FrameData[21]),
    .X(FrameData_O[21]));
 sg13g2_buf_1 _297_ (.A(FrameData[22]),
    .X(FrameData_O[22]));
 sg13g2_buf_1 _298_ (.A(FrameData[23]),
    .X(FrameData_O[23]));
 sg13g2_buf_1 _299_ (.A(FrameData[24]),
    .X(FrameData_O[24]));
 sg13g2_buf_1 _300_ (.A(FrameData[25]),
    .X(FrameData_O[25]));
 sg13g2_buf_1 _301_ (.A(FrameData[26]),
    .X(FrameData_O[26]));
 sg13g2_buf_1 _302_ (.A(FrameData[27]),
    .X(FrameData_O[27]));
 sg13g2_buf_1 _303_ (.A(FrameData[28]),
    .X(FrameData_O[28]));
 sg13g2_buf_1 _304_ (.A(FrameData[29]),
    .X(FrameData_O[29]));
 sg13g2_buf_1 _305_ (.A(FrameData[30]),
    .X(FrameData_O[30]));
 sg13g2_buf_1 _306_ (.A(FrameData[31]),
    .X(FrameData_O[31]));
 sg13g2_buf_1 _307_ (.A(FrameStrobe[0]),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 _308_ (.A(FrameStrobe[1]),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 _309_ (.A(FrameStrobe[2]),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 _310_ (.A(FrameStrobe[3]),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 _311_ (.A(FrameStrobe[4]),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 _312_ (.A(FrameStrobe[5]),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 _313_ (.A(FrameStrobe[6]),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 _314_ (.A(FrameStrobe[7]),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 _315_ (.A(FrameStrobe[8]),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 _316_ (.A(FrameStrobe[9]),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 _317_ (.A(FrameStrobe[10]),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 _318_ (.A(FrameStrobe[11]),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 _319_ (.A(FrameStrobe[12]),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 _320_ (.A(FrameStrobe[13]),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 _321_ (.A(FrameStrobe[14]),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 _322_ (.A(FrameStrobe[15]),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 _323_ (.A(FrameStrobe[16]),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 _324_ (.A(FrameStrobe[17]),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 _325_ (.A(FrameStrobe[18]),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 _326_ (.A(FrameStrobe[19]),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 _327_ (.A(\Inst_S_IO_switch_matrix.N1BEG0 ),
    .X(N1BEG[0]));
 sg13g2_buf_1 _328_ (.A(\Inst_S_IO_switch_matrix.N1BEG1 ),
    .X(N1BEG[1]));
 sg13g2_buf_1 _329_ (.A(\Inst_S_IO_switch_matrix.N1BEG2 ),
    .X(N1BEG[2]));
 sg13g2_buf_1 _330_ (.A(\Inst_S_IO_switch_matrix.N1BEG3 ),
    .X(N1BEG[3]));
 sg13g2_buf_1 _331_ (.A(\Inst_S_IO_switch_matrix.N2BEG0 ),
    .X(N2BEG[0]));
 sg13g2_buf_1 _332_ (.A(\Inst_S_IO_switch_matrix.N2BEG1 ),
    .X(N2BEG[1]));
 sg13g2_buf_1 _333_ (.A(\Inst_S_IO_switch_matrix.N2BEG2 ),
    .X(N2BEG[2]));
 sg13g2_buf_1 _334_ (.A(\Inst_S_IO_switch_matrix.N2BEG3 ),
    .X(N2BEG[3]));
 sg13g2_buf_1 _335_ (.A(\Inst_S_IO_switch_matrix.N2BEG4 ),
    .X(N2BEG[4]));
 sg13g2_buf_1 _336_ (.A(\Inst_S_IO_switch_matrix.N2BEG5 ),
    .X(N2BEG[5]));
 sg13g2_buf_1 _337_ (.A(\Inst_S_IO_switch_matrix.N2BEG6 ),
    .X(N2BEG[6]));
 sg13g2_buf_1 _338_ (.A(\Inst_S_IO_switch_matrix.N2BEG7 ),
    .X(N2BEG[7]));
 sg13g2_buf_1 _339_ (.A(\Inst_S_IO_switch_matrix.N2BEGb0 ),
    .X(N2BEGb[0]));
 sg13g2_buf_1 _340_ (.A(\Inst_S_IO_switch_matrix.N2BEGb1 ),
    .X(N2BEGb[1]));
 sg13g2_buf_1 _341_ (.A(\Inst_S_IO_switch_matrix.N2BEGb2 ),
    .X(N2BEGb[2]));
 sg13g2_buf_1 _342_ (.A(\Inst_S_IO_switch_matrix.N2BEGb3 ),
    .X(N2BEGb[3]));
 sg13g2_buf_1 _343_ (.A(\Inst_S_IO_switch_matrix.N2BEGb4 ),
    .X(N2BEGb[4]));
 sg13g2_buf_1 _344_ (.A(\Inst_S_IO_switch_matrix.N2BEGb5 ),
    .X(N2BEGb[5]));
 sg13g2_buf_1 _345_ (.A(\Inst_S_IO_switch_matrix.N2BEGb6 ),
    .X(N2BEGb[6]));
 sg13g2_buf_1 _346_ (.A(\Inst_S_IO_switch_matrix.N2BEGb7 ),
    .X(N2BEGb[7]));
 sg13g2_buf_1 _347_ (.A(\Inst_S_IO_switch_matrix.N4BEG0 ),
    .X(N4BEG[0]));
 sg13g2_buf_1 _348_ (.A(\Inst_S_IO_switch_matrix.N4BEG1 ),
    .X(N4BEG[1]));
 sg13g2_buf_1 _349_ (.A(\Inst_S_IO_switch_matrix.N4BEG2 ),
    .X(N4BEG[2]));
 sg13g2_buf_1 _350_ (.A(\Inst_S_IO_switch_matrix.N4BEG3 ),
    .X(N4BEG[3]));
 sg13g2_buf_1 _351_ (.A(\Inst_S_IO_switch_matrix.N4BEG4 ),
    .X(N4BEG[4]));
 sg13g2_buf_1 _352_ (.A(\Inst_S_IO_switch_matrix.N4BEG5 ),
    .X(N4BEG[5]));
 sg13g2_buf_1 _353_ (.A(\Inst_S_IO_switch_matrix.N4BEG6 ),
    .X(N4BEG[6]));
 sg13g2_buf_1 _354_ (.A(\Inst_S_IO_switch_matrix.N4BEG7 ),
    .X(N4BEG[7]));
 sg13g2_buf_1 _355_ (.A(\Inst_S_IO_switch_matrix.N4BEG8 ),
    .X(N4BEG[8]));
 sg13g2_buf_1 _356_ (.A(\Inst_S_IO_switch_matrix.N4BEG9 ),
    .X(N4BEG[9]));
 sg13g2_buf_1 _357_ (.A(\Inst_S_IO_switch_matrix.N4BEG10 ),
    .X(N4BEG[10]));
 sg13g2_buf_1 _358_ (.A(\Inst_S_IO_switch_matrix.N4BEG11 ),
    .X(N4BEG[11]));
 sg13g2_buf_1 _359_ (.A(\Inst_S_IO_switch_matrix.N4BEG12 ),
    .X(N4BEG[12]));
 sg13g2_buf_1 _360_ (.A(\Inst_S_IO_switch_matrix.N4BEG13 ),
    .X(N4BEG[13]));
 sg13g2_buf_1 _361_ (.A(\Inst_S_IO_switch_matrix.N4BEG14 ),
    .X(N4BEG[14]));
 sg13g2_buf_1 _362_ (.A(\Inst_S_IO_switch_matrix.N4BEG15 ),
    .X(N4BEG[15]));
 sg13g2_buf_1 _363_ (.A(\Inst_S_IO_switch_matrix.NN4BEG0 ),
    .X(NN4BEG[0]));
 sg13g2_buf_1 _364_ (.A(\Inst_S_IO_switch_matrix.NN4BEG1 ),
    .X(NN4BEG[1]));
 sg13g2_buf_1 _365_ (.A(\Inst_S_IO_switch_matrix.NN4BEG2 ),
    .X(NN4BEG[2]));
 sg13g2_buf_1 _366_ (.A(\Inst_S_IO_switch_matrix.NN4BEG3 ),
    .X(NN4BEG[3]));
 sg13g2_buf_1 _367_ (.A(\Inst_S_IO_switch_matrix.NN4BEG4 ),
    .X(NN4BEG[4]));
 sg13g2_buf_1 _368_ (.A(\Inst_S_IO_switch_matrix.NN4BEG5 ),
    .X(NN4BEG[5]));
 sg13g2_buf_1 _369_ (.A(\Inst_S_IO_switch_matrix.NN4BEG6 ),
    .X(NN4BEG[6]));
 sg13g2_buf_1 _370_ (.A(\Inst_S_IO_switch_matrix.NN4BEG7 ),
    .X(NN4BEG[7]));
 sg13g2_buf_1 _371_ (.A(\Inst_S_IO_switch_matrix.NN4BEG8 ),
    .X(NN4BEG[8]));
 sg13g2_buf_1 _372_ (.A(\Inst_S_IO_switch_matrix.NN4BEG9 ),
    .X(NN4BEG[9]));
 sg13g2_buf_1 _373_ (.A(\Inst_S_IO_switch_matrix.NN4BEG10 ),
    .X(NN4BEG[10]));
 sg13g2_buf_1 _374_ (.A(\Inst_S_IO_switch_matrix.NN4BEG11 ),
    .X(NN4BEG[11]));
 sg13g2_buf_1 _375_ (.A(\Inst_S_IO_switch_matrix.NN4BEG12 ),
    .X(NN4BEG[12]));
 sg13g2_buf_1 _376_ (.A(\Inst_S_IO_switch_matrix.NN4BEG13 ),
    .X(NN4BEG[13]));
 sg13g2_buf_1 _377_ (.A(\Inst_S_IO_switch_matrix.NN4BEG14 ),
    .X(NN4BEG[14]));
 sg13g2_buf_1 _378_ (.A(\Inst_S_IO_switch_matrix.NN4BEG15 ),
    .X(NN4BEG[15]));
 sg13g2_buf_1 _379_ (.A(clknet_1_0__leaf_UserCLK),
    .X(UserCLKo));
 sg13g2_buf_8 clkbuf_regs_0_UserCLK (.A(UserCLK),
    .X(UserCLK_regs));
 sg13g2_buf_8 clkbuf_0_UserCLK (.A(UserCLK),
    .X(clknet_0_UserCLK));
 sg13g2_buf_8 clkbuf_1_0__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_0__leaf_UserCLK));
 sg13g2_buf_8 clkbuf_0_UserCLK_regs (.A(UserCLK_regs),
    .X(clknet_0_UserCLK_regs));
 sg13g2_buf_8 clkbuf_1_0__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_0__leaf_UserCLK_regs));
 sg13g2_buf_8 clkbuf_1_1__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_1__leaf_UserCLK_regs));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_4 FILLER_0_7 ();
 sg13g2_fill_2 FILLER_0_11 ();
 sg13g2_fill_1 FILLER_0_30 ();
 sg13g2_decap_8 FILLER_0_41 ();
 sg13g2_decap_8 FILLER_0_48 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_fill_2 FILLER_0_154 ();
 sg13g2_fill_1 FILLER_0_156 ();
 sg13g2_fill_1 FILLER_0_178 ();
 sg13g2_decap_4 FILLER_0_230 ();
 sg13g2_fill_1 FILLER_0_251 ();
 sg13g2_decap_4 FILLER_0_269 ();
 sg13g2_fill_2 FILLER_0_273 ();
 sg13g2_fill_2 FILLER_0_292 ();
 sg13g2_fill_2 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_4 FILLER_0_404 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_fill_2 FILLER_0_421 ();
 sg13g2_fill_1 FILLER_0_423 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_24 ();
 sg13g2_fill_1 FILLER_1_26 ();
 sg13g2_decap_4 FILLER_1_59 ();
 sg13g2_fill_1 FILLER_1_165 ();
 sg13g2_decap_8 FILLER_1_193 ();
 sg13g2_decap_8 FILLER_1_200 ();
 sg13g2_fill_2 FILLER_1_207 ();
 sg13g2_fill_1 FILLER_1_277 ();
 sg13g2_fill_2 FILLER_1_320 ();
 sg13g2_fill_1 FILLER_1_322 ();
 sg13g2_fill_1 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_389 ();
 sg13g2_fill_1 FILLER_1_412 ();
 sg13g2_fill_2 FILLER_1_421 ();
 sg13g2_fill_1 FILLER_1_423 ();
 sg13g2_decap_4 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_48 ();
 sg13g2_decap_8 FILLER_2_72 ();
 sg13g2_fill_2 FILLER_2_79 ();
 sg13g2_fill_1 FILLER_2_81 ();
 sg13g2_fill_2 FILLER_2_99 ();
 sg13g2_fill_1 FILLER_2_101 ();
 sg13g2_fill_2 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_125 ();
 sg13g2_decap_4 FILLER_2_132 ();
 sg13g2_fill_1 FILLER_2_136 ();
 sg13g2_decap_4 FILLER_2_213 ();
 sg13g2_decap_4 FILLER_2_247 ();
 sg13g2_fill_1 FILLER_2_251 ();
 sg13g2_fill_1 FILLER_2_273 ();
 sg13g2_decap_4 FILLER_2_291 ();
 sg13g2_fill_1 FILLER_2_295 ();
 sg13g2_fill_2 FILLER_2_313 ();
 sg13g2_decap_4 FILLER_2_332 ();
 sg13g2_fill_2 FILLER_2_336 ();
 sg13g2_fill_2 FILLER_2_355 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_fill_2 FILLER_2_421 ();
 sg13g2_fill_1 FILLER_2_423 ();
 sg13g2_decap_4 FILLER_3_0 ();
 sg13g2_decap_4 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_43 ();
 sg13g2_decap_8 FILLER_3_50 ();
 sg13g2_decap_8 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_4 FILLER_3_109 ();
 sg13g2_fill_2 FILLER_3_113 ();
 sg13g2_decap_4 FILLER_3_166 ();
 sg13g2_fill_1 FILLER_3_195 ();
 sg13g2_decap_8 FILLER_3_213 ();
 sg13g2_fill_2 FILLER_3_220 ();
 sg13g2_fill_1 FILLER_3_222 ();
 sg13g2_fill_2 FILLER_3_291 ();
 sg13g2_fill_2 FILLER_3_310 ();
 sg13g2_decap_4 FILLER_3_320 ();
 sg13g2_fill_2 FILLER_3_324 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_fill_1 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_4 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_21 ();
 sg13g2_fill_1 FILLER_4_23 ();
 sg13g2_decap_4 FILLER_4_54 ();
 sg13g2_decap_8 FILLER_4_79 ();
 sg13g2_decap_8 FILLER_4_86 ();
 sg13g2_decap_8 FILLER_4_93 ();
 sg13g2_fill_2 FILLER_4_121 ();
 sg13g2_fill_2 FILLER_4_144 ();
 sg13g2_fill_1 FILLER_4_146 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_4 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_214 ();
 sg13g2_decap_8 FILLER_4_221 ();
 sg13g2_fill_2 FILLER_4_228 ();
 sg13g2_fill_2 FILLER_4_272 ();
 sg13g2_fill_2 FILLER_4_304 ();
 sg13g2_fill_2 FILLER_4_323 ();
 sg13g2_fill_1 FILLER_4_325 ();
 sg13g2_fill_2 FILLER_4_347 ();
 sg13g2_fill_1 FILLER_4_349 ();
 sg13g2_decap_4 FILLER_4_375 ();
 sg13g2_fill_2 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_fill_2 FILLER_4_421 ();
 sg13g2_fill_1 FILLER_4_423 ();
 sg13g2_decap_4 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_4 ();
 sg13g2_fill_2 FILLER_5_22 ();
 sg13g2_fill_1 FILLER_5_24 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_fill_1 FILLER_5_84 ();
 sg13g2_fill_2 FILLER_5_106 ();
 sg13g2_fill_1 FILLER_5_108 ();
 sg13g2_decap_4 FILLER_5_134 ();
 sg13g2_fill_2 FILLER_5_138 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_4 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_170 ();
 sg13g2_fill_1 FILLER_5_177 ();
 sg13g2_decap_8 FILLER_5_195 ();
 sg13g2_fill_2 FILLER_5_202 ();
 sg13g2_fill_1 FILLER_5_204 ();
 sg13g2_decap_4 FILLER_5_230 ();
 sg13g2_fill_2 FILLER_5_234 ();
 sg13g2_decap_8 FILLER_5_253 ();
 sg13g2_decap_8 FILLER_5_260 ();
 sg13g2_fill_2 FILLER_5_267 ();
 sg13g2_decap_8 FILLER_5_311 ();
 sg13g2_fill_2 FILLER_5_318 ();
 sg13g2_fill_1 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_fill_2 FILLER_5_373 ();
 sg13g2_fill_2 FILLER_5_421 ();
 sg13g2_fill_1 FILLER_5_423 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_fill_2 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_30 ();
 sg13g2_fill_2 FILLER_6_39 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_4 FILLER_6_205 ();
 sg13g2_decap_8 FILLER_6_243 ();
 sg13g2_decap_4 FILLER_6_250 ();
 sg13g2_fill_2 FILLER_6_254 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_fill_2 FILLER_6_280 ();
 sg13g2_fill_1 FILLER_6_286 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_fill_1 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_fill_2 FILLER_6_410 ();
 sg13g2_fill_1 FILLER_6_412 ();
 sg13g2_fill_2 FILLER_6_421 ();
 sg13g2_fill_1 FILLER_6_423 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_14 ();
 sg13g2_fill_1 FILLER_7_33 ();
 sg13g2_fill_2 FILLER_7_92 ();
 sg13g2_fill_1 FILLER_7_94 ();
 sg13g2_fill_2 FILLER_7_137 ();
 sg13g2_fill_1 FILLER_7_139 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_fill_2 FILLER_7_168 ();
 sg13g2_fill_1 FILLER_7_170 ();
 sg13g2_fill_2 FILLER_7_188 ();
 sg13g2_decap_4 FILLER_7_232 ();
 sg13g2_decap_8 FILLER_7_257 ();
 sg13g2_decap_4 FILLER_7_264 ();
 sg13g2_fill_1 FILLER_7_268 ();
 sg13g2_fill_2 FILLER_7_311 ();
 sg13g2_fill_1 FILLER_7_313 ();
 sg13g2_decap_8 FILLER_7_352 ();
 sg13g2_decap_8 FILLER_7_363 ();
 sg13g2_decap_8 FILLER_7_370 ();
 sg13g2_fill_2 FILLER_7_377 ();
 sg13g2_fill_2 FILLER_7_383 ();
 sg13g2_fill_2 FILLER_7_410 ();
 sg13g2_fill_1 FILLER_7_412 ();
 sg13g2_fill_2 FILLER_7_421 ();
 sg13g2_fill_1 FILLER_7_423 ();
 sg13g2_decap_4 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_4 ();
 sg13g2_fill_2 FILLER_8_22 ();
 sg13g2_fill_1 FILLER_8_24 ();
 sg13g2_decap_8 FILLER_8_57 ();
 sg13g2_decap_8 FILLER_8_64 ();
 sg13g2_decap_8 FILLER_8_113 ();
 sg13g2_decap_4 FILLER_8_124 ();
 sg13g2_fill_2 FILLER_8_128 ();
 sg13g2_fill_2 FILLER_8_134 ();
 sg13g2_fill_1 FILLER_8_136 ();
 sg13g2_decap_4 FILLER_8_188 ();
 sg13g2_fill_1 FILLER_8_209 ();
 sg13g2_decap_8 FILLER_8_227 ();
 sg13g2_decap_8 FILLER_8_234 ();
 sg13g2_fill_1 FILLER_8_258 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_fill_2 FILLER_8_300 ();
 sg13g2_fill_1 FILLER_8_319 ();
 sg13g2_fill_1 FILLER_8_337 ();
 sg13g2_decap_4 FILLER_8_342 ();
 sg13g2_fill_1 FILLER_8_346 ();
 sg13g2_fill_1 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_4 FILLER_8_389 ();
 sg13g2_fill_2 FILLER_8_410 ();
 sg13g2_fill_1 FILLER_8_412 ();
 sg13g2_fill_2 FILLER_8_421 ();
 sg13g2_fill_1 FILLER_8_423 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_24 ();
 sg13g2_fill_2 FILLER_9_41 ();
 sg13g2_decap_8 FILLER_9_69 ();
 sg13g2_decap_8 FILLER_9_76 ();
 sg13g2_fill_2 FILLER_9_83 ();
 sg13g2_fill_1 FILLER_9_106 ();
 sg13g2_decap_4 FILLER_9_115 ();
 sg13g2_fill_1 FILLER_9_119 ();
 sg13g2_fill_1 FILLER_9_137 ();
 sg13g2_decap_4 FILLER_9_159 ();
 sg13g2_fill_2 FILLER_9_167 ();
 sg13g2_fill_2 FILLER_9_194 ();
 sg13g2_decap_4 FILLER_9_200 ();
 sg13g2_fill_1 FILLER_9_204 ();
 sg13g2_decap_8 FILLER_9_230 ();
 sg13g2_fill_1 FILLER_9_237 ();
 sg13g2_fill_2 FILLER_9_276 ();
 sg13g2_fill_1 FILLER_9_278 ();
 sg13g2_fill_1 FILLER_9_296 ();
 sg13g2_decap_4 FILLER_9_318 ();
 sg13g2_fill_1 FILLER_9_322 ();
 sg13g2_fill_2 FILLER_9_331 ();
 sg13g2_fill_1 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_351 ();
 sg13g2_decap_4 FILLER_9_358 ();
 sg13g2_fill_2 FILLER_9_362 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_fill_2 FILLER_9_421 ();
 sg13g2_fill_1 FILLER_9_423 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_43 ();
 sg13g2_fill_1 FILLER_10_49 ();
 sg13g2_decap_4 FILLER_10_71 ();
 sg13g2_fill_2 FILLER_10_96 ();
 sg13g2_fill_1 FILLER_10_98 ();
 sg13g2_fill_2 FILLER_10_120 ();
 sg13g2_fill_1 FILLER_10_122 ();
 sg13g2_fill_2 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_163 ();
 sg13g2_fill_1 FILLER_10_202 ();
 sg13g2_fill_2 FILLER_10_241 ();
 sg13g2_fill_1 FILLER_10_247 ();
 sg13g2_fill_1 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_fill_1 FILLER_10_322 ();
 sg13g2_fill_1 FILLER_10_344 ();
 sg13g2_fill_2 FILLER_10_355 ();
 sg13g2_fill_1 FILLER_10_357 ();
 sg13g2_decap_4 FILLER_10_396 ();
 sg13g2_fill_1 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_421 ();
 sg13g2_fill_1 FILLER_10_423 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_118 ();
 sg13g2_decap_8 FILLER_11_125 ();
 sg13g2_fill_2 FILLER_11_132 ();
 sg13g2_fill_1 FILLER_11_134 ();
 sg13g2_decap_4 FILLER_11_139 ();
 sg13g2_fill_2 FILLER_11_160 ();
 sg13g2_fill_1 FILLER_11_162 ();
 sg13g2_decap_8 FILLER_11_167 ();
 sg13g2_decap_8 FILLER_11_174 ();
 sg13g2_fill_2 FILLER_11_181 ();
 sg13g2_decap_8 FILLER_11_204 ();
 sg13g2_decap_8 FILLER_11_211 ();
 sg13g2_fill_1 FILLER_11_218 ();
 sg13g2_fill_1 FILLER_11_223 ();
 sg13g2_decap_8 FILLER_11_258 ();
 sg13g2_fill_2 FILLER_11_265 ();
 sg13g2_fill_1 FILLER_11_267 ();
 sg13g2_decap_8 FILLER_11_285 ();
 sg13g2_decap_4 FILLER_11_292 ();
 sg13g2_fill_1 FILLER_11_329 ();
 sg13g2_decap_4 FILLER_11_347 ();
 sg13g2_fill_1 FILLER_11_351 ();
 sg13g2_decap_4 FILLER_11_369 ();
 sg13g2_fill_2 FILLER_11_377 ();
 sg13g2_fill_2 FILLER_11_383 ();
 sg13g2_fill_1 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_410 ();
 sg13g2_fill_1 FILLER_11_412 ();
 sg13g2_fill_2 FILLER_11_421 ();
 sg13g2_fill_1 FILLER_11_423 ();
endmodule
